
module memc_Size16_7 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n214, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1, n2, n3, n4, n5, n6, n7, n8,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n288, n290, n292, n294, n296, n298, n300, n302,
         n304, n306, n308, n310, n312, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1162), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1161), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1160), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1159), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1158), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1157), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1156), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1155), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1154), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1153), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1152), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1151), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1150), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1149), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1148), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1147), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1146), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1145), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1144), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1143), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1142), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1141), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1140), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1139), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1138), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1137), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1136), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1135), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1134), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1133), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1132), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1131), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1130), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1129), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1128), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1127), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1126), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1125), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1124), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1123), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1122), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1121), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1120), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1119), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1118), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1117), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1116), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1115), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1114), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1113), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1112), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1111), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1110), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1109), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1108), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1107), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1106), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1105), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1104), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1103), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1102), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1101), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1100), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1099), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1098), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1097), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1096), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1095), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1094), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1093), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1092), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1091), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1090), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1089), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1088), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1087), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1085), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1083), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1082), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1081), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1080), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1079), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1078), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1077), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1076), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1075), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1074), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1073), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1072), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1071), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1070), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1069), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1068), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1067), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1066), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1065), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1064), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1063), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1062), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1061), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1060), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1059), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1058), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1057), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1056), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1055), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1054), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1053), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1052), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1051), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1050), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1049), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1048), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1047), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1046), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1045), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1044), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1043), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1042), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1041), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1040), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1039), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1038), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1037), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1036), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1035), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1034), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1033), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1032), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1031), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1030), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1029), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1028), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1027), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1026), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1025), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1024), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1023), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1022), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1021), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1020), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1019), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1018), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1017), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1016), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1015), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1014), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1013), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1012), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1011), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1010), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1009), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1008), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1007), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1006), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1005), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1004), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1003), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1002), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1001), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1000), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n999), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n998), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n997), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n996), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n995), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n994), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n993), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n992), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n991), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n990), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n989), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n988), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n987), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n986), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n985), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n984), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n983), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n982), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n981), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n980), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n979), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n978), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n977), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n976), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n975), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n974), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n973), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n972), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n971), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n970), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n969), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n968), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n967), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n966), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n965), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n964), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n963), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n962), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n961), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n960), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n959), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n958), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n957), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n956), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n955), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n954), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n953), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n952), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n951), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n950), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n949), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n948), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n947), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n946), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n945), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n944), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n943), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n942), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n941), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n940), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n939), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n938), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n937), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n936), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n935), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n934), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n933), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n932), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n931), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n930), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n929), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n928), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n927), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n926), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n925), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n924), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n923), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n922), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n921), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n920), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n919), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n918), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n917), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n916), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n915), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n914), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n913), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n912), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n911), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n910), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n909), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n908), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n907), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n906), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n905), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n904), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n903), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n902), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n901), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n900), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n899), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n898), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n897), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n896), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n895), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n894), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n893), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n892), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n891), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n890), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n889), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n888), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n887), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n886), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n885), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n884), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n883), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n882), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n881), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n880), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n879), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n878), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n877), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n876), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n875), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n874), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n873), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n872), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n871), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n870), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n869), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n868), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n867), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n866), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n865), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n864), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n863), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n862), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n861), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n860), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n859), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n858), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n857), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n856), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n855), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n854), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n853), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n852), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n851), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n850), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n849), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n848), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n847), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n846), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n845), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n844), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n843), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n842), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n841), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n840), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n839), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n838), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n837), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n836), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n835), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n834), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n833), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n832), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n831), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n830), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n829), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n828), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n827), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n826), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n825), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n824), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n823), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n822), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n821), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n820), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n819), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n818), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n817), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n816), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n815), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n814), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n813), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n812), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n811), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n810), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n809), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n808), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n807), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n806), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n805), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n804), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n803), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n802), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n801), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n800), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n799), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n798), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n797), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n796), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n795), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n794), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n793), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n792), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n791), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n790), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n789), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n788), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n787), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n786), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n785), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n784), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n783), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n782), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n781), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n780), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n779), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n778), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n777), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n776), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n775), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n774), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n773), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n772), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n771), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n770), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n769), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n768), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n767), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n766), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n765), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n764), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n763), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n762), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n761), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n760), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n759), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n758), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n757), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n756), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n755), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n754), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n753), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n752), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n751), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n750), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n749), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n748), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n747), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n746), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n745), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n744), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n743), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n742), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n741), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n740), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n739), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n738), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n737), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n736), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n735), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n734), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n733), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n732), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n731), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n730), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n729), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n728), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n727), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n726), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n725), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n724), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n723), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n722), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n721), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n720), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n719), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n718), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n717), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n716), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n715), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n714), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n713), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n712), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n711), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n710), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n709), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n708), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n707), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n706), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n705), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n704), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n703), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n702), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n701), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n700), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n699), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n698), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n697), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n696), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n695), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n694), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n693), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n692), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n691), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n690), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n689), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n688), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n687), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n686), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n685), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n684), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n683), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n682), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n681), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n680), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n679), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n678), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n677), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n676), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n675), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n674), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n673), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n672), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n671), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n670), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n669), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n668), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n667), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n666), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n665), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n664), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n663), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n662), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n661), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n660), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n659), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n658), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n657), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n656), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n655), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n654), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n653), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n652), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n651), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n214) );
  INVX1 U2 ( .A(n274), .Y(n1) );
  INVX2 U3 ( .A(n282), .Y(n283) );
  INVX2 U4 ( .A(n284), .Y(n285) );
  INVX2 U5 ( .A(n277), .Y(n278) );
  INVX4 U6 ( .A(n280), .Y(n281) );
  INVX4 U7 ( .A(n623), .Y(n624) );
  INVX4 U8 ( .A(n625), .Y(n626) );
  INVX4 U9 ( .A(n621), .Y(n622) );
  INVX4 U10 ( .A(n627), .Y(n628) );
  INVX4 U11 ( .A(n616), .Y(n617) );
  INVX4 U12 ( .A(n631), .Y(n632) );
  INVX4 U13 ( .A(n629), .Y(n630) );
  INVX4 U14 ( .A(n316), .Y(n317) );
  INVX4 U15 ( .A(n314), .Y(n315) );
  INVX4 U16 ( .A(n275), .Y(n276) );
  INVX1 U17 ( .A(n2338), .Y(n2188) );
  INVX1 U18 ( .A(n2338), .Y(n2187) );
  INVX1 U19 ( .A(n2338), .Y(n2186) );
  INVX1 U20 ( .A(n2342), .Y(n2182) );
  INVX1 U21 ( .A(n2340), .Y(n2183) );
  INVX1 U22 ( .A(n2342), .Y(n2181) );
  INVX1 U23 ( .A(n2337), .Y(n2204) );
  INVX2 U24 ( .A(n2192), .Y(n2193) );
  INVX1 U25 ( .A(n2338), .Y(n2190) );
  INVX1 U26 ( .A(n2338), .Y(n2189) );
  INVX2 U27 ( .A(n2337), .Y(n2199) );
  INVX1 U28 ( .A(n2172), .Y(N25) );
  INVX1 U29 ( .A(n2173), .Y(N24) );
  INVX1 U30 ( .A(n2165), .Y(N32) );
  INVX1 U31 ( .A(n2166), .Y(N31) );
  INVX1 U32 ( .A(n2167), .Y(N30) );
  INVX1 U33 ( .A(n2168), .Y(N29) );
  INVX1 U34 ( .A(n2169), .Y(N28) );
  INVX1 U35 ( .A(n2170), .Y(N27) );
  INVX1 U36 ( .A(n2171), .Y(N26) );
  INVX1 U37 ( .A(n2174), .Y(N23) );
  INVX1 U38 ( .A(n2175), .Y(N22) );
  INVX1 U39 ( .A(n2176), .Y(N21) );
  INVX1 U40 ( .A(n2177), .Y(N20) );
  INVX1 U41 ( .A(n2178), .Y(N19) );
  INVX1 U42 ( .A(n2179), .Y(N18) );
  INVX1 U43 ( .A(n2180), .Y(N17) );
  BUFX2 U44 ( .A(n1630), .Y(n2236) );
  BUFX2 U45 ( .A(n1632), .Y(n2238) );
  BUFX2 U46 ( .A(n1634), .Y(n2240) );
  BUFX2 U47 ( .A(n1636), .Y(n2243) );
  BUFX2 U48 ( .A(n1638), .Y(n2245) );
  BUFX2 U49 ( .A(n1640), .Y(n2247) );
  BUFX2 U50 ( .A(n1642), .Y(n2249) );
  BUFX2 U51 ( .A(n1644), .Y(n2252) );
  BUFX2 U52 ( .A(n1646), .Y(n2254) );
  BUFX2 U53 ( .A(n1648), .Y(n2256) );
  BUFX2 U54 ( .A(n1650), .Y(n2258) );
  BUFX2 U55 ( .A(n1652), .Y(n2260) );
  BUFX2 U56 ( .A(n1654), .Y(n2262) );
  BUFX2 U57 ( .A(n1656), .Y(n2264) );
  BUFX2 U58 ( .A(n1658), .Y(n2268) );
  BUFX2 U59 ( .A(n1660), .Y(n2270) );
  BUFX2 U60 ( .A(n1662), .Y(n2272) );
  BUFX2 U61 ( .A(n1664), .Y(n2274) );
  BUFX2 U62 ( .A(n1666), .Y(n2276) );
  BUFX2 U63 ( .A(n1668), .Y(n2278) );
  BUFX2 U64 ( .A(n1670), .Y(n2280) );
  BUFX2 U65 ( .A(n1672), .Y(n2283) );
  BUFX2 U66 ( .A(n1674), .Y(n2285) );
  BUFX2 U67 ( .A(n1676), .Y(n2287) );
  BUFX2 U68 ( .A(n1678), .Y(n2289) );
  BUFX2 U69 ( .A(n1680), .Y(n2291) );
  BUFX2 U70 ( .A(n1682), .Y(n2293) );
  BUFX2 U71 ( .A(n1684), .Y(n2295) );
  INVX1 U72 ( .A(write), .Y(n2) );
  INVX1 U73 ( .A(write), .Y(n274) );
  INVX1 U74 ( .A(n2338), .Y(n2185) );
  INVX1 U75 ( .A(n2211), .Y(n2212) );
  INVX2 U76 ( .A(N12), .Y(n2338) );
  INVX2 U77 ( .A(n2340), .Y(n2184) );
  INVX4 U78 ( .A(n2334), .Y(n2233) );
  INVX2 U79 ( .A(n2234), .Y(n2205) );
  INVX4 U80 ( .A(n2235), .Y(n2211) );
  BUFX2 U81 ( .A(n1632), .Y(n2239) );
  BUFX2 U82 ( .A(n1636), .Y(n2244) );
  BUFX2 U83 ( .A(n1638), .Y(n2246) );
  INVX1 U84 ( .A(n2342), .Y(n2341) );
  INVX1 U85 ( .A(N14), .Y(n2342) );
  BUFX2 U86 ( .A(n1654), .Y(n2263) );
  BUFX2 U87 ( .A(n1656), .Y(n2265) );
  BUFX2 U88 ( .A(n1674), .Y(n2286) );
  BUFX2 U89 ( .A(n1676), .Y(n2288) );
  INVX1 U90 ( .A(n1627), .Y(n2282) );
  INVX1 U91 ( .A(n1628), .Y(n2297) );
  BUFX2 U92 ( .A(n1652), .Y(n2261) );
  BUFX2 U93 ( .A(n1644), .Y(n2253) );
  BUFX2 U94 ( .A(n1634), .Y(n2241) );
  BUFX2 U95 ( .A(n1640), .Y(n2248) );
  BUFX2 U96 ( .A(n1642), .Y(n2250) );
  BUFX2 U97 ( .A(n1672), .Y(n2284) );
  BUFX2 U98 ( .A(n1678), .Y(n2290) );
  BUFX2 U99 ( .A(n1680), .Y(n2292) );
  BUFX2 U100 ( .A(n1682), .Y(n2294) );
  BUFX2 U101 ( .A(n1684), .Y(n2296) );
  BUFX2 U102 ( .A(n1630), .Y(n2237) );
  BUFX2 U103 ( .A(n1658), .Y(n2269) );
  BUFX2 U104 ( .A(n1660), .Y(n2271) );
  BUFX2 U105 ( .A(n1662), .Y(n2273) );
  BUFX2 U106 ( .A(n1664), .Y(n2275) );
  BUFX2 U107 ( .A(n1666), .Y(n2277) );
  BUFX2 U108 ( .A(n1668), .Y(n2279) );
  BUFX2 U109 ( .A(n1670), .Y(n2281) );
  BUFX2 U110 ( .A(n1646), .Y(n2255) );
  BUFX2 U111 ( .A(n1648), .Y(n2257) );
  BUFX2 U112 ( .A(n1650), .Y(n2259) );
  INVX1 U113 ( .A(n1626), .Y(n2267) );
  INVX1 U114 ( .A(n1625), .Y(n2251) );
  INVX1 U115 ( .A(n2340), .Y(n2339) );
  INVX1 U116 ( .A(N13), .Y(n2340) );
  INVX1 U117 ( .A(rst), .Y(n2333) );
  INVX1 U118 ( .A(n318), .Y(n3) );
  INVX2 U119 ( .A(n639), .Y(n641) );
  INVX2 U120 ( .A(n636), .Y(n638) );
  INVX2 U121 ( .A(n633), .Y(n635) );
  AND2X2 U122 ( .A(\data_in<0> ), .B(n1185), .Y(n4) );
  INVX4 U123 ( .A(n340), .Y(n341) );
  INVX4 U124 ( .A(n338), .Y(n339) );
  INVX2 U125 ( .A(n639), .Y(n640) );
  INVX2 U126 ( .A(n636), .Y(n637) );
  INVX2 U127 ( .A(n633), .Y(n634) );
  INVX1 U128 ( .A(n2323), .Y(n5) );
  INVX8 U129 ( .A(n2323), .Y(n6) );
  INVX8 U130 ( .A(n2332), .Y(n7) );
  INVX1 U131 ( .A(n272), .Y(n8) );
  AND2X2 U132 ( .A(n11), .B(n1608), .Y(\data_out<12> ) );
  AND2X2 U133 ( .A(n1609), .B(n11), .Y(\data_out<13> ) );
  INVX1 U134 ( .A(n272), .Y(n11) );
  INVX1 U135 ( .A(n1205), .Y(n12) );
  INVX1 U136 ( .A(n1205), .Y(n13) );
  INVX1 U137 ( .A(n274), .Y(n1203) );
  INVX1 U138 ( .A(n274), .Y(n14) );
  AND2X2 U139 ( .A(\mem<30><0> ), .B(n617), .Y(n15) );
  INVX1 U140 ( .A(n15), .Y(n16) );
  AND2X2 U141 ( .A(\mem<30><1> ), .B(n617), .Y(n17) );
  INVX1 U142 ( .A(n17), .Y(n18) );
  AND2X2 U143 ( .A(\mem<30><2> ), .B(n617), .Y(n19) );
  INVX1 U144 ( .A(n19), .Y(n20) );
  AND2X2 U145 ( .A(\mem<30><3> ), .B(n617), .Y(n21) );
  INVX1 U146 ( .A(n21), .Y(n22) );
  AND2X2 U147 ( .A(\mem<30><4> ), .B(n617), .Y(n23) );
  INVX1 U148 ( .A(n23), .Y(n24) );
  AND2X2 U149 ( .A(\mem<30><5> ), .B(n617), .Y(n25) );
  INVX1 U150 ( .A(n25), .Y(n26) );
  AND2X2 U151 ( .A(\mem<30><6> ), .B(n617), .Y(n27) );
  INVX1 U152 ( .A(n27), .Y(n28) );
  AND2X2 U153 ( .A(\mem<30><7> ), .B(n617), .Y(n29) );
  INVX1 U154 ( .A(n29), .Y(n30) );
  AND2X2 U155 ( .A(\mem<30><8> ), .B(n617), .Y(n31) );
  INVX1 U156 ( .A(n31), .Y(n32) );
  AND2X2 U157 ( .A(\mem<30><9> ), .B(n617), .Y(n33) );
  INVX1 U158 ( .A(n33), .Y(n34) );
  AND2X2 U159 ( .A(\mem<30><10> ), .B(n617), .Y(n35) );
  INVX1 U160 ( .A(n35), .Y(n36) );
  AND2X2 U161 ( .A(\mem<30><11> ), .B(n617), .Y(n37) );
  INVX1 U162 ( .A(n37), .Y(n38) );
  AND2X2 U163 ( .A(\mem<30><12> ), .B(n617), .Y(n39) );
  INVX1 U164 ( .A(n39), .Y(n40) );
  AND2X2 U165 ( .A(\mem<30><13> ), .B(n617), .Y(n41) );
  INVX1 U166 ( .A(n41), .Y(n42) );
  AND2X2 U167 ( .A(\mem<30><14> ), .B(n617), .Y(n43) );
  INVX1 U168 ( .A(n43), .Y(n44) );
  AND2X2 U169 ( .A(\mem<30><15> ), .B(n617), .Y(n45) );
  INVX1 U170 ( .A(n45), .Y(n46) );
  AND2X2 U171 ( .A(\mem<29><0> ), .B(n2242), .Y(n47) );
  INVX1 U172 ( .A(n47), .Y(n48) );
  AND2X2 U173 ( .A(\mem<29><1> ), .B(n2242), .Y(n49) );
  INVX1 U174 ( .A(n49), .Y(n50) );
  AND2X2 U175 ( .A(\mem<29><2> ), .B(n2242), .Y(n51) );
  INVX1 U176 ( .A(n51), .Y(n52) );
  AND2X2 U177 ( .A(\mem<29><3> ), .B(n2242), .Y(n53) );
  INVX1 U178 ( .A(n53), .Y(n54) );
  AND2X2 U179 ( .A(\mem<29><4> ), .B(n2242), .Y(n55) );
  INVX1 U180 ( .A(n55), .Y(n56) );
  AND2X2 U181 ( .A(\mem<29><5> ), .B(n2242), .Y(n57) );
  INVX1 U182 ( .A(n57), .Y(n58) );
  AND2X2 U183 ( .A(\mem<29><6> ), .B(n2242), .Y(n59) );
  INVX1 U184 ( .A(n59), .Y(n60) );
  AND2X2 U185 ( .A(\mem<29><7> ), .B(n2242), .Y(n61) );
  INVX1 U186 ( .A(n61), .Y(n62) );
  AND2X2 U187 ( .A(\mem<29><8> ), .B(n619), .Y(n63) );
  INVX1 U188 ( .A(n63), .Y(n64) );
  AND2X2 U189 ( .A(\mem<29><9> ), .B(n619), .Y(n65) );
  INVX1 U190 ( .A(n65), .Y(n66) );
  AND2X2 U191 ( .A(\mem<29><10> ), .B(n619), .Y(n67) );
  INVX1 U192 ( .A(n67), .Y(n68) );
  AND2X2 U193 ( .A(\mem<29><11> ), .B(n619), .Y(n69) );
  INVX1 U194 ( .A(n69), .Y(n70) );
  AND2X2 U195 ( .A(\mem<29><12> ), .B(n619), .Y(n71) );
  INVX1 U196 ( .A(n71), .Y(n72) );
  AND2X2 U197 ( .A(\mem<29><13> ), .B(n619), .Y(n73) );
  INVX1 U198 ( .A(n73), .Y(n74) );
  AND2X2 U199 ( .A(\mem<29><14> ), .B(n619), .Y(n75) );
  INVX1 U200 ( .A(n75), .Y(n76) );
  AND2X2 U201 ( .A(\mem<29><15> ), .B(n619), .Y(n77) );
  INVX1 U202 ( .A(n77), .Y(n78) );
  AND2X2 U203 ( .A(\mem<28><0> ), .B(n622), .Y(n79) );
  INVX1 U204 ( .A(n79), .Y(n80) );
  AND2X2 U205 ( .A(\mem<28><1> ), .B(n622), .Y(n81) );
  INVX1 U206 ( .A(n81), .Y(n82) );
  AND2X2 U207 ( .A(\mem<28><2> ), .B(n622), .Y(n83) );
  INVX1 U208 ( .A(n83), .Y(n84) );
  AND2X2 U209 ( .A(\mem<28><3> ), .B(n622), .Y(n85) );
  INVX1 U210 ( .A(n85), .Y(n86) );
  AND2X2 U211 ( .A(\mem<28><4> ), .B(n622), .Y(n87) );
  INVX1 U212 ( .A(n87), .Y(n88) );
  AND2X2 U213 ( .A(\mem<28><5> ), .B(n622), .Y(n89) );
  INVX1 U214 ( .A(n89), .Y(n90) );
  AND2X2 U215 ( .A(\mem<28><6> ), .B(n622), .Y(n91) );
  INVX1 U216 ( .A(n91), .Y(n92) );
  AND2X2 U217 ( .A(\mem<28><7> ), .B(n622), .Y(n93) );
  INVX1 U218 ( .A(n93), .Y(n94) );
  AND2X2 U219 ( .A(\mem<28><8> ), .B(n622), .Y(n95) );
  INVX1 U220 ( .A(n95), .Y(n96) );
  AND2X2 U221 ( .A(\mem<28><9> ), .B(n622), .Y(n97) );
  INVX1 U222 ( .A(n97), .Y(n98) );
  AND2X2 U223 ( .A(\mem<28><10> ), .B(n622), .Y(n99) );
  INVX1 U224 ( .A(n99), .Y(n100) );
  AND2X2 U225 ( .A(\mem<28><11> ), .B(n622), .Y(n101) );
  INVX1 U226 ( .A(n101), .Y(n102) );
  AND2X2 U227 ( .A(\mem<28><12> ), .B(n622), .Y(n103) );
  INVX1 U228 ( .A(n103), .Y(n104) );
  AND2X2 U229 ( .A(\mem<28><13> ), .B(n622), .Y(n105) );
  INVX1 U230 ( .A(n105), .Y(n106) );
  AND2X2 U231 ( .A(\mem<28><14> ), .B(n622), .Y(n107) );
  INVX1 U232 ( .A(n107), .Y(n108) );
  AND2X2 U233 ( .A(\mem<28><15> ), .B(n622), .Y(n109) );
  INVX1 U234 ( .A(n109), .Y(n110) );
  AND2X2 U235 ( .A(\mem<27><0> ), .B(n624), .Y(n111) );
  INVX1 U236 ( .A(n111), .Y(n112) );
  AND2X2 U237 ( .A(\mem<27><1> ), .B(n624), .Y(n113) );
  INVX1 U238 ( .A(n113), .Y(n114) );
  AND2X2 U239 ( .A(\mem<27><2> ), .B(n624), .Y(n115) );
  INVX1 U240 ( .A(n115), .Y(n116) );
  AND2X2 U241 ( .A(\mem<27><3> ), .B(n624), .Y(n117) );
  INVX1 U242 ( .A(n117), .Y(n118) );
  AND2X2 U243 ( .A(\mem<27><4> ), .B(n624), .Y(n119) );
  INVX1 U244 ( .A(n119), .Y(n120) );
  AND2X2 U245 ( .A(\mem<27><5> ), .B(n624), .Y(n121) );
  INVX1 U246 ( .A(n121), .Y(n122) );
  AND2X2 U247 ( .A(\mem<27><6> ), .B(n624), .Y(n123) );
  INVX1 U248 ( .A(n123), .Y(n124) );
  AND2X2 U249 ( .A(\mem<27><7> ), .B(n624), .Y(n125) );
  INVX1 U250 ( .A(n125), .Y(n126) );
  AND2X2 U251 ( .A(\mem<27><8> ), .B(n624), .Y(n127) );
  INVX1 U252 ( .A(n127), .Y(n128) );
  AND2X2 U253 ( .A(\mem<27><9> ), .B(n624), .Y(n129) );
  INVX1 U254 ( .A(n129), .Y(n130) );
  AND2X2 U255 ( .A(\mem<27><10> ), .B(n624), .Y(n131) );
  INVX1 U256 ( .A(n131), .Y(n132) );
  AND2X2 U257 ( .A(\mem<27><11> ), .B(n624), .Y(n133) );
  INVX1 U258 ( .A(n133), .Y(n134) );
  AND2X2 U259 ( .A(\mem<27><12> ), .B(n624), .Y(n135) );
  INVX1 U260 ( .A(n135), .Y(n136) );
  AND2X2 U261 ( .A(\mem<27><13> ), .B(n624), .Y(n137) );
  INVX1 U262 ( .A(n137), .Y(n138) );
  AND2X2 U263 ( .A(\mem<27><14> ), .B(n624), .Y(n139) );
  INVX1 U264 ( .A(n139), .Y(n140) );
  AND2X2 U265 ( .A(\mem<27><15> ), .B(n624), .Y(n141) );
  INVX1 U266 ( .A(n141), .Y(n142) );
  AND2X2 U267 ( .A(\mem<26><8> ), .B(n626), .Y(n143) );
  INVX1 U268 ( .A(n143), .Y(n144) );
  AND2X2 U269 ( .A(\mem<26><9> ), .B(n626), .Y(n145) );
  INVX1 U270 ( .A(n145), .Y(n146) );
  AND2X2 U271 ( .A(\mem<26><10> ), .B(n626), .Y(n147) );
  INVX1 U272 ( .A(n147), .Y(n148) );
  AND2X2 U273 ( .A(\mem<26><11> ), .B(n626), .Y(n149) );
  INVX1 U274 ( .A(n149), .Y(n150) );
  AND2X2 U275 ( .A(\mem<26><12> ), .B(n626), .Y(n151) );
  INVX1 U276 ( .A(n151), .Y(n152) );
  AND2X2 U277 ( .A(\mem<26><13> ), .B(n626), .Y(n153) );
  INVX1 U278 ( .A(n153), .Y(n154) );
  AND2X2 U279 ( .A(\mem<26><14> ), .B(n626), .Y(n155) );
  INVX1 U280 ( .A(n155), .Y(n156) );
  AND2X2 U281 ( .A(\mem<26><15> ), .B(n626), .Y(n157) );
  INVX1 U282 ( .A(n157), .Y(n158) );
  AND2X2 U283 ( .A(\mem<25><8> ), .B(n628), .Y(n159) );
  INVX1 U284 ( .A(n159), .Y(n160) );
  AND2X2 U285 ( .A(\mem<25><9> ), .B(n628), .Y(n161) );
  INVX1 U286 ( .A(n161), .Y(n162) );
  AND2X2 U287 ( .A(\mem<25><10> ), .B(n628), .Y(n163) );
  INVX1 U288 ( .A(n163), .Y(n164) );
  AND2X2 U289 ( .A(\mem<25><11> ), .B(n628), .Y(n165) );
  INVX1 U290 ( .A(n165), .Y(n166) );
  AND2X2 U291 ( .A(\mem<25><12> ), .B(n628), .Y(n167) );
  INVX1 U292 ( .A(n167), .Y(n168) );
  AND2X2 U293 ( .A(\mem<25><13> ), .B(n628), .Y(n169) );
  INVX1 U294 ( .A(n169), .Y(n170) );
  AND2X2 U295 ( .A(\mem<25><14> ), .B(n628), .Y(n171) );
  INVX1 U296 ( .A(n171), .Y(n172) );
  AND2X2 U297 ( .A(\mem<25><15> ), .B(n628), .Y(n173) );
  INVX1 U298 ( .A(n173), .Y(n174) );
  AND2X2 U299 ( .A(\mem<24><0> ), .B(n630), .Y(n175) );
  INVX1 U300 ( .A(n175), .Y(n176) );
  AND2X2 U301 ( .A(\mem<24><1> ), .B(n630), .Y(n177) );
  INVX1 U302 ( .A(n177), .Y(n178) );
  AND2X2 U303 ( .A(\mem<24><2> ), .B(n630), .Y(n179) );
  INVX1 U304 ( .A(n179), .Y(n180) );
  AND2X2 U305 ( .A(\mem<24><3> ), .B(n630), .Y(n181) );
  INVX1 U306 ( .A(n181), .Y(n182) );
  AND2X2 U307 ( .A(\mem<24><4> ), .B(n630), .Y(n183) );
  INVX1 U308 ( .A(n183), .Y(n184) );
  AND2X2 U309 ( .A(\mem<24><5> ), .B(n630), .Y(n185) );
  INVX1 U310 ( .A(n185), .Y(n186) );
  AND2X2 U311 ( .A(\mem<24><6> ), .B(n630), .Y(n187) );
  INVX1 U312 ( .A(n187), .Y(n188) );
  AND2X2 U313 ( .A(\mem<24><7> ), .B(n630), .Y(n189) );
  INVX1 U314 ( .A(n189), .Y(n190) );
  AND2X2 U315 ( .A(\mem<24><8> ), .B(n630), .Y(n191) );
  INVX1 U316 ( .A(n191), .Y(n192) );
  AND2X2 U317 ( .A(\mem<24><9> ), .B(n630), .Y(n193) );
  INVX1 U318 ( .A(n193), .Y(n194) );
  AND2X2 U319 ( .A(\mem<24><10> ), .B(n630), .Y(n195) );
  INVX1 U320 ( .A(n195), .Y(n196) );
  AND2X2 U321 ( .A(\mem<24><11> ), .B(n630), .Y(n197) );
  INVX1 U322 ( .A(n197), .Y(n198) );
  AND2X2 U323 ( .A(\mem<24><12> ), .B(n630), .Y(n199) );
  INVX1 U324 ( .A(n199), .Y(n200) );
  AND2X2 U325 ( .A(\mem<24><13> ), .B(n630), .Y(n201) );
  INVX1 U326 ( .A(n201), .Y(n202) );
  AND2X2 U327 ( .A(\mem<24><14> ), .B(n630), .Y(n203) );
  INVX1 U328 ( .A(n203), .Y(n204) );
  AND2X2 U329 ( .A(\mem<24><15> ), .B(n630), .Y(n205) );
  INVX1 U330 ( .A(n205), .Y(n206) );
  AND2X2 U331 ( .A(\mem<23><8> ), .B(n632), .Y(n207) );
  INVX1 U332 ( .A(n207), .Y(n208) );
  AND2X2 U333 ( .A(\mem<23><9> ), .B(n632), .Y(n209) );
  INVX1 U334 ( .A(n209), .Y(n210) );
  AND2X2 U335 ( .A(\mem<23><10> ), .B(n632), .Y(n211) );
  INVX1 U336 ( .A(n211), .Y(n212) );
  AND2X2 U337 ( .A(\mem<23><11> ), .B(n632), .Y(n213) );
  INVX1 U338 ( .A(n213), .Y(n215) );
  AND2X2 U339 ( .A(\mem<23><12> ), .B(n632), .Y(n216) );
  INVX1 U340 ( .A(n216), .Y(n217) );
  AND2X2 U341 ( .A(\mem<23><13> ), .B(n632), .Y(n218) );
  INVX1 U342 ( .A(n218), .Y(n219) );
  AND2X2 U343 ( .A(\mem<23><14> ), .B(n632), .Y(n220) );
  INVX1 U344 ( .A(n220), .Y(n221) );
  AND2X2 U345 ( .A(\mem<23><15> ), .B(n632), .Y(n222) );
  INVX1 U346 ( .A(n222), .Y(n223) );
  AND2X2 U347 ( .A(\mem<22><8> ), .B(n634), .Y(n224) );
  INVX1 U348 ( .A(n224), .Y(n225) );
  AND2X2 U349 ( .A(\mem<22><9> ), .B(n634), .Y(n226) );
  INVX1 U350 ( .A(n226), .Y(n227) );
  AND2X2 U351 ( .A(\mem<22><10> ), .B(n634), .Y(n228) );
  INVX1 U352 ( .A(n228), .Y(n229) );
  AND2X2 U353 ( .A(\mem<22><11> ), .B(n634), .Y(n230) );
  INVX1 U354 ( .A(n230), .Y(n231) );
  AND2X2 U355 ( .A(\mem<22><12> ), .B(n634), .Y(n232) );
  INVX1 U356 ( .A(n232), .Y(n233) );
  AND2X2 U357 ( .A(\mem<22><13> ), .B(n634), .Y(n234) );
  INVX1 U358 ( .A(n234), .Y(n235) );
  AND2X2 U359 ( .A(\mem<22><14> ), .B(n634), .Y(n236) );
  INVX1 U360 ( .A(n236), .Y(n237) );
  AND2X2 U361 ( .A(\mem<22><15> ), .B(n634), .Y(n238) );
  INVX1 U362 ( .A(n238), .Y(n239) );
  AND2X2 U363 ( .A(\mem<21><8> ), .B(n637), .Y(n240) );
  INVX1 U364 ( .A(n240), .Y(n241) );
  AND2X2 U365 ( .A(\mem<21><9> ), .B(n637), .Y(n242) );
  INVX1 U366 ( .A(n242), .Y(n243) );
  AND2X2 U367 ( .A(\mem<21><10> ), .B(n637), .Y(n244) );
  INVX1 U368 ( .A(n244), .Y(n245) );
  AND2X2 U369 ( .A(\mem<21><11> ), .B(n637), .Y(n246) );
  INVX1 U370 ( .A(n246), .Y(n247) );
  AND2X2 U371 ( .A(\mem<21><12> ), .B(n637), .Y(n248) );
  INVX1 U372 ( .A(n248), .Y(n249) );
  AND2X2 U373 ( .A(\mem<21><13> ), .B(n637), .Y(n250) );
  INVX1 U374 ( .A(n250), .Y(n251) );
  AND2X2 U375 ( .A(\mem<21><14> ), .B(n637), .Y(n252) );
  INVX1 U376 ( .A(n252), .Y(n253) );
  AND2X2 U377 ( .A(\mem<21><15> ), .B(n637), .Y(n254) );
  INVX1 U378 ( .A(n254), .Y(n255) );
  AND2X2 U379 ( .A(\mem<20><8> ), .B(n640), .Y(n256) );
  INVX1 U380 ( .A(n256), .Y(n257) );
  AND2X2 U381 ( .A(\mem<20><9> ), .B(n640), .Y(n258) );
  INVX1 U382 ( .A(n258), .Y(n259) );
  AND2X2 U383 ( .A(\mem<20><10> ), .B(n640), .Y(n260) );
  INVX1 U384 ( .A(n260), .Y(n261) );
  AND2X2 U385 ( .A(\mem<20><11> ), .B(n640), .Y(n262) );
  INVX1 U386 ( .A(n262), .Y(n263) );
  AND2X2 U387 ( .A(\mem<20><12> ), .B(n640), .Y(n264) );
  INVX1 U388 ( .A(n264), .Y(n265) );
  AND2X2 U389 ( .A(\mem<20><13> ), .B(n640), .Y(n266) );
  INVX1 U390 ( .A(n266), .Y(n267) );
  AND2X2 U391 ( .A(\mem<20><14> ), .B(n640), .Y(n268) );
  INVX1 U392 ( .A(n268), .Y(n269) );
  AND2X2 U393 ( .A(\mem<20><15> ), .B(n640), .Y(n270) );
  INVX1 U394 ( .A(n270), .Y(n271) );
  INVX1 U395 ( .A(n2), .Y(n272) );
  INVX1 U396 ( .A(write), .Y(n1205) );
  INVX1 U397 ( .A(n1205), .Y(n273) );
  AND2X2 U398 ( .A(n1195), .B(n1651), .Y(n275) );
  AND2X2 U399 ( .A(n1173), .B(n1653), .Y(n277) );
  INVX1 U400 ( .A(n318), .Y(n279) );
  INVX4 U401 ( .A(n320), .Y(n321) );
  INVX4 U402 ( .A(n322), .Y(n323) );
  INVX4 U403 ( .A(n324), .Y(n325) );
  INVX4 U404 ( .A(n326), .Y(n327) );
  INVX4 U405 ( .A(n328), .Y(n329) );
  INVX4 U406 ( .A(n330), .Y(n331) );
  INVX4 U407 ( .A(n332), .Y(n333) );
  INVX4 U408 ( .A(n334), .Y(n335) );
  AND2X2 U409 ( .A(n1173), .B(n1627), .Y(n280) );
  INVX4 U410 ( .A(n336), .Y(n337) );
  AND2X2 U411 ( .A(n1197), .B(n1673), .Y(n282) );
  AND2X2 U412 ( .A(n1198), .B(n1675), .Y(n284) );
  INVX4 U413 ( .A(n342), .Y(n343) );
  INVX4 U414 ( .A(n344), .Y(n345) );
  INVX4 U415 ( .A(n346), .Y(n347) );
  INVX4 U416 ( .A(n348), .Y(n349) );
  INVX4 U417 ( .A(n350), .Y(n351) );
  OR2X2 U418 ( .A(n1585), .B(n12), .Y(n286) );
  INVX1 U419 ( .A(n286), .Y(\data_out<0> ) );
  OR2X2 U420 ( .A(n1), .B(n1587), .Y(n288) );
  INVX1 U421 ( .A(n288), .Y(\data_out<1> ) );
  OR2X2 U422 ( .A(n273), .B(n1589), .Y(n290) );
  INVX1 U423 ( .A(n290), .Y(\data_out<2> ) );
  OR2X2 U424 ( .A(n13), .B(n1591), .Y(n292) );
  INVX1 U425 ( .A(n292), .Y(\data_out<3> ) );
  OR2X2 U426 ( .A(n273), .B(n1593), .Y(n294) );
  INVX1 U427 ( .A(n294), .Y(\data_out<4> ) );
  OR2X2 U428 ( .A(n14), .B(n1595), .Y(n296) );
  INVX1 U429 ( .A(n296), .Y(\data_out<5> ) );
  OR2X2 U430 ( .A(n1203), .B(n1597), .Y(n298) );
  INVX1 U431 ( .A(n298), .Y(\data_out<6> ) );
  OR2X2 U432 ( .A(n13), .B(n1599), .Y(n300) );
  INVX1 U433 ( .A(n300), .Y(\data_out<7> ) );
  OR2X2 U434 ( .A(n14), .B(n1601), .Y(n302) );
  INVX1 U435 ( .A(n302), .Y(\data_out<8> ) );
  OR2X2 U436 ( .A(n1603), .B(n12), .Y(n304) );
  INVX1 U437 ( .A(n304), .Y(\data_out<9> ) );
  OR2X2 U438 ( .A(n1203), .B(n1605), .Y(n306) );
  INVX1 U439 ( .A(n306), .Y(\data_out<10> ) );
  OR2X2 U440 ( .A(n1), .B(n1607), .Y(n308) );
  INVX1 U441 ( .A(n308), .Y(\data_out<11> ) );
  OR2X2 U442 ( .A(n1204), .B(n1611), .Y(n310) );
  INVX1 U443 ( .A(n310), .Y(\data_out<14> ) );
  OR2X2 U444 ( .A(n1204), .B(n1613), .Y(n312) );
  INVX1 U445 ( .A(n312), .Y(\data_out<15> ) );
  AND2X2 U446 ( .A(n1194), .B(n1629), .Y(n314) );
  AND2X2 U447 ( .A(n1191), .B(n1653), .Y(n316) );
  AND2X2 U448 ( .A(n1192), .B(n1655), .Y(n318) );
  INVX1 U449 ( .A(n318), .Y(n319) );
  AND2X2 U450 ( .A(n1193), .B(n1626), .Y(n320) );
  AND2X2 U451 ( .A(n1190), .B(n1657), .Y(n322) );
  AND2X2 U452 ( .A(n1191), .B(n1659), .Y(n324) );
  AND2X2 U453 ( .A(n1189), .B(n1661), .Y(n326) );
  AND2X2 U454 ( .A(n1189), .B(n1663), .Y(n328) );
  AND2X2 U455 ( .A(n1189), .B(n1665), .Y(n330) );
  AND2X2 U456 ( .A(n1190), .B(n1667), .Y(n332) );
  AND2X2 U457 ( .A(n1172), .B(n1669), .Y(n334) );
  AND2X2 U458 ( .A(n1195), .B(n1671), .Y(n336) );
  AND2X2 U459 ( .A(n1194), .B(n1673), .Y(n338) );
  AND2X2 U460 ( .A(n1178), .B(n1675), .Y(n340) );
  AND2X2 U461 ( .A(n1201), .B(n1677), .Y(n342) );
  AND2X2 U462 ( .A(n1202), .B(n1679), .Y(n344) );
  AND2X2 U463 ( .A(n1201), .B(n1681), .Y(n346) );
  AND2X2 U464 ( .A(n1202), .B(n1683), .Y(n348) );
  AND2X2 U465 ( .A(n1192), .B(n1628), .Y(n350) );
  AND2X2 U466 ( .A(\mem<19><0> ), .B(n276), .Y(n352) );
  INVX1 U467 ( .A(n352), .Y(n353) );
  AND2X2 U468 ( .A(\mem<19><1> ), .B(n276), .Y(n354) );
  INVX1 U469 ( .A(n354), .Y(n355) );
  AND2X2 U470 ( .A(\mem<19><2> ), .B(n276), .Y(n356) );
  INVX1 U471 ( .A(n356), .Y(n357) );
  AND2X2 U472 ( .A(\mem<19><3> ), .B(n276), .Y(n358) );
  INVX1 U473 ( .A(n358), .Y(n359) );
  AND2X2 U474 ( .A(\mem<19><4> ), .B(n276), .Y(n360) );
  INVX1 U475 ( .A(n360), .Y(n361) );
  AND2X2 U476 ( .A(\mem<19><5> ), .B(n276), .Y(n362) );
  INVX1 U477 ( .A(n362), .Y(n363) );
  AND2X2 U478 ( .A(\mem<19><6> ), .B(n276), .Y(n364) );
  INVX1 U479 ( .A(n364), .Y(n365) );
  AND2X2 U480 ( .A(\mem<19><7> ), .B(n276), .Y(n366) );
  INVX1 U481 ( .A(n366), .Y(n367) );
  AND2X2 U482 ( .A(\mem<19><8> ), .B(n276), .Y(n368) );
  INVX1 U483 ( .A(n368), .Y(n369) );
  AND2X2 U484 ( .A(\mem<19><9> ), .B(n276), .Y(n370) );
  INVX1 U485 ( .A(n370), .Y(n371) );
  AND2X2 U486 ( .A(\mem<19><10> ), .B(n276), .Y(n372) );
  INVX1 U487 ( .A(n372), .Y(n373) );
  AND2X2 U488 ( .A(\mem<18><0> ), .B(n317), .Y(n374) );
  INVX1 U489 ( .A(n374), .Y(n375) );
  AND2X2 U490 ( .A(\mem<18><1> ), .B(n317), .Y(n376) );
  INVX1 U491 ( .A(n376), .Y(n377) );
  AND2X2 U492 ( .A(\mem<18><2> ), .B(n317), .Y(n378) );
  INVX1 U493 ( .A(n378), .Y(n379) );
  AND2X2 U494 ( .A(\mem<18><3> ), .B(n317), .Y(n380) );
  INVX1 U495 ( .A(n380), .Y(n381) );
  AND2X2 U496 ( .A(\mem<18><4> ), .B(n317), .Y(n382) );
  INVX1 U497 ( .A(n382), .Y(n383) );
  AND2X2 U498 ( .A(\mem<18><5> ), .B(n317), .Y(n384) );
  INVX1 U499 ( .A(n384), .Y(n385) );
  AND2X2 U500 ( .A(\mem<18><6> ), .B(n317), .Y(n386) );
  INVX1 U501 ( .A(n386), .Y(n387) );
  AND2X2 U502 ( .A(\mem<18><7> ), .B(n317), .Y(n388) );
  INVX1 U503 ( .A(n388), .Y(n389) );
  AND2X2 U504 ( .A(\mem<18><8> ), .B(n278), .Y(n390) );
  INVX1 U505 ( .A(n390), .Y(n391) );
  AND2X2 U506 ( .A(\mem<18><9> ), .B(n278), .Y(n392) );
  INVX1 U507 ( .A(n392), .Y(n393) );
  AND2X2 U508 ( .A(\mem<18><10> ), .B(n317), .Y(n394) );
  INVX1 U509 ( .A(n394), .Y(n395) );
  AND2X2 U510 ( .A(\mem<17><0> ), .B(n319), .Y(n396) );
  INVX1 U511 ( .A(n396), .Y(n397) );
  AND2X2 U512 ( .A(\mem<17><1> ), .B(n319), .Y(n398) );
  INVX1 U513 ( .A(n398), .Y(n399) );
  AND2X2 U514 ( .A(\mem<17><2> ), .B(n319), .Y(n400) );
  INVX1 U515 ( .A(n400), .Y(n401) );
  AND2X2 U516 ( .A(\mem<17><3> ), .B(n319), .Y(n402) );
  INVX1 U517 ( .A(n402), .Y(n403) );
  AND2X2 U518 ( .A(\mem<17><4> ), .B(n319), .Y(n404) );
  INVX1 U519 ( .A(n404), .Y(n405) );
  AND2X2 U520 ( .A(\mem<17><5> ), .B(n319), .Y(n406) );
  INVX1 U521 ( .A(n406), .Y(n407) );
  AND2X2 U522 ( .A(\mem<17><6> ), .B(n319), .Y(n408) );
  INVX1 U523 ( .A(n408), .Y(n409) );
  AND2X2 U524 ( .A(\mem<17><7> ), .B(n319), .Y(n410) );
  INVX1 U525 ( .A(n410), .Y(n411) );
  AND2X2 U526 ( .A(\mem<17><8> ), .B(n2266), .Y(n412) );
  INVX1 U527 ( .A(n412), .Y(n413) );
  AND2X2 U528 ( .A(\mem<17><9> ), .B(n2266), .Y(n414) );
  INVX1 U529 ( .A(n414), .Y(n415) );
  AND2X2 U530 ( .A(\mem<17><10> ), .B(n3), .Y(n416) );
  INVX1 U531 ( .A(n416), .Y(n417) );
  AND2X2 U532 ( .A(\mem<16><0> ), .B(n321), .Y(n418) );
  INVX1 U533 ( .A(n418), .Y(n419) );
  AND2X2 U534 ( .A(\mem<16><1> ), .B(n321), .Y(n420) );
  INVX1 U535 ( .A(n420), .Y(n421) );
  AND2X2 U536 ( .A(\mem<16><2> ), .B(n321), .Y(n422) );
  INVX1 U537 ( .A(n422), .Y(n423) );
  AND2X2 U538 ( .A(\mem<16><3> ), .B(n321), .Y(n424) );
  INVX1 U539 ( .A(n424), .Y(n425) );
  AND2X2 U540 ( .A(\mem<16><4> ), .B(n321), .Y(n426) );
  INVX1 U541 ( .A(n426), .Y(n427) );
  AND2X2 U542 ( .A(\mem<16><5> ), .B(n321), .Y(n428) );
  INVX1 U543 ( .A(n428), .Y(n429) );
  AND2X2 U544 ( .A(\mem<16><6> ), .B(n321), .Y(n430) );
  INVX1 U545 ( .A(n430), .Y(n431) );
  AND2X2 U546 ( .A(\mem<16><7> ), .B(n321), .Y(n432) );
  INVX1 U547 ( .A(n432), .Y(n433) );
  AND2X2 U548 ( .A(\mem<16><8> ), .B(n321), .Y(n434) );
  INVX1 U549 ( .A(n434), .Y(n435) );
  AND2X2 U550 ( .A(\mem<16><9> ), .B(n321), .Y(n436) );
  INVX1 U551 ( .A(n436), .Y(n437) );
  AND2X2 U552 ( .A(\mem<16><10> ), .B(n321), .Y(n438) );
  INVX1 U553 ( .A(n438), .Y(n439) );
  AND2X2 U554 ( .A(\mem<15><0> ), .B(n323), .Y(n440) );
  INVX1 U555 ( .A(n440), .Y(n441) );
  AND2X2 U556 ( .A(\mem<15><1> ), .B(n323), .Y(n442) );
  INVX1 U557 ( .A(n442), .Y(n443) );
  AND2X2 U558 ( .A(\mem<15><2> ), .B(n323), .Y(n444) );
  INVX1 U559 ( .A(n444), .Y(n445) );
  AND2X2 U560 ( .A(\mem<15><3> ), .B(n323), .Y(n446) );
  INVX1 U561 ( .A(n446), .Y(n447) );
  AND2X2 U562 ( .A(\mem<15><4> ), .B(n323), .Y(n448) );
  INVX1 U563 ( .A(n448), .Y(n449) );
  AND2X2 U564 ( .A(\mem<15><5> ), .B(n323), .Y(n450) );
  INVX1 U565 ( .A(n450), .Y(n451) );
  AND2X2 U566 ( .A(\mem<15><6> ), .B(n323), .Y(n452) );
  INVX1 U567 ( .A(n452), .Y(n453) );
  AND2X2 U568 ( .A(\mem<15><7> ), .B(n323), .Y(n454) );
  INVX1 U569 ( .A(n454), .Y(n455) );
  AND2X2 U570 ( .A(\mem<15><8> ), .B(n323), .Y(n456) );
  INVX1 U571 ( .A(n456), .Y(n457) );
  AND2X2 U572 ( .A(\mem<15><9> ), .B(n323), .Y(n458) );
  INVX1 U573 ( .A(n458), .Y(n459) );
  AND2X2 U574 ( .A(\mem<15><10> ), .B(n323), .Y(n460) );
  INVX1 U575 ( .A(n460), .Y(n461) );
  AND2X2 U576 ( .A(\mem<14><0> ), .B(n325), .Y(n462) );
  INVX1 U577 ( .A(n462), .Y(n463) );
  AND2X2 U578 ( .A(\mem<14><1> ), .B(n325), .Y(n464) );
  INVX1 U579 ( .A(n464), .Y(n465) );
  AND2X2 U580 ( .A(\mem<14><2> ), .B(n325), .Y(n466) );
  INVX1 U581 ( .A(n466), .Y(n467) );
  AND2X2 U582 ( .A(\mem<14><3> ), .B(n325), .Y(n468) );
  INVX1 U583 ( .A(n468), .Y(n469) );
  AND2X2 U584 ( .A(\mem<14><4> ), .B(n325), .Y(n470) );
  INVX1 U585 ( .A(n470), .Y(n471) );
  AND2X2 U586 ( .A(\mem<14><5> ), .B(n325), .Y(n472) );
  INVX1 U587 ( .A(n472), .Y(n473) );
  AND2X2 U588 ( .A(\mem<14><6> ), .B(n325), .Y(n474) );
  INVX1 U589 ( .A(n474), .Y(n475) );
  AND2X2 U590 ( .A(\mem<14><7> ), .B(n325), .Y(n476) );
  INVX1 U591 ( .A(n476), .Y(n477) );
  AND2X2 U592 ( .A(\mem<14><8> ), .B(n325), .Y(n478) );
  INVX1 U593 ( .A(n478), .Y(n479) );
  AND2X2 U594 ( .A(\mem<14><9> ), .B(n325), .Y(n480) );
  INVX1 U595 ( .A(n480), .Y(n481) );
  AND2X2 U596 ( .A(\mem<14><10> ), .B(n325), .Y(n482) );
  INVX1 U597 ( .A(n482), .Y(n483) );
  AND2X2 U598 ( .A(\mem<13><0> ), .B(n327), .Y(n484) );
  INVX1 U599 ( .A(n484), .Y(n485) );
  AND2X2 U600 ( .A(\mem<13><1> ), .B(n327), .Y(n486) );
  INVX1 U601 ( .A(n486), .Y(n487) );
  AND2X2 U602 ( .A(\mem<13><2> ), .B(n327), .Y(n488) );
  INVX1 U603 ( .A(n488), .Y(n489) );
  AND2X2 U604 ( .A(\mem<13><3> ), .B(n327), .Y(n490) );
  INVX1 U605 ( .A(n490), .Y(n491) );
  AND2X2 U606 ( .A(\mem<13><4> ), .B(n327), .Y(n492) );
  INVX1 U607 ( .A(n492), .Y(n493) );
  AND2X2 U608 ( .A(\mem<13><5> ), .B(n327), .Y(n494) );
  INVX1 U609 ( .A(n494), .Y(n495) );
  AND2X2 U610 ( .A(\mem<13><6> ), .B(n327), .Y(n496) );
  INVX1 U611 ( .A(n496), .Y(n497) );
  AND2X2 U612 ( .A(\mem<13><7> ), .B(n327), .Y(n498) );
  INVX1 U613 ( .A(n498), .Y(n499) );
  AND2X2 U614 ( .A(\mem<13><8> ), .B(n327), .Y(n500) );
  INVX1 U615 ( .A(n500), .Y(n501) );
  AND2X2 U616 ( .A(\mem<13><9> ), .B(n327), .Y(n502) );
  INVX1 U617 ( .A(n502), .Y(n503) );
  AND2X2 U618 ( .A(\mem<13><10> ), .B(n327), .Y(n504) );
  INVX1 U619 ( .A(n504), .Y(n505) );
  AND2X2 U620 ( .A(\mem<12><0> ), .B(n329), .Y(n506) );
  INVX1 U621 ( .A(n506), .Y(n507) );
  AND2X2 U622 ( .A(\mem<12><1> ), .B(n329), .Y(n508) );
  INVX1 U623 ( .A(n508), .Y(n509) );
  AND2X2 U624 ( .A(\mem<12><2> ), .B(n329), .Y(n510) );
  INVX1 U625 ( .A(n510), .Y(n511) );
  AND2X2 U626 ( .A(\mem<12><3> ), .B(n329), .Y(n512) );
  INVX1 U627 ( .A(n512), .Y(n513) );
  AND2X2 U628 ( .A(\mem<12><4> ), .B(n329), .Y(n514) );
  INVX1 U629 ( .A(n514), .Y(n515) );
  AND2X2 U630 ( .A(\mem<12><5> ), .B(n329), .Y(n516) );
  INVX1 U631 ( .A(n516), .Y(n517) );
  AND2X2 U632 ( .A(\mem<12><6> ), .B(n329), .Y(n518) );
  INVX1 U633 ( .A(n518), .Y(n519) );
  AND2X2 U634 ( .A(\mem<12><7> ), .B(n329), .Y(n520) );
  INVX1 U635 ( .A(n520), .Y(n521) );
  AND2X2 U636 ( .A(\mem<12><8> ), .B(n329), .Y(n522) );
  INVX1 U637 ( .A(n522), .Y(n523) );
  AND2X2 U638 ( .A(\mem<12><9> ), .B(n329), .Y(n524) );
  INVX1 U639 ( .A(n524), .Y(n525) );
  AND2X2 U640 ( .A(\mem<12><10> ), .B(n329), .Y(n526) );
  INVX1 U641 ( .A(n526), .Y(n527) );
  AND2X2 U642 ( .A(\mem<11><0> ), .B(n331), .Y(n528) );
  INVX1 U643 ( .A(n528), .Y(n529) );
  AND2X2 U644 ( .A(\mem<11><1> ), .B(n331), .Y(n530) );
  INVX1 U645 ( .A(n530), .Y(n531) );
  AND2X2 U646 ( .A(\mem<11><2> ), .B(n331), .Y(n532) );
  INVX1 U647 ( .A(n532), .Y(n533) );
  AND2X2 U648 ( .A(\mem<11><3> ), .B(n331), .Y(n534) );
  INVX1 U649 ( .A(n534), .Y(n535) );
  AND2X2 U650 ( .A(\mem<11><4> ), .B(n331), .Y(n536) );
  INVX1 U651 ( .A(n536), .Y(n537) );
  AND2X2 U652 ( .A(\mem<11><5> ), .B(n331), .Y(n538) );
  INVX1 U653 ( .A(n538), .Y(n539) );
  AND2X2 U654 ( .A(\mem<11><6> ), .B(n331), .Y(n540) );
  INVX1 U655 ( .A(n540), .Y(n541) );
  AND2X2 U656 ( .A(\mem<11><7> ), .B(n331), .Y(n542) );
  INVX1 U657 ( .A(n542), .Y(n543) );
  AND2X2 U658 ( .A(\mem<11><8> ), .B(n331), .Y(n544) );
  INVX1 U659 ( .A(n544), .Y(n545) );
  AND2X2 U660 ( .A(\mem<11><9> ), .B(n331), .Y(n546) );
  INVX1 U661 ( .A(n546), .Y(n547) );
  AND2X2 U662 ( .A(\mem<11><10> ), .B(n331), .Y(n548) );
  INVX1 U663 ( .A(n548), .Y(n549) );
  AND2X2 U664 ( .A(\mem<10><0> ), .B(n333), .Y(n550) );
  INVX1 U665 ( .A(n550), .Y(n551) );
  AND2X2 U666 ( .A(\mem<10><1> ), .B(n333), .Y(n552) );
  INVX1 U667 ( .A(n552), .Y(n553) );
  AND2X2 U668 ( .A(\mem<10><2> ), .B(n333), .Y(n554) );
  INVX1 U669 ( .A(n554), .Y(n555) );
  AND2X2 U670 ( .A(\mem<10><3> ), .B(n333), .Y(n556) );
  INVX1 U671 ( .A(n556), .Y(n557) );
  AND2X2 U672 ( .A(\mem<10><4> ), .B(n333), .Y(n558) );
  INVX1 U673 ( .A(n558), .Y(n559) );
  AND2X2 U674 ( .A(\mem<10><5> ), .B(n333), .Y(n560) );
  INVX1 U675 ( .A(n560), .Y(n561) );
  AND2X2 U676 ( .A(\mem<10><6> ), .B(n333), .Y(n562) );
  INVX1 U677 ( .A(n562), .Y(n563) );
  AND2X2 U678 ( .A(\mem<10><7> ), .B(n333), .Y(n564) );
  INVX1 U679 ( .A(n564), .Y(n565) );
  AND2X2 U680 ( .A(\mem<10><8> ), .B(n333), .Y(n566) );
  INVX1 U681 ( .A(n566), .Y(n567) );
  AND2X2 U682 ( .A(\mem<10><9> ), .B(n333), .Y(n568) );
  INVX1 U683 ( .A(n568), .Y(n569) );
  AND2X2 U684 ( .A(\mem<10><10> ), .B(n333), .Y(n570) );
  INVX1 U685 ( .A(n570), .Y(n571) );
  AND2X2 U686 ( .A(\mem<9><0> ), .B(n335), .Y(n572) );
  INVX1 U687 ( .A(n572), .Y(n573) );
  AND2X2 U688 ( .A(\mem<9><1> ), .B(n335), .Y(n574) );
  INVX1 U689 ( .A(n574), .Y(n575) );
  AND2X2 U690 ( .A(\mem<9><2> ), .B(n335), .Y(n576) );
  INVX1 U691 ( .A(n576), .Y(n577) );
  AND2X2 U692 ( .A(\mem<9><3> ), .B(n335), .Y(n578) );
  INVX1 U693 ( .A(n578), .Y(n579) );
  AND2X2 U694 ( .A(\mem<9><4> ), .B(n335), .Y(n580) );
  INVX1 U695 ( .A(n580), .Y(n581) );
  AND2X2 U696 ( .A(\mem<9><5> ), .B(n335), .Y(n582) );
  INVX1 U697 ( .A(n582), .Y(n583) );
  AND2X2 U698 ( .A(\mem<9><6> ), .B(n335), .Y(n584) );
  INVX1 U699 ( .A(n584), .Y(n585) );
  AND2X2 U700 ( .A(\mem<9><7> ), .B(n335), .Y(n586) );
  INVX1 U701 ( .A(n586), .Y(n587) );
  AND2X2 U702 ( .A(\mem<9><8> ), .B(n335), .Y(n588) );
  INVX1 U703 ( .A(n588), .Y(n589) );
  AND2X2 U704 ( .A(\mem<9><9> ), .B(n335), .Y(n590) );
  INVX1 U705 ( .A(n590), .Y(n591) );
  AND2X2 U706 ( .A(\mem<9><10> ), .B(n335), .Y(n592) );
  INVX1 U707 ( .A(n592), .Y(n593) );
  AND2X2 U708 ( .A(\mem<0><0> ), .B(n351), .Y(n594) );
  INVX1 U709 ( .A(n594), .Y(n595) );
  AND2X2 U710 ( .A(\mem<0><1> ), .B(n351), .Y(n596) );
  INVX1 U711 ( .A(n596), .Y(n597) );
  AND2X2 U712 ( .A(\mem<0><2> ), .B(n351), .Y(n598) );
  INVX1 U713 ( .A(n598), .Y(n599) );
  AND2X2 U714 ( .A(\mem<0><3> ), .B(n351), .Y(n600) );
  INVX1 U715 ( .A(n600), .Y(n601) );
  AND2X2 U716 ( .A(\mem<0><4> ), .B(n351), .Y(n602) );
  INVX1 U717 ( .A(n602), .Y(n603) );
  AND2X2 U718 ( .A(\mem<0><5> ), .B(n351), .Y(n604) );
  INVX1 U719 ( .A(n604), .Y(n605) );
  AND2X2 U720 ( .A(\mem<0><6> ), .B(n351), .Y(n606) );
  INVX1 U721 ( .A(n606), .Y(n607) );
  AND2X2 U722 ( .A(\mem<0><7> ), .B(n351), .Y(n608) );
  INVX1 U723 ( .A(n608), .Y(n609) );
  AND2X2 U724 ( .A(\mem<0><8> ), .B(n351), .Y(n610) );
  INVX1 U725 ( .A(n610), .Y(n611) );
  AND2X2 U726 ( .A(\mem<0><9> ), .B(n351), .Y(n612) );
  INVX1 U727 ( .A(n612), .Y(n613) );
  AND2X2 U728 ( .A(\mem<0><10> ), .B(n351), .Y(n614) );
  INVX1 U729 ( .A(n614), .Y(n615) );
  AND2X2 U730 ( .A(n1195), .B(n1631), .Y(n616) );
  AND2X2 U731 ( .A(n1180), .B(n1633), .Y(n618) );
  INVX1 U732 ( .A(n618), .Y(n619) );
  INVX1 U733 ( .A(n618), .Y(n620) );
  AND2X2 U734 ( .A(n1179), .B(n1635), .Y(n621) );
  AND2X2 U735 ( .A(n1178), .B(n1637), .Y(n623) );
  AND2X2 U736 ( .A(n1178), .B(n1639), .Y(n625) );
  AND2X2 U737 ( .A(n1179), .B(n1641), .Y(n627) );
  AND2X2 U738 ( .A(n1181), .B(n1625), .Y(n629) );
  AND2X2 U739 ( .A(n1194), .B(n1643), .Y(n631) );
  AND2X2 U740 ( .A(n1181), .B(n1645), .Y(n633) );
  AND2X2 U741 ( .A(n1193), .B(n1647), .Y(n636) );
  AND2X2 U742 ( .A(n1193), .B(n1649), .Y(n639) );
  AND2X2 U743 ( .A(\data_in<0> ), .B(n1185), .Y(n642) );
  AND2X2 U744 ( .A(n1187), .B(\data_in<1> ), .Y(n643) );
  AND2X2 U745 ( .A(n1187), .B(\data_in<2> ), .Y(n644) );
  AND2X2 U746 ( .A(n1192), .B(\data_in<3> ), .Y(n645) );
  AND2X2 U747 ( .A(\data_in<4> ), .B(n2423), .Y(n646) );
  AND2X2 U748 ( .A(n1188), .B(\data_in<5> ), .Y(n647) );
  AND2X2 U749 ( .A(n1188), .B(\data_in<6> ), .Y(n648) );
  AND2X2 U750 ( .A(\data_in<7> ), .B(n1184), .Y(n649) );
  AND2X2 U751 ( .A(\data_in<8> ), .B(n2423), .Y(n650) );
  AND2X2 U752 ( .A(n1186), .B(\data_in<9> ), .Y(n1163) );
  AND2X2 U753 ( .A(n1186), .B(\data_in<10> ), .Y(n1164) );
  AND2X2 U754 ( .A(\data_in<11> ), .B(n1182), .Y(n1165) );
  INVX1 U755 ( .A(n1165), .Y(n1166) );
  AND2X2 U756 ( .A(\data_in<12> ), .B(n1183), .Y(n1167) );
  AND2X2 U757 ( .A(\data_in<13> ), .B(n1183), .Y(n1168) );
  AND2X2 U758 ( .A(\data_in<14> ), .B(n1184), .Y(n1169) );
  AND2X2 U759 ( .A(\data_in<15> ), .B(n1182), .Y(n1170) );
  INVX1 U760 ( .A(n1170), .Y(n1171) );
  INVX1 U761 ( .A(n2298), .Y(n1172) );
  INVX1 U762 ( .A(n2298), .Y(n1173) );
  BUFX2 U763 ( .A(n2343), .Y(n1174) );
  BUFX2 U764 ( .A(n2343), .Y(n1175) );
  BUFX2 U765 ( .A(n2343), .Y(n1176) );
  BUFX2 U766 ( .A(n2343), .Y(n1177) );
  INVX1 U767 ( .A(n1174), .Y(n1178) );
  INVX1 U768 ( .A(n1174), .Y(n1179) );
  INVX1 U769 ( .A(n1174), .Y(n1180) );
  INVX1 U770 ( .A(n1174), .Y(n1181) );
  INVX1 U771 ( .A(n1175), .Y(n1182) );
  INVX1 U772 ( .A(n1175), .Y(n1183) );
  INVX1 U773 ( .A(n1175), .Y(n1184) );
  INVX1 U774 ( .A(n1176), .Y(n1185) );
  INVX1 U775 ( .A(n1176), .Y(n1186) );
  INVX1 U776 ( .A(n1177), .Y(n1187) );
  INVX1 U777 ( .A(n1177), .Y(n1188) );
  INVX1 U778 ( .A(n1177), .Y(n1189) );
  INVX1 U779 ( .A(n1200), .Y(n1190) );
  INVX1 U780 ( .A(n1200), .Y(n1191) );
  INVX1 U781 ( .A(n1176), .Y(n1192) );
  INVX1 U782 ( .A(n1177), .Y(n1193) );
  INVX1 U783 ( .A(n1174), .Y(n1194) );
  INVX1 U784 ( .A(n1174), .Y(n1195) );
  INVX1 U785 ( .A(n1172), .Y(n1196) );
  INVX1 U786 ( .A(n1196), .Y(n1197) );
  INVX1 U787 ( .A(n1196), .Y(n1198) );
  INVX1 U788 ( .A(n1172), .Y(n1199) );
  INVX1 U789 ( .A(n1173), .Y(n1200) );
  INVX1 U790 ( .A(n1199), .Y(n1201) );
  INVX1 U791 ( .A(n1199), .Y(n1202) );
  INVX1 U792 ( .A(n2343), .Y(n2423) );
  INVX1 U793 ( .A(n2), .Y(n1204) );
  OR2X2 U794 ( .A(n8), .B(rst), .Y(n2343) );
  AND2X2 U795 ( .A(\mem<19><11> ), .B(n276), .Y(n1206) );
  INVX1 U796 ( .A(n1206), .Y(n1207) );
  AND2X2 U797 ( .A(\mem<19><12> ), .B(n276), .Y(n1208) );
  INVX1 U798 ( .A(n1208), .Y(n1209) );
  AND2X2 U799 ( .A(\mem<19><13> ), .B(n276), .Y(n1210) );
  INVX1 U800 ( .A(n1210), .Y(n1211) );
  AND2X2 U801 ( .A(\mem<19><14> ), .B(n276), .Y(n1212) );
  INVX1 U802 ( .A(n1212), .Y(n1213) );
  AND2X2 U803 ( .A(\mem<19><15> ), .B(n276), .Y(n1214) );
  INVX1 U804 ( .A(n1214), .Y(n1215) );
  AND2X2 U805 ( .A(\mem<18><11> ), .B(n278), .Y(n1216) );
  INVX1 U806 ( .A(n1216), .Y(n1217) );
  AND2X2 U807 ( .A(\mem<18><12> ), .B(n317), .Y(n1218) );
  INVX1 U808 ( .A(n1218), .Y(n1219) );
  AND2X2 U809 ( .A(\mem<18><13> ), .B(n278), .Y(n1220) );
  INVX1 U810 ( .A(n1220), .Y(n1221) );
  AND2X2 U811 ( .A(\mem<18><14> ), .B(n317), .Y(n1222) );
  INVX1 U812 ( .A(n1222), .Y(n1223) );
  AND2X2 U813 ( .A(\mem<18><15> ), .B(n278), .Y(n1224) );
  INVX1 U814 ( .A(n1224), .Y(n1225) );
  AND2X2 U815 ( .A(\mem<17><11> ), .B(n3), .Y(n1226) );
  INVX1 U816 ( .A(n1226), .Y(n1227) );
  AND2X2 U817 ( .A(\mem<17><12> ), .B(n3), .Y(n1228) );
  INVX1 U818 ( .A(n1228), .Y(n1229) );
  AND2X2 U819 ( .A(\mem<17><13> ), .B(n3), .Y(n1230) );
  INVX1 U820 ( .A(n1230), .Y(n1231) );
  AND2X2 U821 ( .A(\mem<17><14> ), .B(n3), .Y(n1232) );
  INVX1 U822 ( .A(n1232), .Y(n1233) );
  AND2X2 U823 ( .A(\mem<17><15> ), .B(n3), .Y(n1234) );
  INVX1 U824 ( .A(n1234), .Y(n1235) );
  AND2X2 U825 ( .A(\mem<16><11> ), .B(n321), .Y(n1236) );
  INVX1 U826 ( .A(n1236), .Y(n1237) );
  AND2X2 U827 ( .A(\mem<16><12> ), .B(n321), .Y(n1238) );
  INVX1 U828 ( .A(n1238), .Y(n1239) );
  AND2X2 U829 ( .A(\mem<16><13> ), .B(n321), .Y(n1240) );
  INVX1 U830 ( .A(n1240), .Y(n1241) );
  AND2X2 U831 ( .A(\mem<16><14> ), .B(n321), .Y(n1242) );
  INVX1 U832 ( .A(n1242), .Y(n1243) );
  AND2X2 U833 ( .A(\mem<16><15> ), .B(n321), .Y(n1244) );
  INVX1 U834 ( .A(n1244), .Y(n1245) );
  AND2X2 U835 ( .A(\mem<15><11> ), .B(n323), .Y(n1246) );
  INVX1 U836 ( .A(n1246), .Y(n1247) );
  AND2X2 U837 ( .A(\mem<15><12> ), .B(n323), .Y(n1248) );
  INVX1 U838 ( .A(n1248), .Y(n1249) );
  AND2X2 U839 ( .A(\mem<15><13> ), .B(n323), .Y(n1250) );
  INVX1 U840 ( .A(n1250), .Y(n1251) );
  AND2X2 U841 ( .A(\mem<15><14> ), .B(n323), .Y(n1252) );
  INVX1 U842 ( .A(n1252), .Y(n1253) );
  AND2X2 U843 ( .A(\mem<15><15> ), .B(n323), .Y(n1254) );
  INVX1 U844 ( .A(n1254), .Y(n1255) );
  AND2X2 U845 ( .A(\mem<14><11> ), .B(n325), .Y(n1256) );
  INVX1 U846 ( .A(n1256), .Y(n1257) );
  AND2X2 U847 ( .A(\mem<14><12> ), .B(n325), .Y(n1258) );
  INVX1 U848 ( .A(n1258), .Y(n1259) );
  AND2X2 U849 ( .A(\mem<14><13> ), .B(n325), .Y(n1260) );
  INVX1 U850 ( .A(n1260), .Y(n1261) );
  AND2X2 U851 ( .A(\mem<14><14> ), .B(n325), .Y(n1262) );
  INVX1 U852 ( .A(n1262), .Y(n1263) );
  AND2X2 U853 ( .A(\mem<14><15> ), .B(n325), .Y(n1264) );
  INVX1 U854 ( .A(n1264), .Y(n1265) );
  AND2X2 U855 ( .A(\mem<13><11> ), .B(n327), .Y(n1266) );
  INVX1 U856 ( .A(n1266), .Y(n1267) );
  AND2X2 U857 ( .A(\mem<13><12> ), .B(n327), .Y(n1268) );
  INVX1 U858 ( .A(n1268), .Y(n1269) );
  AND2X2 U859 ( .A(\mem<13><13> ), .B(n327), .Y(n1270) );
  INVX1 U860 ( .A(n1270), .Y(n1271) );
  AND2X2 U861 ( .A(\mem<13><14> ), .B(n327), .Y(n1272) );
  INVX1 U862 ( .A(n1272), .Y(n1273) );
  AND2X2 U863 ( .A(\mem<13><15> ), .B(n327), .Y(n1274) );
  INVX1 U864 ( .A(n1274), .Y(n1275) );
  AND2X2 U865 ( .A(\mem<12><11> ), .B(n329), .Y(n1276) );
  INVX1 U866 ( .A(n1276), .Y(n1277) );
  AND2X2 U867 ( .A(\mem<12><12> ), .B(n329), .Y(n1278) );
  INVX1 U868 ( .A(n1278), .Y(n1279) );
  AND2X2 U869 ( .A(\mem<12><13> ), .B(n329), .Y(n1280) );
  INVX1 U870 ( .A(n1280), .Y(n1281) );
  AND2X2 U871 ( .A(\mem<12><14> ), .B(n329), .Y(n1282) );
  INVX1 U872 ( .A(n1282), .Y(n1283) );
  AND2X2 U873 ( .A(\mem<12><15> ), .B(n329), .Y(n1284) );
  INVX1 U874 ( .A(n1284), .Y(n1285) );
  AND2X2 U875 ( .A(\mem<11><11> ), .B(n331), .Y(n1286) );
  INVX1 U876 ( .A(n1286), .Y(n1287) );
  AND2X2 U877 ( .A(\mem<11><12> ), .B(n331), .Y(n1288) );
  INVX1 U878 ( .A(n1288), .Y(n1289) );
  AND2X2 U879 ( .A(\mem<11><13> ), .B(n331), .Y(n1290) );
  INVX1 U880 ( .A(n1290), .Y(n1291) );
  AND2X2 U881 ( .A(\mem<11><14> ), .B(n331), .Y(n1292) );
  INVX1 U882 ( .A(n1292), .Y(n1293) );
  AND2X2 U883 ( .A(\mem<11><15> ), .B(n331), .Y(n1294) );
  INVX1 U884 ( .A(n1294), .Y(n1295) );
  AND2X2 U885 ( .A(\mem<10><11> ), .B(n333), .Y(n1296) );
  INVX1 U886 ( .A(n1296), .Y(n1297) );
  AND2X2 U887 ( .A(\mem<10><12> ), .B(n333), .Y(n1298) );
  INVX1 U888 ( .A(n1298), .Y(n1299) );
  AND2X2 U889 ( .A(\mem<10><13> ), .B(n333), .Y(n1300) );
  INVX1 U890 ( .A(n1300), .Y(n1301) );
  AND2X2 U891 ( .A(\mem<10><14> ), .B(n333), .Y(n1302) );
  INVX1 U892 ( .A(n1302), .Y(n1303) );
  AND2X2 U893 ( .A(\mem<10><15> ), .B(n333), .Y(n1304) );
  INVX1 U894 ( .A(n1304), .Y(n1305) );
  AND2X2 U895 ( .A(\mem<9><11> ), .B(n335), .Y(n1306) );
  INVX1 U896 ( .A(n1306), .Y(n1307) );
  AND2X2 U897 ( .A(\mem<9><12> ), .B(n335), .Y(n1308) );
  INVX1 U898 ( .A(n1308), .Y(n1309) );
  AND2X2 U899 ( .A(\mem<9><13> ), .B(n335), .Y(n1310) );
  INVX1 U900 ( .A(n1310), .Y(n1311) );
  AND2X2 U901 ( .A(\mem<9><14> ), .B(n335), .Y(n1312) );
  INVX1 U902 ( .A(n1312), .Y(n1313) );
  AND2X2 U903 ( .A(\mem<9><15> ), .B(n335), .Y(n1314) );
  INVX1 U904 ( .A(n1314), .Y(n1315) );
  AND2X2 U905 ( .A(\mem<8><0> ), .B(n281), .Y(n1316) );
  INVX1 U906 ( .A(n1316), .Y(n1317) );
  AND2X2 U907 ( .A(\mem<8><1> ), .B(n281), .Y(n1318) );
  INVX1 U908 ( .A(n1318), .Y(n1319) );
  AND2X2 U909 ( .A(\mem<8><2> ), .B(n281), .Y(n1320) );
  INVX1 U910 ( .A(n1320), .Y(n1321) );
  AND2X2 U911 ( .A(\mem<8><3> ), .B(n281), .Y(n1322) );
  INVX1 U912 ( .A(n1322), .Y(n1323) );
  AND2X2 U913 ( .A(\mem<8><4> ), .B(n281), .Y(n1324) );
  INVX1 U914 ( .A(n1324), .Y(n1325) );
  AND2X2 U915 ( .A(\mem<8><5> ), .B(n281), .Y(n1326) );
  INVX1 U916 ( .A(n1326), .Y(n1327) );
  AND2X2 U917 ( .A(\mem<8><6> ), .B(n281), .Y(n1328) );
  INVX1 U918 ( .A(n1328), .Y(n1329) );
  AND2X2 U919 ( .A(\mem<8><7> ), .B(n281), .Y(n1330) );
  INVX1 U920 ( .A(n1330), .Y(n1331) );
  AND2X2 U921 ( .A(\mem<8><8> ), .B(n281), .Y(n1332) );
  INVX1 U922 ( .A(n1332), .Y(n1333) );
  AND2X2 U923 ( .A(\mem<8><9> ), .B(n281), .Y(n1334) );
  INVX1 U924 ( .A(n1334), .Y(n1335) );
  AND2X2 U925 ( .A(\mem<8><10> ), .B(n281), .Y(n1336) );
  INVX1 U926 ( .A(n1336), .Y(n1337) );
  AND2X2 U927 ( .A(\mem<7><0> ), .B(n337), .Y(n1338) );
  INVX1 U928 ( .A(n1338), .Y(n1339) );
  AND2X2 U929 ( .A(\mem<7><1> ), .B(n337), .Y(n1340) );
  INVX1 U930 ( .A(n1340), .Y(n1341) );
  AND2X2 U931 ( .A(\mem<7><2> ), .B(n337), .Y(n1342) );
  INVX1 U932 ( .A(n1342), .Y(n1343) );
  AND2X2 U933 ( .A(\mem<7><3> ), .B(n337), .Y(n1344) );
  INVX1 U934 ( .A(n1344), .Y(n1345) );
  AND2X2 U935 ( .A(\mem<7><4> ), .B(n337), .Y(n1346) );
  INVX1 U936 ( .A(n1346), .Y(n1347) );
  AND2X2 U937 ( .A(\mem<7><5> ), .B(n337), .Y(n1348) );
  INVX1 U938 ( .A(n1348), .Y(n1349) );
  AND2X2 U939 ( .A(\mem<7><6> ), .B(n337), .Y(n1350) );
  INVX1 U940 ( .A(n1350), .Y(n1351) );
  AND2X2 U941 ( .A(\mem<7><7> ), .B(n337), .Y(n1352) );
  INVX1 U942 ( .A(n1352), .Y(n1353) );
  AND2X2 U943 ( .A(\mem<7><8> ), .B(n337), .Y(n1354) );
  INVX1 U944 ( .A(n1354), .Y(n1355) );
  AND2X2 U945 ( .A(\mem<7><9> ), .B(n337), .Y(n1356) );
  INVX1 U946 ( .A(n1356), .Y(n1357) );
  AND2X2 U947 ( .A(\mem<7><10> ), .B(n337), .Y(n1358) );
  INVX1 U948 ( .A(n1358), .Y(n1359) );
  AND2X2 U949 ( .A(\mem<6><0> ), .B(n339), .Y(n1360) );
  INVX1 U950 ( .A(n1360), .Y(n1361) );
  AND2X2 U951 ( .A(\mem<6><1> ), .B(n339), .Y(n1362) );
  INVX1 U952 ( .A(n1362), .Y(n1363) );
  AND2X2 U953 ( .A(\mem<6><2> ), .B(n339), .Y(n1364) );
  INVX1 U954 ( .A(n1364), .Y(n1365) );
  AND2X2 U955 ( .A(\mem<6><3> ), .B(n339), .Y(n1366) );
  INVX1 U956 ( .A(n1366), .Y(n1367) );
  AND2X2 U957 ( .A(\mem<6><4> ), .B(n339), .Y(n1368) );
  INVX1 U958 ( .A(n1368), .Y(n1369) );
  AND2X2 U959 ( .A(\mem<6><5> ), .B(n339), .Y(n1370) );
  INVX1 U960 ( .A(n1370), .Y(n1371) );
  AND2X2 U961 ( .A(\mem<6><6> ), .B(n339), .Y(n1372) );
  INVX1 U962 ( .A(n1372), .Y(n1373) );
  AND2X2 U963 ( .A(\mem<6><7> ), .B(n339), .Y(n1374) );
  INVX1 U964 ( .A(n1374), .Y(n1375) );
  AND2X2 U965 ( .A(\mem<6><8> ), .B(n283), .Y(n1376) );
  INVX1 U966 ( .A(n1376), .Y(n1377) );
  AND2X2 U967 ( .A(\mem<6><9> ), .B(n283), .Y(n1378) );
  INVX1 U968 ( .A(n1378), .Y(n1379) );
  AND2X2 U969 ( .A(\mem<6><10> ), .B(n283), .Y(n1380) );
  INVX1 U970 ( .A(n1380), .Y(n1381) );
  AND2X2 U971 ( .A(\mem<5><0> ), .B(n341), .Y(n1382) );
  INVX1 U972 ( .A(n1382), .Y(n1383) );
  AND2X2 U973 ( .A(\mem<5><1> ), .B(n341), .Y(n1384) );
  INVX1 U974 ( .A(n1384), .Y(n1385) );
  AND2X2 U975 ( .A(\mem<5><2> ), .B(n341), .Y(n1386) );
  INVX1 U976 ( .A(n1386), .Y(n1387) );
  AND2X2 U977 ( .A(\mem<5><3> ), .B(n341), .Y(n1388) );
  INVX1 U978 ( .A(n1388), .Y(n1389) );
  AND2X2 U979 ( .A(\mem<5><4> ), .B(n341), .Y(n1390) );
  INVX1 U980 ( .A(n1390), .Y(n1391) );
  AND2X2 U981 ( .A(\mem<5><5> ), .B(n341), .Y(n1392) );
  INVX1 U982 ( .A(n1392), .Y(n1393) );
  AND2X2 U983 ( .A(\mem<5><6> ), .B(n341), .Y(n1394) );
  INVX1 U984 ( .A(n1394), .Y(n1395) );
  AND2X2 U985 ( .A(\mem<5><7> ), .B(n341), .Y(n1396) );
  INVX1 U986 ( .A(n1396), .Y(n1397) );
  AND2X2 U987 ( .A(\mem<5><8> ), .B(n285), .Y(n1398) );
  INVX1 U988 ( .A(n1398), .Y(n1399) );
  AND2X2 U989 ( .A(\mem<5><9> ), .B(n285), .Y(n1400) );
  INVX1 U990 ( .A(n1400), .Y(n1401) );
  AND2X2 U991 ( .A(\mem<5><10> ), .B(n285), .Y(n1402) );
  INVX1 U992 ( .A(n1402), .Y(n1403) );
  AND2X2 U993 ( .A(\mem<4><0> ), .B(n343), .Y(n1404) );
  INVX1 U994 ( .A(n1404), .Y(n1405) );
  AND2X2 U995 ( .A(\mem<4><1> ), .B(n343), .Y(n1406) );
  INVX1 U996 ( .A(n1406), .Y(n1407) );
  AND2X2 U997 ( .A(\mem<4><2> ), .B(n343), .Y(n1408) );
  INVX1 U998 ( .A(n1408), .Y(n1409) );
  AND2X2 U999 ( .A(\mem<4><3> ), .B(n343), .Y(n1410) );
  INVX1 U1000 ( .A(n1410), .Y(n1411) );
  AND2X2 U1001 ( .A(\mem<4><4> ), .B(n343), .Y(n1412) );
  INVX1 U1002 ( .A(n1412), .Y(n1413) );
  AND2X2 U1003 ( .A(\mem<4><5> ), .B(n343), .Y(n1414) );
  INVX1 U1004 ( .A(n1414), .Y(n1415) );
  AND2X2 U1005 ( .A(\mem<4><6> ), .B(n343), .Y(n1416) );
  INVX1 U1006 ( .A(n1416), .Y(n1417) );
  AND2X2 U1007 ( .A(\mem<4><7> ), .B(n343), .Y(n1418) );
  INVX1 U1008 ( .A(n1418), .Y(n1419) );
  AND2X2 U1009 ( .A(\mem<4><8> ), .B(n343), .Y(n1420) );
  INVX1 U1010 ( .A(n1420), .Y(n1421) );
  AND2X2 U1011 ( .A(\mem<4><9> ), .B(n343), .Y(n1422) );
  INVX1 U1012 ( .A(n1422), .Y(n1423) );
  AND2X2 U1013 ( .A(\mem<4><10> ), .B(n343), .Y(n1424) );
  INVX1 U1014 ( .A(n1424), .Y(n1425) );
  AND2X2 U1015 ( .A(\mem<3><0> ), .B(n345), .Y(n1426) );
  INVX1 U1016 ( .A(n1426), .Y(n1427) );
  AND2X2 U1017 ( .A(\mem<3><1> ), .B(n345), .Y(n1428) );
  INVX1 U1018 ( .A(n1428), .Y(n1429) );
  AND2X2 U1019 ( .A(\mem<3><2> ), .B(n345), .Y(n1430) );
  INVX1 U1020 ( .A(n1430), .Y(n1431) );
  AND2X2 U1021 ( .A(\mem<3><3> ), .B(n345), .Y(n1432) );
  INVX1 U1022 ( .A(n1432), .Y(n1433) );
  AND2X2 U1023 ( .A(\mem<3><4> ), .B(n345), .Y(n1434) );
  INVX1 U1024 ( .A(n1434), .Y(n1435) );
  AND2X2 U1025 ( .A(\mem<3><5> ), .B(n345), .Y(n1436) );
  INVX1 U1026 ( .A(n1436), .Y(n1437) );
  AND2X2 U1027 ( .A(\mem<3><6> ), .B(n345), .Y(n1438) );
  INVX1 U1028 ( .A(n1438), .Y(n1439) );
  AND2X2 U1029 ( .A(\mem<3><7> ), .B(n345), .Y(n1440) );
  INVX1 U1030 ( .A(n1440), .Y(n1441) );
  AND2X2 U1031 ( .A(\mem<3><8> ), .B(n345), .Y(n1442) );
  INVX1 U1032 ( .A(n1442), .Y(n1443) );
  AND2X2 U1033 ( .A(\mem<3><9> ), .B(n345), .Y(n1444) );
  INVX1 U1034 ( .A(n1444), .Y(n1445) );
  AND2X2 U1035 ( .A(\mem<3><10> ), .B(n345), .Y(n1446) );
  INVX1 U1036 ( .A(n1446), .Y(n1447) );
  AND2X2 U1037 ( .A(\mem<2><0> ), .B(n347), .Y(n1448) );
  INVX1 U1038 ( .A(n1448), .Y(n1449) );
  AND2X2 U1039 ( .A(\mem<2><1> ), .B(n347), .Y(n1450) );
  INVX1 U1040 ( .A(n1450), .Y(n1451) );
  AND2X2 U1041 ( .A(\mem<2><2> ), .B(n347), .Y(n1452) );
  INVX1 U1042 ( .A(n1452), .Y(n1453) );
  AND2X2 U1043 ( .A(\mem<2><3> ), .B(n347), .Y(n1454) );
  INVX1 U1044 ( .A(n1454), .Y(n1455) );
  AND2X2 U1045 ( .A(\mem<2><4> ), .B(n347), .Y(n1456) );
  INVX1 U1046 ( .A(n1456), .Y(n1457) );
  AND2X2 U1047 ( .A(\mem<2><5> ), .B(n347), .Y(n1458) );
  INVX1 U1048 ( .A(n1458), .Y(n1459) );
  AND2X2 U1049 ( .A(\mem<2><6> ), .B(n347), .Y(n1460) );
  INVX1 U1050 ( .A(n1460), .Y(n1461) );
  AND2X2 U1051 ( .A(\mem<2><7> ), .B(n347), .Y(n1462) );
  INVX1 U1052 ( .A(n1462), .Y(n1463) );
  AND2X2 U1053 ( .A(\mem<2><8> ), .B(n347), .Y(n1464) );
  INVX1 U1054 ( .A(n1464), .Y(n1465) );
  AND2X2 U1055 ( .A(\mem<2><9> ), .B(n347), .Y(n1466) );
  INVX1 U1056 ( .A(n1466), .Y(n1467) );
  AND2X2 U1057 ( .A(\mem<2><10> ), .B(n347), .Y(n1468) );
  INVX1 U1058 ( .A(n1468), .Y(n1469) );
  AND2X2 U1059 ( .A(\mem<1><0> ), .B(n349), .Y(n1470) );
  INVX1 U1060 ( .A(n1470), .Y(n1471) );
  AND2X2 U1061 ( .A(\mem<1><1> ), .B(n349), .Y(n1472) );
  INVX1 U1062 ( .A(n1472), .Y(n1473) );
  AND2X2 U1063 ( .A(\mem<1><2> ), .B(n349), .Y(n1474) );
  INVX1 U1064 ( .A(n1474), .Y(n1475) );
  AND2X2 U1065 ( .A(\mem<1><3> ), .B(n349), .Y(n1476) );
  INVX1 U1066 ( .A(n1476), .Y(n1477) );
  AND2X2 U1067 ( .A(\mem<1><4> ), .B(n349), .Y(n1478) );
  INVX1 U1068 ( .A(n1478), .Y(n1479) );
  AND2X2 U1069 ( .A(\mem<1><5> ), .B(n349), .Y(n1480) );
  INVX1 U1070 ( .A(n1480), .Y(n1481) );
  AND2X2 U1071 ( .A(\mem<1><6> ), .B(n349), .Y(n1482) );
  INVX1 U1072 ( .A(n1482), .Y(n1483) );
  AND2X2 U1073 ( .A(\mem<1><7> ), .B(n349), .Y(n1484) );
  INVX1 U1074 ( .A(n1484), .Y(n1485) );
  AND2X2 U1075 ( .A(\mem<1><8> ), .B(n349), .Y(n1486) );
  INVX1 U1076 ( .A(n1486), .Y(n1487) );
  AND2X2 U1077 ( .A(\mem<1><9> ), .B(n349), .Y(n1488) );
  INVX1 U1078 ( .A(n1488), .Y(n1489) );
  AND2X2 U1079 ( .A(\mem<1><10> ), .B(n349), .Y(n1490) );
  INVX1 U1080 ( .A(n1490), .Y(n1491) );
  AND2X2 U1081 ( .A(\mem<0><11> ), .B(n351), .Y(n1492) );
  INVX1 U1082 ( .A(n1492), .Y(n1493) );
  AND2X2 U1083 ( .A(\mem<0><12> ), .B(n351), .Y(n1494) );
  INVX1 U1084 ( .A(n1494), .Y(n1495) );
  AND2X2 U1085 ( .A(\mem<0><13> ), .B(n351), .Y(n1496) );
  INVX1 U1086 ( .A(n1496), .Y(n1497) );
  AND2X2 U1087 ( .A(\mem<0><14> ), .B(n351), .Y(n1498) );
  INVX1 U1088 ( .A(n1498), .Y(n1499) );
  AND2X2 U1089 ( .A(\mem<0><15> ), .B(n351), .Y(n1500) );
  INVX1 U1090 ( .A(n1500), .Y(n1501) );
  INVX1 U1091 ( .A(n2335), .Y(n2334) );
  AND2X1 U1092 ( .A(n2185), .B(n2336), .Y(n1502) );
  INVX1 U1093 ( .A(n2337), .Y(n2336) );
  AND2X1 U1094 ( .A(n214), .B(n2341), .Y(n1503) );
  AND2X2 U1095 ( .A(\mem<8><11> ), .B(n281), .Y(n1504) );
  INVX1 U1096 ( .A(n1504), .Y(n1505) );
  AND2X2 U1097 ( .A(\mem<8><12> ), .B(n281), .Y(n1506) );
  INVX1 U1098 ( .A(n1506), .Y(n1507) );
  AND2X2 U1099 ( .A(\mem<8><13> ), .B(n281), .Y(n1508) );
  INVX1 U1100 ( .A(n1508), .Y(n1509) );
  AND2X2 U1101 ( .A(\mem<8><14> ), .B(n281), .Y(n1510) );
  INVX1 U1102 ( .A(n1510), .Y(n1511) );
  AND2X2 U1103 ( .A(\mem<8><15> ), .B(n281), .Y(n1512) );
  INVX1 U1104 ( .A(n1512), .Y(n1513) );
  AND2X2 U1105 ( .A(\mem<7><11> ), .B(n337), .Y(n1514) );
  INVX1 U1106 ( .A(n1514), .Y(n1515) );
  AND2X2 U1107 ( .A(\mem<7><12> ), .B(n337), .Y(n1516) );
  INVX1 U1108 ( .A(n1516), .Y(n1517) );
  AND2X2 U1109 ( .A(\mem<7><13> ), .B(n337), .Y(n1518) );
  INVX1 U1110 ( .A(n1518), .Y(n1519) );
  AND2X2 U1111 ( .A(\mem<7><14> ), .B(n337), .Y(n1520) );
  INVX1 U1112 ( .A(n1520), .Y(n1521) );
  AND2X2 U1113 ( .A(\mem<7><15> ), .B(n337), .Y(n1522) );
  INVX1 U1114 ( .A(n1522), .Y(n1523) );
  AND2X2 U1115 ( .A(\mem<6><11> ), .B(n283), .Y(n1524) );
  INVX1 U1116 ( .A(n1524), .Y(n1525) );
  AND2X2 U1117 ( .A(\mem<6><12> ), .B(n283), .Y(n1526) );
  INVX1 U1118 ( .A(n1526), .Y(n1527) );
  AND2X2 U1119 ( .A(\mem<6><13> ), .B(n339), .Y(n1528) );
  INVX1 U1120 ( .A(n1528), .Y(n1529) );
  AND2X2 U1121 ( .A(\mem<6><14> ), .B(n339), .Y(n1530) );
  INVX1 U1122 ( .A(n1530), .Y(n1531) );
  AND2X2 U1123 ( .A(\mem<6><15> ), .B(n339), .Y(n1532) );
  INVX1 U1124 ( .A(n1532), .Y(n1533) );
  AND2X2 U1125 ( .A(\mem<5><11> ), .B(n285), .Y(n1534) );
  INVX1 U1126 ( .A(n1534), .Y(n1535) );
  AND2X2 U1127 ( .A(\mem<5><12> ), .B(n285), .Y(n1536) );
  INVX1 U1128 ( .A(n1536), .Y(n1537) );
  AND2X2 U1129 ( .A(\mem<5><13> ), .B(n341), .Y(n1538) );
  INVX1 U1130 ( .A(n1538), .Y(n1539) );
  AND2X2 U1131 ( .A(\mem<5><14> ), .B(n341), .Y(n1540) );
  INVX1 U1132 ( .A(n1540), .Y(n1541) );
  AND2X2 U1133 ( .A(\mem<5><15> ), .B(n341), .Y(n1542) );
  INVX1 U1134 ( .A(n1542), .Y(n1543) );
  AND2X2 U1135 ( .A(\mem<4><11> ), .B(n343), .Y(n1544) );
  INVX1 U1136 ( .A(n1544), .Y(n1545) );
  AND2X2 U1137 ( .A(\mem<4><12> ), .B(n343), .Y(n1546) );
  INVX1 U1138 ( .A(n1546), .Y(n1547) );
  AND2X2 U1139 ( .A(\mem<4><13> ), .B(n343), .Y(n1548) );
  INVX1 U1140 ( .A(n1548), .Y(n1549) );
  AND2X2 U1141 ( .A(\mem<4><14> ), .B(n343), .Y(n1550) );
  INVX1 U1142 ( .A(n1550), .Y(n1551) );
  AND2X2 U1143 ( .A(\mem<4><15> ), .B(n343), .Y(n1552) );
  INVX1 U1144 ( .A(n1552), .Y(n1553) );
  AND2X2 U1145 ( .A(\mem<3><11> ), .B(n345), .Y(n1554) );
  INVX1 U1146 ( .A(n1554), .Y(n1555) );
  AND2X2 U1147 ( .A(\mem<3><12> ), .B(n345), .Y(n1556) );
  INVX1 U1148 ( .A(n1556), .Y(n1557) );
  AND2X2 U1149 ( .A(\mem<3><13> ), .B(n345), .Y(n1558) );
  INVX1 U1150 ( .A(n1558), .Y(n1559) );
  AND2X2 U1151 ( .A(\mem<3><14> ), .B(n345), .Y(n1560) );
  INVX1 U1152 ( .A(n1560), .Y(n1561) );
  AND2X2 U1153 ( .A(\mem<3><15> ), .B(n345), .Y(n1562) );
  INVX1 U1154 ( .A(n1562), .Y(n1563) );
  AND2X2 U1155 ( .A(\mem<2><11> ), .B(n347), .Y(n1564) );
  INVX1 U1156 ( .A(n1564), .Y(n1565) );
  AND2X2 U1157 ( .A(\mem<2><12> ), .B(n347), .Y(n1566) );
  INVX1 U1158 ( .A(n1566), .Y(n1567) );
  AND2X2 U1159 ( .A(\mem<2><13> ), .B(n347), .Y(n1568) );
  INVX1 U1160 ( .A(n1568), .Y(n1569) );
  AND2X2 U1161 ( .A(\mem<2><14> ), .B(n347), .Y(n1570) );
  INVX1 U1162 ( .A(n1570), .Y(n1571) );
  AND2X2 U1163 ( .A(\mem<2><15> ), .B(n347), .Y(n1572) );
  INVX1 U1164 ( .A(n1572), .Y(n1573) );
  AND2X2 U1165 ( .A(\mem<1><11> ), .B(n349), .Y(n1574) );
  INVX1 U1166 ( .A(n1574), .Y(n1575) );
  AND2X2 U1167 ( .A(\mem<1><12> ), .B(n349), .Y(n1576) );
  INVX1 U1168 ( .A(n1576), .Y(n1577) );
  AND2X2 U1169 ( .A(\mem<1><13> ), .B(n349), .Y(n1578) );
  INVX1 U1170 ( .A(n1578), .Y(n1579) );
  AND2X2 U1171 ( .A(\mem<1><14> ), .B(n349), .Y(n1580) );
  INVX1 U1172 ( .A(n1580), .Y(n1581) );
  AND2X2 U1173 ( .A(\mem<1><15> ), .B(n349), .Y(n1582) );
  INVX1 U1174 ( .A(n1582), .Y(n1583) );
  AND2X1 U1175 ( .A(N32), .B(n2333), .Y(n1584) );
  INVX1 U1177 ( .A(n1584), .Y(n1585) );
  AND2X1 U1178 ( .A(N31), .B(n2333), .Y(n1586) );
  INVX1 U1179 ( .A(n1586), .Y(n1587) );
  AND2X1 U1180 ( .A(N30), .B(n2333), .Y(n1588) );
  INVX1 U1181 ( .A(n1588), .Y(n1589) );
  AND2X1 U1182 ( .A(N29), .B(n2333), .Y(n1590) );
  INVX1 U1183 ( .A(n1590), .Y(n1591) );
  AND2X1 U1184 ( .A(N28), .B(n2333), .Y(n1592) );
  INVX1 U1185 ( .A(n1592), .Y(n1593) );
  AND2X1 U1186 ( .A(N27), .B(n2333), .Y(n1594) );
  INVX1 U1187 ( .A(n1594), .Y(n1595) );
  AND2X1 U1188 ( .A(N26), .B(n2333), .Y(n1596) );
  INVX1 U1189 ( .A(n1596), .Y(n1597) );
  AND2X1 U1190 ( .A(N25), .B(n2333), .Y(n1598) );
  INVX1 U1191 ( .A(n1598), .Y(n1599) );
  AND2X1 U1192 ( .A(N24), .B(n2333), .Y(n1600) );
  INVX1 U1193 ( .A(n1600), .Y(n1601) );
  AND2X1 U1194 ( .A(N23), .B(n2333), .Y(n1602) );
  INVX1 U1195 ( .A(n1602), .Y(n1603) );
  AND2X1 U1196 ( .A(N22), .B(n2333), .Y(n1604) );
  INVX1 U1197 ( .A(n1604), .Y(n1605) );
  AND2X1 U1198 ( .A(N21), .B(n2333), .Y(n1606) );
  INVX1 U1199 ( .A(n1606), .Y(n1607) );
  AND2X1 U1200 ( .A(N20), .B(n2333), .Y(n1608) );
  AND2X1 U1201 ( .A(N19), .B(n2333), .Y(n1609) );
  AND2X1 U1202 ( .A(N18), .B(n2333), .Y(n1610) );
  INVX1 U1203 ( .A(n1610), .Y(n1611) );
  AND2X1 U1204 ( .A(N17), .B(n2333), .Y(n1612) );
  INVX1 U1205 ( .A(n1612), .Y(n1613) );
  BUFX2 U1206 ( .A(n2360), .Y(n1614) );
  INVX1 U1207 ( .A(n1614), .Y(n2416) );
  BUFX2 U1208 ( .A(n2361), .Y(n1615) );
  INVX1 U1209 ( .A(n1615), .Y(n2417) );
  BUFX2 U1210 ( .A(n2362), .Y(n1616) );
  INVX1 U1211 ( .A(n1616), .Y(n2418) );
  BUFX2 U1212 ( .A(n2363), .Y(n1617) );
  INVX1 U1213 ( .A(n1617), .Y(n2419) );
  BUFX2 U1214 ( .A(n2372), .Y(n1618) );
  INVX1 U1215 ( .A(n1618), .Y(n2420) );
  BUFX2 U1216 ( .A(n2413), .Y(n1619) );
  INVX1 U1217 ( .A(n1619), .Y(n2414) );
  BUFX2 U1218 ( .A(n2415), .Y(n1620) );
  INVX1 U1219 ( .A(n1620), .Y(n2421) );
  AND2X1 U1220 ( .A(n2334), .B(n1502), .Y(n1621) );
  AND2X1 U1221 ( .A(n2339), .B(n1503), .Y(n1622) );
  AND2X1 U1222 ( .A(n2335), .B(n1502), .Y(n1623) );
  AND2X1 U1223 ( .A(n2340), .B(n1503), .Y(n1624) );
  AND2X1 U1224 ( .A(n1622), .B(n2422), .Y(n1625) );
  AND2X1 U1225 ( .A(n2422), .B(n1624), .Y(n1626) );
  AND2X1 U1226 ( .A(n2422), .B(n2414), .Y(n1627) );
  AND2X1 U1227 ( .A(n2422), .B(n2421), .Y(n1628) );
  AND2X1 U1228 ( .A(n1621), .B(n1622), .Y(n1629) );
  INVX1 U1229 ( .A(n1629), .Y(n1630) );
  AND2X1 U1230 ( .A(n1622), .B(n1623), .Y(n1631) );
  INVX1 U1231 ( .A(n1631), .Y(n1632) );
  AND2X1 U1232 ( .A(n1622), .B(n2416), .Y(n1633) );
  INVX1 U1233 ( .A(n1633), .Y(n1634) );
  BUFX2 U1234 ( .A(n620), .Y(n2242) );
  AND2X1 U1235 ( .A(n1622), .B(n2417), .Y(n1635) );
  INVX1 U1236 ( .A(n1635), .Y(n1636) );
  AND2X1 U1237 ( .A(n1622), .B(n2418), .Y(n1637) );
  INVX1 U1238 ( .A(n1637), .Y(n1638) );
  AND2X1 U1239 ( .A(n1622), .B(n2419), .Y(n1639) );
  INVX1 U1240 ( .A(n1639), .Y(n1640) );
  AND2X1 U1241 ( .A(n1622), .B(n2420), .Y(n1641) );
  INVX1 U1242 ( .A(n1641), .Y(n1642) );
  AND2X1 U1243 ( .A(n1621), .B(n1624), .Y(n1643) );
  INVX1 U1244 ( .A(n1643), .Y(n1644) );
  AND2X1 U1245 ( .A(n1623), .B(n1624), .Y(n1645) );
  INVX1 U1246 ( .A(n1645), .Y(n1646) );
  AND2X1 U1247 ( .A(n2416), .B(n1624), .Y(n1647) );
  INVX1 U1248 ( .A(n1647), .Y(n1648) );
  AND2X1 U1249 ( .A(n2417), .B(n1624), .Y(n1649) );
  INVX1 U1250 ( .A(n1649), .Y(n1650) );
  AND2X1 U1251 ( .A(n2418), .B(n1624), .Y(n1651) );
  INVX1 U1252 ( .A(n1651), .Y(n1652) );
  AND2X1 U1253 ( .A(n2419), .B(n1624), .Y(n1653) );
  INVX1 U1254 ( .A(n1653), .Y(n1654) );
  AND2X1 U1255 ( .A(n2420), .B(n1624), .Y(n1655) );
  INVX1 U1256 ( .A(n1655), .Y(n1656) );
  BUFX2 U1257 ( .A(n279), .Y(n2266) );
  AND2X1 U1258 ( .A(n1621), .B(n2414), .Y(n1657) );
  INVX1 U1259 ( .A(n1657), .Y(n1658) );
  AND2X1 U1260 ( .A(n1623), .B(n2414), .Y(n1659) );
  INVX1 U1261 ( .A(n1659), .Y(n1660) );
  AND2X1 U1262 ( .A(n2416), .B(n2414), .Y(n1661) );
  INVX1 U1263 ( .A(n1661), .Y(n1662) );
  AND2X1 U1264 ( .A(n2417), .B(n2414), .Y(n1663) );
  INVX1 U1265 ( .A(n1663), .Y(n1664) );
  AND2X1 U1266 ( .A(n2418), .B(n2414), .Y(n1665) );
  INVX1 U1267 ( .A(n1665), .Y(n1666) );
  AND2X1 U1268 ( .A(n2419), .B(n2414), .Y(n1667) );
  INVX1 U1269 ( .A(n1667), .Y(n1668) );
  AND2X1 U1270 ( .A(n2420), .B(n2414), .Y(n1669) );
  INVX1 U1271 ( .A(n1669), .Y(n1670) );
  AND2X1 U1272 ( .A(n1621), .B(n2421), .Y(n1671) );
  INVX1 U1273 ( .A(n1671), .Y(n1672) );
  AND2X1 U1274 ( .A(n1623), .B(n2421), .Y(n1673) );
  INVX1 U1275 ( .A(n1673), .Y(n1674) );
  AND2X1 U1276 ( .A(n2416), .B(n2421), .Y(n1675) );
  INVX1 U1277 ( .A(n1675), .Y(n1676) );
  AND2X1 U1278 ( .A(n2417), .B(n2421), .Y(n1677) );
  INVX1 U1279 ( .A(n1677), .Y(n1678) );
  AND2X1 U1280 ( .A(n2418), .B(n2421), .Y(n1679) );
  INVX1 U1281 ( .A(n1679), .Y(n1680) );
  AND2X1 U1282 ( .A(n2419), .B(n2421), .Y(n1681) );
  INVX1 U1283 ( .A(n1681), .Y(n1682) );
  AND2X1 U1284 ( .A(n2420), .B(n2421), .Y(n1683) );
  INVX1 U1285 ( .A(n1683), .Y(n1684) );
  INVX1 U1286 ( .A(N11), .Y(n2337) );
  MUX2X1 U1287 ( .B(n1686), .A(n1687), .S(n2193), .Y(n1685) );
  MUX2X1 U1288 ( .B(n1689), .A(n1690), .S(n2193), .Y(n1688) );
  MUX2X1 U1289 ( .B(n1692), .A(n1693), .S(n2193), .Y(n1691) );
  MUX2X1 U1290 ( .B(n1695), .A(n1696), .S(n2193), .Y(n1694) );
  MUX2X1 U1291 ( .B(n1698), .A(n1699), .S(n2184), .Y(n1697) );
  MUX2X1 U1292 ( .B(n1701), .A(n1702), .S(n2193), .Y(n1700) );
  MUX2X1 U1293 ( .B(n1704), .A(n1705), .S(n2193), .Y(n1703) );
  MUX2X1 U1294 ( .B(n1707), .A(n1708), .S(n2193), .Y(n1706) );
  MUX2X1 U1295 ( .B(n1710), .A(n1711), .S(n2193), .Y(n1709) );
  MUX2X1 U1296 ( .B(n1713), .A(n1714), .S(n2184), .Y(n1712) );
  MUX2X1 U1297 ( .B(n1716), .A(n1717), .S(n2194), .Y(n1715) );
  MUX2X1 U1298 ( .B(n1719), .A(n1720), .S(n2194), .Y(n1718) );
  MUX2X1 U1299 ( .B(n1722), .A(n1723), .S(n2194), .Y(n1721) );
  MUX2X1 U1300 ( .B(n1725), .A(n1726), .S(n2194), .Y(n1724) );
  MUX2X1 U1301 ( .B(n1728), .A(n1729), .S(n2184), .Y(n1727) );
  MUX2X1 U1302 ( .B(n1731), .A(n1732), .S(n2194), .Y(n1730) );
  MUX2X1 U1303 ( .B(n1734), .A(n1735), .S(n2194), .Y(n1733) );
  MUX2X1 U1304 ( .B(n1737), .A(n1738), .S(n2194), .Y(n1736) );
  MUX2X1 U1305 ( .B(n1740), .A(n1741), .S(n2194), .Y(n1739) );
  MUX2X1 U1306 ( .B(n1743), .A(n1744), .S(n2184), .Y(n1742) );
  MUX2X1 U1307 ( .B(n1746), .A(n1747), .S(n2194), .Y(n1745) );
  MUX2X1 U1308 ( .B(n1749), .A(n1750), .S(n2194), .Y(n1748) );
  MUX2X1 U1309 ( .B(n1752), .A(n1753), .S(n2194), .Y(n1751) );
  MUX2X1 U1310 ( .B(n1755), .A(n1756), .S(n2194), .Y(n1754) );
  MUX2X1 U1311 ( .B(n1758), .A(n1759), .S(n2184), .Y(n1757) );
  MUX2X1 U1312 ( .B(n1761), .A(n1762), .S(n2195), .Y(n1760) );
  MUX2X1 U1313 ( .B(n1764), .A(n1765), .S(n2195), .Y(n1763) );
  MUX2X1 U1314 ( .B(n1767), .A(n1768), .S(n2195), .Y(n1766) );
  MUX2X1 U1315 ( .B(n1770), .A(n1771), .S(n2195), .Y(n1769) );
  MUX2X1 U1316 ( .B(n1773), .A(n1774), .S(n2184), .Y(n1772) );
  MUX2X1 U1317 ( .B(n1776), .A(n1777), .S(n2195), .Y(n1775) );
  MUX2X1 U1318 ( .B(n1779), .A(n1780), .S(n2195), .Y(n1778) );
  MUX2X1 U1319 ( .B(n1782), .A(n1783), .S(n2195), .Y(n1781) );
  MUX2X1 U1320 ( .B(n1785), .A(n1786), .S(n2195), .Y(n1784) );
  MUX2X1 U1321 ( .B(n1788), .A(n1789), .S(n2184), .Y(n1787) );
  MUX2X1 U1322 ( .B(n1791), .A(n1792), .S(n2195), .Y(n1790) );
  MUX2X1 U1323 ( .B(n1794), .A(n1795), .S(n2195), .Y(n1793) );
  MUX2X1 U1324 ( .B(n1797), .A(n1798), .S(n2195), .Y(n1796) );
  MUX2X1 U1325 ( .B(n1800), .A(n1801), .S(n2195), .Y(n1799) );
  MUX2X1 U1326 ( .B(n1803), .A(n1804), .S(n2184), .Y(n1802) );
  MUX2X1 U1327 ( .B(n1806), .A(n1807), .S(n2196), .Y(n1805) );
  MUX2X1 U1328 ( .B(n1809), .A(n1810), .S(n2196), .Y(n1808) );
  MUX2X1 U1329 ( .B(n1812), .A(n1813), .S(n2196), .Y(n1811) );
  MUX2X1 U1330 ( .B(n1815), .A(n1816), .S(n2196), .Y(n1814) );
  MUX2X1 U1331 ( .B(n1818), .A(n1819), .S(n2184), .Y(n1817) );
  MUX2X1 U1332 ( .B(n1821), .A(n1822), .S(n2196), .Y(n1820) );
  MUX2X1 U1333 ( .B(n1824), .A(n1825), .S(n2196), .Y(n1823) );
  MUX2X1 U1334 ( .B(n1827), .A(n1828), .S(n2196), .Y(n1826) );
  MUX2X1 U1335 ( .B(n1830), .A(n1831), .S(n2196), .Y(n1829) );
  MUX2X1 U1336 ( .B(n1833), .A(n1834), .S(n2184), .Y(n1832) );
  MUX2X1 U1337 ( .B(n1836), .A(n1837), .S(n2196), .Y(n1835) );
  MUX2X1 U1338 ( .B(n1839), .A(n1840), .S(n2196), .Y(n1838) );
  MUX2X1 U1339 ( .B(n1842), .A(n1843), .S(n2196), .Y(n1841) );
  MUX2X1 U1340 ( .B(n1845), .A(n1846), .S(n2196), .Y(n1844) );
  MUX2X1 U1341 ( .B(n1848), .A(n1849), .S(n2184), .Y(n1847) );
  MUX2X1 U1342 ( .B(n1851), .A(n1852), .S(n2197), .Y(n1850) );
  MUX2X1 U1343 ( .B(n1854), .A(n1855), .S(n2197), .Y(n1853) );
  MUX2X1 U1344 ( .B(n1857), .A(n1858), .S(n2197), .Y(n1856) );
  MUX2X1 U1345 ( .B(n1860), .A(n1861), .S(n2197), .Y(n1859) );
  MUX2X1 U1346 ( .B(n1863), .A(n1864), .S(n2184), .Y(n1862) );
  MUX2X1 U1347 ( .B(n1866), .A(n1867), .S(n2197), .Y(n1865) );
  MUX2X1 U1348 ( .B(n1869), .A(n1870), .S(n2197), .Y(n1868) );
  MUX2X1 U1349 ( .B(n1872), .A(n1873), .S(n2197), .Y(n1871) );
  MUX2X1 U1350 ( .B(n1875), .A(n1876), .S(n2197), .Y(n1874) );
  MUX2X1 U1351 ( .B(n1878), .A(n1879), .S(n2183), .Y(n1877) );
  MUX2X1 U1352 ( .B(n1881), .A(n1882), .S(n2197), .Y(n1880) );
  MUX2X1 U1353 ( .B(n1884), .A(n1885), .S(n2197), .Y(n1883) );
  MUX2X1 U1354 ( .B(n1887), .A(n1888), .S(n2197), .Y(n1886) );
  MUX2X1 U1355 ( .B(n1890), .A(n1891), .S(n2197), .Y(n1889) );
  MUX2X1 U1356 ( .B(n1893), .A(n1894), .S(n2183), .Y(n1892) );
  MUX2X1 U1357 ( .B(n1896), .A(n1897), .S(n2198), .Y(n1895) );
  MUX2X1 U1358 ( .B(n1899), .A(n1900), .S(n2198), .Y(n1898) );
  MUX2X1 U1359 ( .B(n1902), .A(n1903), .S(n2198), .Y(n1901) );
  MUX2X1 U1360 ( .B(n1905), .A(n1906), .S(n2198), .Y(n1904) );
  MUX2X1 U1361 ( .B(n1908), .A(n1909), .S(n2183), .Y(n1907) );
  MUX2X1 U1362 ( .B(n1911), .A(n1912), .S(n2198), .Y(n1910) );
  MUX2X1 U1363 ( .B(n1914), .A(n1915), .S(n2198), .Y(n1913) );
  MUX2X1 U1364 ( .B(n1917), .A(n1918), .S(n2198), .Y(n1916) );
  MUX2X1 U1365 ( .B(n1920), .A(n1921), .S(n2198), .Y(n1919) );
  MUX2X1 U1366 ( .B(n1923), .A(n1924), .S(n2183), .Y(n1922) );
  MUX2X1 U1367 ( .B(n1926), .A(n1927), .S(n2198), .Y(n1925) );
  MUX2X1 U1368 ( .B(n1929), .A(n1930), .S(n2198), .Y(n1928) );
  MUX2X1 U1369 ( .B(n1932), .A(n1933), .S(n2198), .Y(n1931) );
  MUX2X1 U1370 ( .B(n1935), .A(n1936), .S(n2198), .Y(n1934) );
  MUX2X1 U1371 ( .B(n1938), .A(n1939), .S(n2183), .Y(n1937) );
  MUX2X1 U1372 ( .B(n1941), .A(n1942), .S(n2199), .Y(n1940) );
  MUX2X1 U1373 ( .B(n1944), .A(n1945), .S(n2199), .Y(n1943) );
  MUX2X1 U1374 ( .B(n1947), .A(n1948), .S(n2199), .Y(n1946) );
  MUX2X1 U1375 ( .B(n1950), .A(n1951), .S(n2199), .Y(n1949) );
  MUX2X1 U1376 ( .B(n1953), .A(n1954), .S(n2183), .Y(n1952) );
  MUX2X1 U1377 ( .B(n1956), .A(n1957), .S(n2199), .Y(n1955) );
  MUX2X1 U1378 ( .B(n1959), .A(n1960), .S(n2199), .Y(n1958) );
  MUX2X1 U1379 ( .B(n1962), .A(n1963), .S(n2199), .Y(n1961) );
  MUX2X1 U1380 ( .B(n1965), .A(n1966), .S(n2199), .Y(n1964) );
  MUX2X1 U1381 ( .B(n1968), .A(n1969), .S(n2183), .Y(n1967) );
  MUX2X1 U1382 ( .B(n1971), .A(n1972), .S(n2199), .Y(n1970) );
  MUX2X1 U1383 ( .B(n1974), .A(n1975), .S(n2199), .Y(n1973) );
  MUX2X1 U1384 ( .B(n1977), .A(n1978), .S(n2199), .Y(n1976) );
  MUX2X1 U1385 ( .B(n1980), .A(n1981), .S(n2199), .Y(n1979) );
  MUX2X1 U1386 ( .B(n1983), .A(n1984), .S(n2183), .Y(n1982) );
  MUX2X1 U1387 ( .B(n1986), .A(n1987), .S(n2200), .Y(n1985) );
  MUX2X1 U1388 ( .B(n1989), .A(n1990), .S(n2200), .Y(n1988) );
  MUX2X1 U1389 ( .B(n1992), .A(n1993), .S(n2200), .Y(n1991) );
  MUX2X1 U1390 ( .B(n1995), .A(n1996), .S(n2200), .Y(n1994) );
  MUX2X1 U1391 ( .B(n1998), .A(n1999), .S(n2183), .Y(n1997) );
  MUX2X1 U1392 ( .B(n2001), .A(n2002), .S(n2200), .Y(n2000) );
  MUX2X1 U1393 ( .B(n2004), .A(n2005), .S(n2200), .Y(n2003) );
  MUX2X1 U1394 ( .B(n2007), .A(n2008), .S(n2200), .Y(n2006) );
  MUX2X1 U1395 ( .B(n2010), .A(n2011), .S(n2200), .Y(n2009) );
  MUX2X1 U1396 ( .B(n2013), .A(n2014), .S(n2183), .Y(n2012) );
  MUX2X1 U1397 ( .B(n2016), .A(n2017), .S(n2200), .Y(n2015) );
  MUX2X1 U1398 ( .B(n2019), .A(n2020), .S(n2200), .Y(n2018) );
  MUX2X1 U1399 ( .B(n2022), .A(n2023), .S(n2200), .Y(n2021) );
  MUX2X1 U1400 ( .B(n2025), .A(n2026), .S(n2200), .Y(n2024) );
  MUX2X1 U1401 ( .B(n2028), .A(n2029), .S(n2183), .Y(n2027) );
  MUX2X1 U1402 ( .B(n2031), .A(n2032), .S(n2201), .Y(n2030) );
  MUX2X1 U1403 ( .B(n2034), .A(n2035), .S(n2201), .Y(n2033) );
  MUX2X1 U1404 ( .B(n2037), .A(n2038), .S(n2201), .Y(n2036) );
  MUX2X1 U1405 ( .B(n2040), .A(n2041), .S(n2201), .Y(n2039) );
  MUX2X1 U1406 ( .B(n2043), .A(n2044), .S(n2183), .Y(n2042) );
  MUX2X1 U1407 ( .B(n2046), .A(n2047), .S(n2201), .Y(n2045) );
  MUX2X1 U1408 ( .B(n2049), .A(n2050), .S(n2201), .Y(n2048) );
  MUX2X1 U1409 ( .B(n2052), .A(n2053), .S(n2201), .Y(n2051) );
  MUX2X1 U1410 ( .B(n2055), .A(n2056), .S(n2201), .Y(n2054) );
  MUX2X1 U1411 ( .B(n2058), .A(n2059), .S(n2184), .Y(n2057) );
  MUX2X1 U1412 ( .B(n2061), .A(n2062), .S(n2201), .Y(n2060) );
  MUX2X1 U1413 ( .B(n2064), .A(n2065), .S(n2201), .Y(n2063) );
  MUX2X1 U1414 ( .B(n2067), .A(n2068), .S(n2201), .Y(n2066) );
  MUX2X1 U1415 ( .B(n2070), .A(n2071), .S(n2201), .Y(n2069) );
  MUX2X1 U1416 ( .B(n2073), .A(n2074), .S(n2184), .Y(n2072) );
  MUX2X1 U1417 ( .B(n2076), .A(n2077), .S(n2202), .Y(n2075) );
  MUX2X1 U1418 ( .B(n2079), .A(n2080), .S(n2202), .Y(n2078) );
  MUX2X1 U1419 ( .B(n2082), .A(n2083), .S(n2202), .Y(n2081) );
  MUX2X1 U1420 ( .B(n2085), .A(n2086), .S(n2202), .Y(n2084) );
  MUX2X1 U1421 ( .B(n2088), .A(n2089), .S(n2339), .Y(n2087) );
  MUX2X1 U1422 ( .B(n2091), .A(n2092), .S(n2202), .Y(n2090) );
  MUX2X1 U1423 ( .B(n2094), .A(n2095), .S(n2202), .Y(n2093) );
  MUX2X1 U1424 ( .B(n2097), .A(n2098), .S(n2202), .Y(n2096) );
  MUX2X1 U1425 ( .B(n2100), .A(n2101), .S(n2202), .Y(n2099) );
  MUX2X1 U1426 ( .B(n2103), .A(n2104), .S(n2184), .Y(n2102) );
  MUX2X1 U1427 ( .B(n2106), .A(n2107), .S(n2202), .Y(n2105) );
  MUX2X1 U1428 ( .B(n2109), .A(n2110), .S(n2202), .Y(n2108) );
  MUX2X1 U1429 ( .B(n2112), .A(n2113), .S(n2202), .Y(n2111) );
  MUX2X1 U1430 ( .B(n2115), .A(n2116), .S(n2202), .Y(n2114) );
  MUX2X1 U1431 ( .B(n2118), .A(n2119), .S(n2184), .Y(n2117) );
  MUX2X1 U1432 ( .B(n2121), .A(n2122), .S(n2203), .Y(n2120) );
  MUX2X1 U1433 ( .B(n2124), .A(n2125), .S(n2203), .Y(n2123) );
  MUX2X1 U1434 ( .B(n2127), .A(n2128), .S(n2203), .Y(n2126) );
  MUX2X1 U1435 ( .B(n2130), .A(n2131), .S(n2203), .Y(n2129) );
  MUX2X1 U1436 ( .B(n2133), .A(n2134), .S(n2184), .Y(n2132) );
  MUX2X1 U1437 ( .B(n2136), .A(n2137), .S(n2203), .Y(n2135) );
  MUX2X1 U1438 ( .B(n2139), .A(n2140), .S(n2203), .Y(n2138) );
  MUX2X1 U1439 ( .B(n2142), .A(n2143), .S(n2203), .Y(n2141) );
  MUX2X1 U1440 ( .B(n2145), .A(n2146), .S(n2203), .Y(n2144) );
  MUX2X1 U1441 ( .B(n2148), .A(n2149), .S(n2339), .Y(n2147) );
  MUX2X1 U1442 ( .B(n2151), .A(n2152), .S(n2203), .Y(n2150) );
  MUX2X1 U1443 ( .B(n2154), .A(n2155), .S(n2203), .Y(n2153) );
  MUX2X1 U1444 ( .B(n2157), .A(n2158), .S(n2203), .Y(n2156) );
  MUX2X1 U1445 ( .B(n2160), .A(n2161), .S(n2203), .Y(n2159) );
  MUX2X1 U1446 ( .B(n2163), .A(n2164), .S(n2184), .Y(n2162) );
  MUX2X1 U1447 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n2212), .Y(n1687) );
  MUX2X1 U1448 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n2212), .Y(n1686) );
  MUX2X1 U1449 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n2212), .Y(n1690) );
  MUX2X1 U1450 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n2212), .Y(n1689) );
  MUX2X1 U1451 ( .B(n1688), .A(n1685), .S(n2190), .Y(n1699) );
  MUX2X1 U1452 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n2213), .Y(n1693) );
  MUX2X1 U1453 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n2213), .Y(n1692) );
  MUX2X1 U1454 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n2213), .Y(n1696) );
  MUX2X1 U1455 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n2213), .Y(n1695) );
  MUX2X1 U1456 ( .B(n1694), .A(n1691), .S(n2190), .Y(n1698) );
  MUX2X1 U1457 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n2213), .Y(n1702) );
  MUX2X1 U1458 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n2213), .Y(n1701) );
  MUX2X1 U1459 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n2213), .Y(n1705) );
  MUX2X1 U1460 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n2213), .Y(n1704) );
  MUX2X1 U1461 ( .B(n1703), .A(n1700), .S(n2190), .Y(n1714) );
  MUX2X1 U1462 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n2213), .Y(n1708) );
  MUX2X1 U1463 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n2213), .Y(n1707) );
  MUX2X1 U1464 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n2213), .Y(n1711) );
  MUX2X1 U1465 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n2213), .Y(n1710) );
  MUX2X1 U1466 ( .B(n1709), .A(n1706), .S(n2190), .Y(n1713) );
  MUX2X1 U1467 ( .B(n1712), .A(n1697), .S(n2182), .Y(n2165) );
  MUX2X1 U1468 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n2214), .Y(n1717) );
  MUX2X1 U1469 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n2214), .Y(n1716) );
  MUX2X1 U1470 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n2214), .Y(n1720) );
  MUX2X1 U1471 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n2214), .Y(n1719) );
  MUX2X1 U1472 ( .B(n1718), .A(n1715), .S(n2190), .Y(n1729) );
  MUX2X1 U1473 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n2214), .Y(n1723) );
  MUX2X1 U1474 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n2214), .Y(n1722) );
  MUX2X1 U1475 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n2214), .Y(n1726) );
  MUX2X1 U1476 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n2214), .Y(n1725) );
  MUX2X1 U1477 ( .B(n1724), .A(n1721), .S(n2190), .Y(n1728) );
  MUX2X1 U1478 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n2214), .Y(n1732) );
  MUX2X1 U1479 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n2214), .Y(n1731) );
  MUX2X1 U1480 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n2214), .Y(n1735) );
  MUX2X1 U1481 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n2214), .Y(n1734) );
  MUX2X1 U1482 ( .B(n1733), .A(n1730), .S(n2190), .Y(n1744) );
  MUX2X1 U1483 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n2215), .Y(n1738) );
  MUX2X1 U1484 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n2215), .Y(n1737) );
  MUX2X1 U1485 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n2215), .Y(n1741) );
  MUX2X1 U1486 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n2215), .Y(n1740) );
  MUX2X1 U1487 ( .B(n1739), .A(n1736), .S(n2190), .Y(n1743) );
  MUX2X1 U1488 ( .B(n1742), .A(n1727), .S(n2182), .Y(n2166) );
  MUX2X1 U1489 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n2215), .Y(n1747) );
  MUX2X1 U1490 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n2215), .Y(n1746) );
  MUX2X1 U1491 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n2215), .Y(n1750) );
  MUX2X1 U1492 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n2215), .Y(n1749) );
  MUX2X1 U1493 ( .B(n1748), .A(n1745), .S(n2190), .Y(n1759) );
  MUX2X1 U1494 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n2215), .Y(n1753) );
  MUX2X1 U1495 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n2215), .Y(n1752) );
  MUX2X1 U1496 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n2215), .Y(n1756) );
  MUX2X1 U1497 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n2215), .Y(n1755) );
  MUX2X1 U1498 ( .B(n1754), .A(n1751), .S(n2190), .Y(n1758) );
  MUX2X1 U1499 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n2216), .Y(n1762) );
  MUX2X1 U1500 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n2216), .Y(n1761) );
  MUX2X1 U1501 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n2216), .Y(n1765) );
  MUX2X1 U1502 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n2216), .Y(n1764) );
  MUX2X1 U1503 ( .B(n1763), .A(n1760), .S(n2190), .Y(n1774) );
  MUX2X1 U1504 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n2216), .Y(n1768) );
  MUX2X1 U1505 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n2216), .Y(n1767) );
  MUX2X1 U1506 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n2216), .Y(n1771) );
  MUX2X1 U1507 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n2216), .Y(n1770) );
  MUX2X1 U1508 ( .B(n1769), .A(n1766), .S(n2190), .Y(n1773) );
  MUX2X1 U1509 ( .B(n1772), .A(n1757), .S(n2182), .Y(n2167) );
  MUX2X1 U1510 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n2216), .Y(n1777) );
  MUX2X1 U1511 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n2216), .Y(n1776) );
  MUX2X1 U1512 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n2216), .Y(n1780) );
  MUX2X1 U1513 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n2216), .Y(n1779) );
  MUX2X1 U1514 ( .B(n1778), .A(n1775), .S(n2189), .Y(n1789) );
  MUX2X1 U1515 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n2217), .Y(n1783) );
  MUX2X1 U1516 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n2217), .Y(n1782) );
  MUX2X1 U1517 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n2217), .Y(n1786) );
  MUX2X1 U1518 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n2217), .Y(n1785) );
  MUX2X1 U1519 ( .B(n1784), .A(n1781), .S(n2189), .Y(n1788) );
  MUX2X1 U1520 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n2217), .Y(n1792) );
  MUX2X1 U1521 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n2217), .Y(n1791) );
  MUX2X1 U1522 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n2217), .Y(n1795) );
  MUX2X1 U1523 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n2217), .Y(n1794) );
  MUX2X1 U1524 ( .B(n1793), .A(n1790), .S(n2189), .Y(n1804) );
  MUX2X1 U1525 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n2217), .Y(n1798) );
  MUX2X1 U1526 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n2217), .Y(n1797) );
  MUX2X1 U1527 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n2217), .Y(n1801) );
  MUX2X1 U1528 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n2217), .Y(n1800) );
  MUX2X1 U1529 ( .B(n1799), .A(n1796), .S(n2189), .Y(n1803) );
  MUX2X1 U1530 ( .B(n1802), .A(n1787), .S(n2182), .Y(n2168) );
  MUX2X1 U1531 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n2218), .Y(n1807) );
  MUX2X1 U1532 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n2218), .Y(n1806) );
  MUX2X1 U1533 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n2218), .Y(n1810) );
  MUX2X1 U1534 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n2218), .Y(n1809) );
  MUX2X1 U1535 ( .B(n1808), .A(n1805), .S(n2189), .Y(n1819) );
  MUX2X1 U1536 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n2218), .Y(n1813) );
  MUX2X1 U1537 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n2218), .Y(n1812) );
  MUX2X1 U1538 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n2218), .Y(n1816) );
  MUX2X1 U1539 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n2218), .Y(n1815) );
  MUX2X1 U1540 ( .B(n1814), .A(n1811), .S(n2189), .Y(n1818) );
  MUX2X1 U1541 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n2218), .Y(n1822) );
  MUX2X1 U1542 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n2218), .Y(n1821) );
  MUX2X1 U1543 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n2218), .Y(n1825) );
  MUX2X1 U1544 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n2218), .Y(n1824) );
  MUX2X1 U1545 ( .B(n1823), .A(n1820), .S(n2189), .Y(n1834) );
  MUX2X1 U1546 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n2223), .Y(n1828) );
  MUX2X1 U1547 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n2223), .Y(n1827) );
  MUX2X1 U1548 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n2223), .Y(n1831) );
  MUX2X1 U1549 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n2223), .Y(n1830) );
  MUX2X1 U1550 ( .B(n1829), .A(n1826), .S(n2189), .Y(n1833) );
  MUX2X1 U1551 ( .B(n1832), .A(n1817), .S(n2182), .Y(n2169) );
  MUX2X1 U1552 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n2228), .Y(n1837) );
  MUX2X1 U1553 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n2212), .Y(n1836) );
  MUX2X1 U1554 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n2223), .Y(n1840) );
  MUX2X1 U1555 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n2223), .Y(n1839) );
  MUX2X1 U1556 ( .B(n1838), .A(n1835), .S(n2189), .Y(n1849) );
  MUX2X1 U1557 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n2228), .Y(n1843) );
  MUX2X1 U1558 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n2229), .Y(n1842) );
  MUX2X1 U1559 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n2223), .Y(n1846) );
  MUX2X1 U1560 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n2223), .Y(n1845) );
  MUX2X1 U1561 ( .B(n1844), .A(n1841), .S(n2189), .Y(n1848) );
  MUX2X1 U1562 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n2219), .Y(n1852) );
  MUX2X1 U1563 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n2219), .Y(n1851) );
  MUX2X1 U1564 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n2219), .Y(n1855) );
  MUX2X1 U1565 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n2219), .Y(n1854) );
  MUX2X1 U1566 ( .B(n1853), .A(n1850), .S(n2189), .Y(n1864) );
  MUX2X1 U1567 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n2219), .Y(n1858) );
  MUX2X1 U1568 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n2219), .Y(n1857) );
  MUX2X1 U1569 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n2219), .Y(n1861) );
  MUX2X1 U1570 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n2219), .Y(n1860) );
  MUX2X1 U1571 ( .B(n1859), .A(n1856), .S(n2189), .Y(n1863) );
  MUX2X1 U1572 ( .B(n1862), .A(n1847), .S(n2182), .Y(n2170) );
  MUX2X1 U1573 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n2219), .Y(n1867) );
  MUX2X1 U1574 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n2219), .Y(n1866) );
  MUX2X1 U1575 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n2219), .Y(n1870) );
  MUX2X1 U1576 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n2219), .Y(n1869) );
  MUX2X1 U1577 ( .B(n1868), .A(n1865), .S(n2188), .Y(n1879) );
  MUX2X1 U1578 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n2220), .Y(n1873) );
  MUX2X1 U1579 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n2220), .Y(n1872) );
  MUX2X1 U1580 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n2220), .Y(n1876) );
  MUX2X1 U1581 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n2220), .Y(n1875) );
  MUX2X1 U1582 ( .B(n1874), .A(n1871), .S(n2188), .Y(n1878) );
  MUX2X1 U1583 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n2220), .Y(n1882) );
  MUX2X1 U1584 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n2220), .Y(n1881) );
  MUX2X1 U1585 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n2220), .Y(n1885) );
  MUX2X1 U1586 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n2220), .Y(n1884) );
  MUX2X1 U1587 ( .B(n1883), .A(n1880), .S(n2188), .Y(n1894) );
  MUX2X1 U1588 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n2220), .Y(n1888) );
  MUX2X1 U1589 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n2220), .Y(n1887) );
  MUX2X1 U1590 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n2220), .Y(n1891) );
  MUX2X1 U1591 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n2220), .Y(n1890) );
  MUX2X1 U1592 ( .B(n1889), .A(n1886), .S(n2188), .Y(n1893) );
  MUX2X1 U1593 ( .B(n1892), .A(n1877), .S(n2182), .Y(n2171) );
  MUX2X1 U1594 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n2221), .Y(n1897) );
  MUX2X1 U1595 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n2221), .Y(n1896) );
  MUX2X1 U1596 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n2221), .Y(n1900) );
  MUX2X1 U1597 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n2221), .Y(n1899) );
  MUX2X1 U1598 ( .B(n1898), .A(n1895), .S(n2188), .Y(n1909) );
  MUX2X1 U1599 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n2221), .Y(n1903) );
  MUX2X1 U1600 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n2221), .Y(n1902) );
  MUX2X1 U1601 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n2221), .Y(n1906) );
  MUX2X1 U1602 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n2221), .Y(n1905) );
  MUX2X1 U1603 ( .B(n1904), .A(n1901), .S(n2188), .Y(n1908) );
  MUX2X1 U1604 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n2221), .Y(n1912) );
  MUX2X1 U1605 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n2221), .Y(n1911) );
  MUX2X1 U1606 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n2221), .Y(n1915) );
  MUX2X1 U1607 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n2221), .Y(n1914) );
  MUX2X1 U1608 ( .B(n1913), .A(n1910), .S(n2188), .Y(n1924) );
  MUX2X1 U1609 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n2222), .Y(n1918) );
  MUX2X1 U1610 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n2222), .Y(n1917) );
  MUX2X1 U1611 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n2222), .Y(n1921) );
  MUX2X1 U1612 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n2222), .Y(n1920) );
  MUX2X1 U1613 ( .B(n1919), .A(n1916), .S(n2188), .Y(n1923) );
  MUX2X1 U1614 ( .B(n1922), .A(n1907), .S(n2182), .Y(n2172) );
  MUX2X1 U1615 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n2222), .Y(n1927) );
  MUX2X1 U1616 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n2222), .Y(n1926) );
  MUX2X1 U1617 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n2222), .Y(n1930) );
  MUX2X1 U1618 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n2222), .Y(n1929) );
  MUX2X1 U1619 ( .B(n1928), .A(n1925), .S(n2188), .Y(n1939) );
  MUX2X1 U1620 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n2222), .Y(n1933) );
  MUX2X1 U1621 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n2222), .Y(n1932) );
  MUX2X1 U1622 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n2222), .Y(n1936) );
  MUX2X1 U1623 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n2222), .Y(n1935) );
  MUX2X1 U1624 ( .B(n1934), .A(n1931), .S(n2188), .Y(n1938) );
  MUX2X1 U1625 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n2223), .Y(n1942) );
  MUX2X1 U1626 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n2223), .Y(n1941) );
  MUX2X1 U1627 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n2223), .Y(n1945) );
  MUX2X1 U1628 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n2223), .Y(n1944) );
  MUX2X1 U1629 ( .B(n1943), .A(n1940), .S(n2188), .Y(n1954) );
  MUX2X1 U1630 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n2223), .Y(n1948) );
  MUX2X1 U1631 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n2223), .Y(n1947) );
  MUX2X1 U1632 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n2223), .Y(n1951) );
  MUX2X1 U1633 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n2223), .Y(n1950) );
  MUX2X1 U1634 ( .B(n1949), .A(n1946), .S(n2188), .Y(n1953) );
  MUX2X1 U1635 ( .B(n1952), .A(n1937), .S(n2182), .Y(n2173) );
  MUX2X1 U1636 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n2223), .Y(n1957) );
  MUX2X1 U1637 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n2223), .Y(n1956) );
  MUX2X1 U1638 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n2223), .Y(n1960) );
  MUX2X1 U1639 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n2223), .Y(n1959) );
  MUX2X1 U1640 ( .B(n1958), .A(n1955), .S(n2187), .Y(n1969) );
  MUX2X1 U1641 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n2224), .Y(n1963) );
  MUX2X1 U1642 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n2224), .Y(n1962) );
  MUX2X1 U1643 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n2224), .Y(n1966) );
  MUX2X1 U1644 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n2224), .Y(n1965) );
  MUX2X1 U1645 ( .B(n1964), .A(n1961), .S(n2187), .Y(n1968) );
  MUX2X1 U1646 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n2224), .Y(n1972) );
  MUX2X1 U1647 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n2224), .Y(n1971) );
  MUX2X1 U1648 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n2224), .Y(n1975) );
  MUX2X1 U1649 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n2224), .Y(n1974) );
  MUX2X1 U1650 ( .B(n1973), .A(n1970), .S(n2187), .Y(n1984) );
  MUX2X1 U1651 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n2224), .Y(n1978) );
  MUX2X1 U1652 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n2224), .Y(n1977) );
  MUX2X1 U1653 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n2224), .Y(n1981) );
  MUX2X1 U1654 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n2224), .Y(n1980) );
  MUX2X1 U1655 ( .B(n1979), .A(n1976), .S(n2187), .Y(n1983) );
  MUX2X1 U1656 ( .B(n1982), .A(n1967), .S(n2182), .Y(n2174) );
  MUX2X1 U1657 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n2225), .Y(n1987) );
  MUX2X1 U1658 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n2225), .Y(n1986) );
  MUX2X1 U1659 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n2225), .Y(n1990) );
  MUX2X1 U1660 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n2225), .Y(n1989) );
  MUX2X1 U1661 ( .B(n1988), .A(n1985), .S(n2187), .Y(n1999) );
  MUX2X1 U1662 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n2225), .Y(n1993) );
  MUX2X1 U1663 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n2225), .Y(n1992) );
  MUX2X1 U1664 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n2225), .Y(n1996) );
  MUX2X1 U1665 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n2225), .Y(n1995) );
  MUX2X1 U1666 ( .B(n1994), .A(n1991), .S(n2187), .Y(n1998) );
  MUX2X1 U1667 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n2225), .Y(n2002) );
  MUX2X1 U1668 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n2225), .Y(n2001) );
  MUX2X1 U1669 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n2225), .Y(n2005) );
  MUX2X1 U1670 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n2225), .Y(n2004) );
  MUX2X1 U1671 ( .B(n2003), .A(n2000), .S(n2187), .Y(n2014) );
  MUX2X1 U1672 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n2226), .Y(n2008) );
  MUX2X1 U1673 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n2226), .Y(n2007) );
  MUX2X1 U1674 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n2226), .Y(n2011) );
  MUX2X1 U1675 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n2226), .Y(n2010) );
  MUX2X1 U1676 ( .B(n2009), .A(n2006), .S(n2187), .Y(n2013) );
  MUX2X1 U1677 ( .B(n2012), .A(n1997), .S(n2182), .Y(n2175) );
  MUX2X1 U1678 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n2226), .Y(n2017) );
  MUX2X1 U1679 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n2226), .Y(n2016) );
  MUX2X1 U1680 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n2226), .Y(n2020) );
  MUX2X1 U1681 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n2226), .Y(n2019) );
  MUX2X1 U1682 ( .B(n2018), .A(n2015), .S(n2187), .Y(n2029) );
  MUX2X1 U1683 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n2226), .Y(n2023) );
  MUX2X1 U1684 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n2226), .Y(n2022) );
  MUX2X1 U1685 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n2226), .Y(n2026) );
  MUX2X1 U1686 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n2226), .Y(n2025) );
  MUX2X1 U1687 ( .B(n2024), .A(n2021), .S(n2187), .Y(n2028) );
  MUX2X1 U1688 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n2227), .Y(n2032) );
  MUX2X1 U1689 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n2227), .Y(n2031) );
  MUX2X1 U1690 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n2227), .Y(n2035) );
  MUX2X1 U1691 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n2227), .Y(n2034) );
  MUX2X1 U1692 ( .B(n2033), .A(n2030), .S(n2187), .Y(n2044) );
  MUX2X1 U1693 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n2227), .Y(n2038) );
  MUX2X1 U1694 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n2227), .Y(n2037) );
  MUX2X1 U1695 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n2227), .Y(n2041) );
  MUX2X1 U1696 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n2227), .Y(n2040) );
  MUX2X1 U1697 ( .B(n2039), .A(n2036), .S(n2187), .Y(n2043) );
  MUX2X1 U1698 ( .B(n2042), .A(n2027), .S(n2182), .Y(n2176) );
  MUX2X1 U1699 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n2227), .Y(n2047) );
  MUX2X1 U1700 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n2227), .Y(n2046) );
  MUX2X1 U1701 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n2227), .Y(n2050) );
  MUX2X1 U1702 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n2227), .Y(n2049) );
  MUX2X1 U1703 ( .B(n2048), .A(n2045), .S(n2186), .Y(n2059) );
  MUX2X1 U1704 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n2228), .Y(n2053) );
  MUX2X1 U1705 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n2228), .Y(n2052) );
  MUX2X1 U1706 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n2228), .Y(n2056) );
  MUX2X1 U1707 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n2228), .Y(n2055) );
  MUX2X1 U1708 ( .B(n2054), .A(n2051), .S(n2186), .Y(n2058) );
  MUX2X1 U1709 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n2228), .Y(n2062) );
  MUX2X1 U1710 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n2228), .Y(n2061) );
  MUX2X1 U1711 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n2228), .Y(n2065) );
  MUX2X1 U1712 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n2228), .Y(n2064) );
  MUX2X1 U1713 ( .B(n2063), .A(n2060), .S(n2186), .Y(n2074) );
  MUX2X1 U1714 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n2228), .Y(n2068) );
  MUX2X1 U1715 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n2228), .Y(n2067) );
  MUX2X1 U1716 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n2228), .Y(n2071) );
  MUX2X1 U1717 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n2228), .Y(n2070) );
  MUX2X1 U1718 ( .B(n2069), .A(n2066), .S(n2186), .Y(n2073) );
  MUX2X1 U1719 ( .B(n2072), .A(n2057), .S(n2181), .Y(n2177) );
  MUX2X1 U1720 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n2229), .Y(n2077) );
  MUX2X1 U1721 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n2229), .Y(n2076) );
  MUX2X1 U1722 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n2229), .Y(n2080) );
  MUX2X1 U1723 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n2229), .Y(n2079) );
  MUX2X1 U1724 ( .B(n2078), .A(n2075), .S(n2186), .Y(n2089) );
  MUX2X1 U1725 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n2229), .Y(n2083) );
  MUX2X1 U1726 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n2229), .Y(n2082) );
  MUX2X1 U1727 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n2229), .Y(n2086) );
  MUX2X1 U1728 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n2229), .Y(n2085) );
  MUX2X1 U1729 ( .B(n2084), .A(n2081), .S(n2186), .Y(n2088) );
  MUX2X1 U1730 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n2229), .Y(n2092) );
  MUX2X1 U1731 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n2229), .Y(n2091) );
  MUX2X1 U1732 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n2229), .Y(n2095) );
  MUX2X1 U1733 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n2229), .Y(n2094) );
  MUX2X1 U1734 ( .B(n2093), .A(n2090), .S(n2186), .Y(n2104) );
  MUX2X1 U1735 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n2230), .Y(n2098) );
  MUX2X1 U1736 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n2230), .Y(n2097) );
  MUX2X1 U1737 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n2230), .Y(n2101) );
  MUX2X1 U1738 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n2230), .Y(n2100) );
  MUX2X1 U1739 ( .B(n2099), .A(n2096), .S(n2186), .Y(n2103) );
  MUX2X1 U1740 ( .B(n2102), .A(n2087), .S(n2181), .Y(n2178) );
  MUX2X1 U1741 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n2230), .Y(n2107) );
  MUX2X1 U1742 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n2230), .Y(n2106) );
  MUX2X1 U1743 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n2230), .Y(n2110) );
  MUX2X1 U1744 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n2230), .Y(n2109) );
  MUX2X1 U1745 ( .B(n2108), .A(n2105), .S(n2186), .Y(n2119) );
  MUX2X1 U1746 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n2230), .Y(n2113) );
  MUX2X1 U1747 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n2230), .Y(n2112) );
  MUX2X1 U1748 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n2230), .Y(n2116) );
  MUX2X1 U1749 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n2230), .Y(n2115) );
  MUX2X1 U1750 ( .B(n2114), .A(n2111), .S(n2186), .Y(n2118) );
  MUX2X1 U1751 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n2231), .Y(n2122) );
  MUX2X1 U1752 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n2231), .Y(n2121) );
  MUX2X1 U1753 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n2231), .Y(n2125) );
  MUX2X1 U1754 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n2231), .Y(n2124) );
  MUX2X1 U1755 ( .B(n2123), .A(n2120), .S(n2186), .Y(n2134) );
  MUX2X1 U1756 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n2231), .Y(n2128) );
  MUX2X1 U1757 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n2231), .Y(n2127) );
  MUX2X1 U1758 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n2231), .Y(n2131) );
  MUX2X1 U1759 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n2231), .Y(n2130) );
  MUX2X1 U1760 ( .B(n2129), .A(n2126), .S(n2186), .Y(n2133) );
  MUX2X1 U1761 ( .B(n2132), .A(n2117), .S(n2181), .Y(n2179) );
  MUX2X1 U1762 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n2231), .Y(n2137) );
  MUX2X1 U1763 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n2231), .Y(n2136) );
  MUX2X1 U1764 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n2231), .Y(n2140) );
  MUX2X1 U1765 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n2231), .Y(n2139) );
  MUX2X1 U1766 ( .B(n2138), .A(n2135), .S(n2185), .Y(n2149) );
  MUX2X1 U1767 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n2232), .Y(n2143) );
  MUX2X1 U1768 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n2232), .Y(n2142) );
  MUX2X1 U1769 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n2232), .Y(n2146) );
  MUX2X1 U1770 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n2232), .Y(n2145) );
  MUX2X1 U1771 ( .B(n2144), .A(n2141), .S(n2185), .Y(n2148) );
  MUX2X1 U1772 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n2232), .Y(n2152) );
  MUX2X1 U1773 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n2232), .Y(n2151) );
  MUX2X1 U1774 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n2232), .Y(n2155) );
  MUX2X1 U1775 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n2232), .Y(n2154) );
  MUX2X1 U1776 ( .B(n2153), .A(n2150), .S(n2185), .Y(n2164) );
  MUX2X1 U1777 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n2232), .Y(n2158) );
  MUX2X1 U1778 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n2232), .Y(n2157) );
  MUX2X1 U1779 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n2232), .Y(n2161) );
  MUX2X1 U1780 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n2232), .Y(n2160) );
  MUX2X1 U1781 ( .B(n2159), .A(n2156), .S(n2185), .Y(n2163) );
  MUX2X1 U1782 ( .B(n2162), .A(n2147), .S(n2181), .Y(n2180) );
  INVX8 U1783 ( .A(n2204), .Y(n2191) );
  INVX8 U1784 ( .A(n2204), .Y(n2192) );
  INVX8 U1785 ( .A(n2192), .Y(n2194) );
  INVX8 U1786 ( .A(n2192), .Y(n2195) );
  INVX8 U1787 ( .A(n2191), .Y(n2196) );
  INVX8 U1788 ( .A(n2191), .Y(n2197) );
  INVX8 U1789 ( .A(n2191), .Y(n2198) );
  INVX8 U1790 ( .A(n2192), .Y(n2200) );
  INVX8 U1791 ( .A(n2191), .Y(n2201) );
  INVX8 U1792 ( .A(n2191), .Y(n2202) );
  INVX8 U1793 ( .A(n2192), .Y(n2203) );
  INVX8 U1794 ( .A(n2234), .Y(n2206) );
  INVX8 U1795 ( .A(n2234), .Y(n2207) );
  INVX8 U1796 ( .A(n2234), .Y(n2208) );
  INVX8 U1797 ( .A(n2235), .Y(n2209) );
  INVX8 U1798 ( .A(n2235), .Y(n2210) );
  INVX8 U1799 ( .A(n2211), .Y(n2213) );
  INVX8 U1800 ( .A(n2211), .Y(n2214) );
  INVX8 U1801 ( .A(n2210), .Y(n2215) );
  INVX8 U1802 ( .A(n2210), .Y(n2216) );
  INVX8 U1803 ( .A(n2210), .Y(n2217) );
  INVX8 U1804 ( .A(n2209), .Y(n2218) );
  INVX8 U1805 ( .A(n2209), .Y(n2219) );
  INVX8 U1806 ( .A(n2208), .Y(n2220) );
  INVX8 U1807 ( .A(n2208), .Y(n2221) );
  INVX8 U1808 ( .A(n2208), .Y(n2222) );
  INVX8 U1809 ( .A(n2233), .Y(n2223) );
  INVX8 U1810 ( .A(n2211), .Y(n2224) );
  INVX8 U1811 ( .A(n2205), .Y(n2225) );
  INVX8 U1812 ( .A(n2207), .Y(n2226) );
  INVX8 U1813 ( .A(n2207), .Y(n2227) );
  INVX8 U1814 ( .A(n2207), .Y(n2228) );
  INVX8 U1815 ( .A(n2206), .Y(n2229) );
  INVX8 U1816 ( .A(n2206), .Y(n2230) );
  INVX8 U1817 ( .A(n2206), .Y(n2231) );
  INVX8 U1818 ( .A(n2205), .Y(n2232) );
  INVX8 U1819 ( .A(n2233), .Y(n2234) );
  INVX8 U1820 ( .A(n2233), .Y(n2235) );
  INVX1 U1821 ( .A(N10), .Y(n2335) );
  INVX1 U1822 ( .A(n2423), .Y(n2298) );
  INVX4 U1823 ( .A(n1171), .Y(n2332) );
  INVX4 U1824 ( .A(n1166), .Y(n2323) );
  INVX8 U1825 ( .A(n4), .Y(n2299) );
  INVX8 U1826 ( .A(n642), .Y(n2300) );
  INVX8 U1827 ( .A(n643), .Y(n2301) );
  INVX8 U1828 ( .A(n643), .Y(n2302) );
  INVX8 U1829 ( .A(n644), .Y(n2303) );
  INVX8 U1830 ( .A(n644), .Y(n2304) );
  INVX8 U1831 ( .A(n645), .Y(n2305) );
  INVX8 U1832 ( .A(n645), .Y(n2306) );
  INVX8 U1833 ( .A(n646), .Y(n2307) );
  INVX8 U1834 ( .A(n646), .Y(n2308) );
  INVX8 U1835 ( .A(n647), .Y(n2309) );
  INVX8 U1836 ( .A(n647), .Y(n2310) );
  INVX8 U1837 ( .A(n648), .Y(n2311) );
  INVX8 U1838 ( .A(n648), .Y(n2312) );
  INVX8 U1839 ( .A(n649), .Y(n2313) );
  INVX8 U1840 ( .A(n649), .Y(n2314) );
  INVX8 U1841 ( .A(n650), .Y(n2315) );
  INVX8 U1842 ( .A(n650), .Y(n2316) );
  INVX8 U1843 ( .A(n1163), .Y(n2317) );
  INVX8 U1844 ( .A(n1163), .Y(n2318) );
  INVX8 U1845 ( .A(n1164), .Y(n2319) );
  INVX8 U1846 ( .A(n1164), .Y(n2320) );
  INVX8 U1847 ( .A(n2323), .Y(n2321) );
  INVX8 U1848 ( .A(n2323), .Y(n2322) );
  INVX8 U1849 ( .A(n1167), .Y(n2324) );
  INVX8 U1850 ( .A(n1167), .Y(n2325) );
  INVX8 U1851 ( .A(n1168), .Y(n2326) );
  INVX8 U1852 ( .A(n1168), .Y(n2327) );
  INVX8 U1853 ( .A(n1169), .Y(n2328) );
  INVX8 U1854 ( .A(n1169), .Y(n2329) );
  INVX8 U1855 ( .A(n2332), .Y(n2330) );
  INVX8 U1856 ( .A(n2332), .Y(n2331) );
  NAND2X1 U1857 ( .A(\mem<31><0> ), .B(n315), .Y(n2344) );
  OAI21X1 U1858 ( .A(n2237), .B(n2299), .C(n2344), .Y(n651) );
  NAND2X1 U1859 ( .A(\mem<31><1> ), .B(n315), .Y(n2345) );
  OAI21X1 U1860 ( .A(n2302), .B(n2236), .C(n2345), .Y(n652) );
  NAND2X1 U1861 ( .A(\mem<31><2> ), .B(n315), .Y(n2346) );
  OAI21X1 U1862 ( .A(n2304), .B(n2236), .C(n2346), .Y(n653) );
  NAND2X1 U1863 ( .A(\mem<31><3> ), .B(n315), .Y(n2347) );
  OAI21X1 U1864 ( .A(n2306), .B(n2236), .C(n2347), .Y(n654) );
  NAND2X1 U1865 ( .A(\mem<31><4> ), .B(n315), .Y(n2348) );
  OAI21X1 U1866 ( .A(n2308), .B(n2236), .C(n2348), .Y(n655) );
  NAND2X1 U1867 ( .A(\mem<31><5> ), .B(n315), .Y(n2349) );
  OAI21X1 U1868 ( .A(n2310), .B(n2236), .C(n2349), .Y(n656) );
  NAND2X1 U1869 ( .A(\mem<31><6> ), .B(n315), .Y(n2350) );
  OAI21X1 U1870 ( .A(n2312), .B(n2236), .C(n2350), .Y(n657) );
  NAND2X1 U1871 ( .A(\mem<31><7> ), .B(n315), .Y(n2351) );
  OAI21X1 U1872 ( .A(n2314), .B(n2236), .C(n2351), .Y(n658) );
  NAND2X1 U1873 ( .A(\mem<31><8> ), .B(n315), .Y(n2352) );
  OAI21X1 U1874 ( .A(n2316), .B(n2236), .C(n2352), .Y(n659) );
  NAND2X1 U1875 ( .A(\mem<31><9> ), .B(n315), .Y(n2353) );
  OAI21X1 U1876 ( .A(n2317), .B(n2237), .C(n2353), .Y(n660) );
  NAND2X1 U1877 ( .A(\mem<31><10> ), .B(n315), .Y(n2354) );
  OAI21X1 U1878 ( .A(n2319), .B(n2237), .C(n2354), .Y(n661) );
  NAND2X1 U1879 ( .A(\mem<31><11> ), .B(n315), .Y(n2355) );
  OAI21X1 U1880 ( .A(n2321), .B(n2237), .C(n2355), .Y(n662) );
  NAND2X1 U1881 ( .A(\mem<31><12> ), .B(n315), .Y(n2356) );
  OAI21X1 U1882 ( .A(n2324), .B(n2237), .C(n2356), .Y(n663) );
  NAND2X1 U1883 ( .A(\mem<31><13> ), .B(n315), .Y(n2357) );
  OAI21X1 U1884 ( .A(n2326), .B(n2237), .C(n2357), .Y(n664) );
  NAND2X1 U1885 ( .A(\mem<31><14> ), .B(n315), .Y(n2358) );
  OAI21X1 U1886 ( .A(n2329), .B(n2237), .C(n2358), .Y(n665) );
  NAND2X1 U1887 ( .A(\mem<31><15> ), .B(n315), .Y(n2359) );
  OAI21X1 U1888 ( .A(n2330), .B(n2237), .C(n2359), .Y(n666) );
  OAI21X1 U1889 ( .A(n2238), .B(n2299), .C(n16), .Y(n667) );
  OAI21X1 U1890 ( .A(n2238), .B(n2302), .C(n18), .Y(n668) );
  OAI21X1 U1891 ( .A(n2238), .B(n2304), .C(n20), .Y(n669) );
  OAI21X1 U1892 ( .A(n2238), .B(n2306), .C(n22), .Y(n670) );
  OAI21X1 U1893 ( .A(n2238), .B(n2308), .C(n24), .Y(n671) );
  OAI21X1 U1894 ( .A(n2238), .B(n2310), .C(n26), .Y(n672) );
  OAI21X1 U1895 ( .A(n2238), .B(n2312), .C(n28), .Y(n673) );
  OAI21X1 U1896 ( .A(n2238), .B(n2314), .C(n30), .Y(n674) );
  OAI21X1 U1897 ( .A(n2239), .B(n2315), .C(n32), .Y(n675) );
  OAI21X1 U1898 ( .A(n2239), .B(n2318), .C(n34), .Y(n676) );
  OAI21X1 U1899 ( .A(n2239), .B(n2320), .C(n36), .Y(n677) );
  OAI21X1 U1900 ( .A(n2239), .B(n6), .C(n38), .Y(n678) );
  OAI21X1 U1901 ( .A(n2239), .B(n2325), .C(n40), .Y(n679) );
  OAI21X1 U1902 ( .A(n2239), .B(n2327), .C(n42), .Y(n680) );
  OAI21X1 U1903 ( .A(n2239), .B(n2328), .C(n44), .Y(n681) );
  OAI21X1 U1904 ( .A(n2239), .B(n2331), .C(n46), .Y(n682) );
  NAND3X1 U1905 ( .A(n2334), .B(n2185), .C(n2337), .Y(n2360) );
  OAI21X1 U1906 ( .A(n2299), .B(n2240), .C(n48), .Y(n683) );
  OAI21X1 U1907 ( .A(n2240), .B(n2301), .C(n50), .Y(n684) );
  OAI21X1 U1908 ( .A(n2240), .B(n2303), .C(n52), .Y(n685) );
  OAI21X1 U1909 ( .A(n2240), .B(n2305), .C(n54), .Y(n686) );
  OAI21X1 U1910 ( .A(n2240), .B(n2307), .C(n56), .Y(n687) );
  OAI21X1 U1911 ( .A(n2240), .B(n2309), .C(n58), .Y(n688) );
  OAI21X1 U1912 ( .A(n2240), .B(n2311), .C(n60), .Y(n689) );
  OAI21X1 U1913 ( .A(n2240), .B(n2313), .C(n62), .Y(n690) );
  OAI21X1 U1914 ( .A(n2241), .B(n2316), .C(n64), .Y(n691) );
  OAI21X1 U1915 ( .A(n2241), .B(n2317), .C(n66), .Y(n692) );
  OAI21X1 U1916 ( .A(n2241), .B(n2320), .C(n68), .Y(n693) );
  OAI21X1 U1917 ( .A(n2241), .B(n2321), .C(n70), .Y(n694) );
  OAI21X1 U1918 ( .A(n2241), .B(n2325), .C(n72), .Y(n695) );
  OAI21X1 U1919 ( .A(n2241), .B(n2326), .C(n74), .Y(n696) );
  OAI21X1 U1920 ( .A(n2241), .B(n2329), .C(n76), .Y(n697) );
  OAI21X1 U1921 ( .A(n2241), .B(n2330), .C(n78), .Y(n698) );
  NAND3X1 U1922 ( .A(n2185), .B(n2337), .C(n2335), .Y(n2361) );
  OAI21X1 U1923 ( .A(n2243), .B(n2299), .C(n80), .Y(n699) );
  OAI21X1 U1924 ( .A(n2243), .B(n2302), .C(n82), .Y(n700) );
  OAI21X1 U1925 ( .A(n2243), .B(n2304), .C(n84), .Y(n701) );
  OAI21X1 U1926 ( .A(n2243), .B(n2306), .C(n86), .Y(n702) );
  OAI21X1 U1927 ( .A(n2243), .B(n2308), .C(n88), .Y(n703) );
  OAI21X1 U1928 ( .A(n2243), .B(n2310), .C(n90), .Y(n704) );
  OAI21X1 U1929 ( .A(n2243), .B(n2312), .C(n92), .Y(n705) );
  OAI21X1 U1930 ( .A(n2243), .B(n2314), .C(n94), .Y(n706) );
  OAI21X1 U1931 ( .A(n2244), .B(n2315), .C(n96), .Y(n707) );
  OAI21X1 U1932 ( .A(n2244), .B(n2317), .C(n98), .Y(n708) );
  OAI21X1 U1933 ( .A(n2244), .B(n2319), .C(n100), .Y(n709) );
  OAI21X1 U1934 ( .A(n2244), .B(n2322), .C(n102), .Y(n710) );
  OAI21X1 U1935 ( .A(n2244), .B(n2324), .C(n104), .Y(n711) );
  OAI21X1 U1936 ( .A(n2244), .B(n2326), .C(n106), .Y(n712) );
  OAI21X1 U1937 ( .A(n2244), .B(n2328), .C(n108), .Y(n713) );
  OAI21X1 U1938 ( .A(n2244), .B(n2330), .C(n110), .Y(n714) );
  NAND3X1 U1939 ( .A(n2334), .B(n2336), .C(n2338), .Y(n2362) );
  OAI21X1 U1940 ( .A(n2245), .B(n2299), .C(n112), .Y(n715) );
  OAI21X1 U1941 ( .A(n2245), .B(n2301), .C(n114), .Y(n716) );
  OAI21X1 U1942 ( .A(n2245), .B(n2303), .C(n116), .Y(n717) );
  OAI21X1 U1943 ( .A(n2245), .B(n2305), .C(n118), .Y(n718) );
  OAI21X1 U1944 ( .A(n2245), .B(n2307), .C(n120), .Y(n719) );
  OAI21X1 U1945 ( .A(n2245), .B(n2309), .C(n122), .Y(n720) );
  OAI21X1 U1946 ( .A(n2245), .B(n2311), .C(n124), .Y(n721) );
  OAI21X1 U1947 ( .A(n2245), .B(n2313), .C(n126), .Y(n722) );
  OAI21X1 U1948 ( .A(n2246), .B(n2316), .C(n128), .Y(n723) );
  OAI21X1 U1949 ( .A(n2246), .B(n2317), .C(n130), .Y(n724) );
  OAI21X1 U1950 ( .A(n2246), .B(n2319), .C(n132), .Y(n725) );
  OAI21X1 U1951 ( .A(n2246), .B(n2321), .C(n134), .Y(n726) );
  OAI21X1 U1952 ( .A(n2246), .B(n2324), .C(n136), .Y(n727) );
  OAI21X1 U1953 ( .A(n2246), .B(n2327), .C(n138), .Y(n728) );
  OAI21X1 U1954 ( .A(n2246), .B(n2329), .C(n140), .Y(n729) );
  OAI21X1 U1955 ( .A(n2246), .B(n7), .C(n142), .Y(n730) );
  NAND3X1 U1956 ( .A(n2338), .B(n2336), .C(n2335), .Y(n2363) );
  NAND2X1 U1957 ( .A(\mem<26><0> ), .B(n626), .Y(n2364) );
  OAI21X1 U1958 ( .A(n2247), .B(n2299), .C(n2364), .Y(n731) );
  NAND2X1 U1959 ( .A(\mem<26><1> ), .B(n626), .Y(n2365) );
  OAI21X1 U1960 ( .A(n2247), .B(n2302), .C(n2365), .Y(n732) );
  NAND2X1 U1961 ( .A(\mem<26><2> ), .B(n626), .Y(n2366) );
  OAI21X1 U1962 ( .A(n2247), .B(n2304), .C(n2366), .Y(n733) );
  NAND2X1 U1963 ( .A(\mem<26><3> ), .B(n626), .Y(n2367) );
  OAI21X1 U1964 ( .A(n2247), .B(n2306), .C(n2367), .Y(n734) );
  NAND2X1 U1965 ( .A(\mem<26><4> ), .B(n626), .Y(n2368) );
  OAI21X1 U1966 ( .A(n2247), .B(n2308), .C(n2368), .Y(n735) );
  NAND2X1 U1967 ( .A(\mem<26><5> ), .B(n626), .Y(n2369) );
  OAI21X1 U1968 ( .A(n2247), .B(n2310), .C(n2369), .Y(n736) );
  NAND2X1 U1969 ( .A(\mem<26><6> ), .B(n626), .Y(n2370) );
  OAI21X1 U1970 ( .A(n2247), .B(n2312), .C(n2370), .Y(n737) );
  NAND2X1 U1971 ( .A(\mem<26><7> ), .B(n626), .Y(n2371) );
  OAI21X1 U1972 ( .A(n2247), .B(n2314), .C(n2371), .Y(n738) );
  OAI21X1 U1973 ( .A(n2248), .B(n2315), .C(n144), .Y(n739) );
  OAI21X1 U1974 ( .A(n2248), .B(n2317), .C(n146), .Y(n740) );
  OAI21X1 U1975 ( .A(n2248), .B(n2319), .C(n148), .Y(n741) );
  OAI21X1 U1976 ( .A(n2248), .B(n2322), .C(n150), .Y(n742) );
  OAI21X1 U1977 ( .A(n2248), .B(n2324), .C(n152), .Y(n743) );
  OAI21X1 U1978 ( .A(n2248), .B(n2326), .C(n154), .Y(n744) );
  OAI21X1 U1979 ( .A(n2248), .B(n2328), .C(n156), .Y(n745) );
  OAI21X1 U1980 ( .A(n2248), .B(n2330), .C(n158), .Y(n746) );
  NAND3X1 U1981 ( .A(n2334), .B(n2338), .C(n2337), .Y(n2372) );
  NAND2X1 U1982 ( .A(\mem<25><0> ), .B(n628), .Y(n2373) );
  OAI21X1 U1983 ( .A(n2249), .B(n2299), .C(n2373), .Y(n747) );
  NAND2X1 U1984 ( .A(\mem<25><1> ), .B(n628), .Y(n2374) );
  OAI21X1 U1985 ( .A(n2249), .B(n2301), .C(n2374), .Y(n748) );
  NAND2X1 U1986 ( .A(\mem<25><2> ), .B(n628), .Y(n2375) );
  OAI21X1 U1987 ( .A(n2249), .B(n2303), .C(n2375), .Y(n749) );
  NAND2X1 U1988 ( .A(\mem<25><3> ), .B(n628), .Y(n2376) );
  OAI21X1 U1989 ( .A(n2249), .B(n2305), .C(n2376), .Y(n750) );
  NAND2X1 U1990 ( .A(\mem<25><4> ), .B(n628), .Y(n2377) );
  OAI21X1 U1991 ( .A(n2249), .B(n2307), .C(n2377), .Y(n751) );
  NAND2X1 U1992 ( .A(\mem<25><5> ), .B(n628), .Y(n2378) );
  OAI21X1 U1993 ( .A(n2249), .B(n2309), .C(n2378), .Y(n752) );
  NAND2X1 U1994 ( .A(\mem<25><6> ), .B(n628), .Y(n2379) );
  OAI21X1 U1995 ( .A(n2249), .B(n2311), .C(n2379), .Y(n753) );
  NAND2X1 U1996 ( .A(\mem<25><7> ), .B(n628), .Y(n2380) );
  OAI21X1 U1997 ( .A(n2249), .B(n2313), .C(n2380), .Y(n754) );
  OAI21X1 U1998 ( .A(n2250), .B(n2316), .C(n160), .Y(n755) );
  OAI21X1 U1999 ( .A(n2250), .B(n2317), .C(n162), .Y(n756) );
  OAI21X1 U2000 ( .A(n2250), .B(n2320), .C(n164), .Y(n757) );
  OAI21X1 U2001 ( .A(n2250), .B(n6), .C(n166), .Y(n758) );
  OAI21X1 U2002 ( .A(n2250), .B(n2325), .C(n168), .Y(n759) );
  OAI21X1 U2003 ( .A(n2250), .B(n2326), .C(n170), .Y(n760) );
  OAI21X1 U2004 ( .A(n2250), .B(n2329), .C(n172), .Y(n761) );
  OAI21X1 U2005 ( .A(n2250), .B(n7), .C(n174), .Y(n762) );
  NOR3X1 U2006 ( .A(n2334), .B(n2336), .C(n2185), .Y(n2422) );
  OAI21X1 U2007 ( .A(n2251), .B(n2299), .C(n176), .Y(n763) );
  OAI21X1 U2008 ( .A(n2251), .B(n2301), .C(n178), .Y(n764) );
  OAI21X1 U2009 ( .A(n2251), .B(n2303), .C(n180), .Y(n765) );
  OAI21X1 U2010 ( .A(n2251), .B(n2305), .C(n182), .Y(n766) );
  OAI21X1 U2011 ( .A(n2251), .B(n2307), .C(n184), .Y(n767) );
  OAI21X1 U2012 ( .A(n2251), .B(n2309), .C(n186), .Y(n768) );
  OAI21X1 U2013 ( .A(n2251), .B(n2311), .C(n188), .Y(n769) );
  OAI21X1 U2014 ( .A(n2251), .B(n2313), .C(n190), .Y(n770) );
  OAI21X1 U2015 ( .A(n2251), .B(n2315), .C(n192), .Y(n771) );
  OAI21X1 U2016 ( .A(n2251), .B(n2317), .C(n194), .Y(n772) );
  OAI21X1 U2017 ( .A(n2251), .B(n2319), .C(n196), .Y(n773) );
  OAI21X1 U2018 ( .A(n2251), .B(n2321), .C(n198), .Y(n774) );
  OAI21X1 U2019 ( .A(n2251), .B(n2324), .C(n200), .Y(n775) );
  OAI21X1 U2020 ( .A(n2251), .B(n2326), .C(n202), .Y(n776) );
  OAI21X1 U2021 ( .A(n2251), .B(n2328), .C(n204), .Y(n777) );
  OAI21X1 U2022 ( .A(n2251), .B(n2330), .C(n206), .Y(n778) );
  NAND2X1 U2023 ( .A(\mem<23><0> ), .B(n632), .Y(n2381) );
  OAI21X1 U2024 ( .A(n2252), .B(n2299), .C(n2381), .Y(n779) );
  NAND2X1 U2025 ( .A(\mem<23><1> ), .B(n632), .Y(n2382) );
  OAI21X1 U2026 ( .A(n2252), .B(n2302), .C(n2382), .Y(n780) );
  NAND2X1 U2027 ( .A(\mem<23><2> ), .B(n632), .Y(n2383) );
  OAI21X1 U2028 ( .A(n2252), .B(n2304), .C(n2383), .Y(n781) );
  NAND2X1 U2029 ( .A(\mem<23><3> ), .B(n632), .Y(n2384) );
  OAI21X1 U2030 ( .A(n2252), .B(n2306), .C(n2384), .Y(n782) );
  NAND2X1 U2031 ( .A(\mem<23><4> ), .B(n632), .Y(n2385) );
  OAI21X1 U2032 ( .A(n2252), .B(n2308), .C(n2385), .Y(n783) );
  NAND2X1 U2033 ( .A(\mem<23><5> ), .B(n632), .Y(n2386) );
  OAI21X1 U2034 ( .A(n2252), .B(n2310), .C(n2386), .Y(n784) );
  NAND2X1 U2035 ( .A(\mem<23><6> ), .B(n632), .Y(n2387) );
  OAI21X1 U2036 ( .A(n2252), .B(n2312), .C(n2387), .Y(n785) );
  NAND2X1 U2037 ( .A(\mem<23><7> ), .B(n632), .Y(n2388) );
  OAI21X1 U2038 ( .A(n2252), .B(n2314), .C(n2388), .Y(n786) );
  OAI21X1 U2039 ( .A(n2253), .B(n2316), .C(n208), .Y(n787) );
  OAI21X1 U2040 ( .A(n2253), .B(n2318), .C(n210), .Y(n788) );
  OAI21X1 U2041 ( .A(n2253), .B(n2319), .C(n212), .Y(n789) );
  OAI21X1 U2042 ( .A(n2253), .B(n2321), .C(n215), .Y(n790) );
  OAI21X1 U2043 ( .A(n2253), .B(n2325), .C(n217), .Y(n791) );
  OAI21X1 U2044 ( .A(n2253), .B(n2327), .C(n219), .Y(n792) );
  OAI21X1 U2045 ( .A(n2253), .B(n2329), .C(n221), .Y(n793) );
  OAI21X1 U2046 ( .A(n2253), .B(n2331), .C(n223), .Y(n794) );
  NAND2X1 U2047 ( .A(\mem<22><0> ), .B(n635), .Y(n2389) );
  OAI21X1 U2048 ( .A(n2254), .B(n2299), .C(n2389), .Y(n795) );
  NAND2X1 U2049 ( .A(\mem<22><1> ), .B(n635), .Y(n2390) );
  OAI21X1 U2050 ( .A(n2254), .B(n2302), .C(n2390), .Y(n796) );
  NAND2X1 U2051 ( .A(\mem<22><2> ), .B(n635), .Y(n2391) );
  OAI21X1 U2052 ( .A(n2254), .B(n2304), .C(n2391), .Y(n797) );
  NAND2X1 U2053 ( .A(\mem<22><3> ), .B(n635), .Y(n2392) );
  OAI21X1 U2054 ( .A(n2254), .B(n2306), .C(n2392), .Y(n798) );
  NAND2X1 U2055 ( .A(\mem<22><4> ), .B(n635), .Y(n2393) );
  OAI21X1 U2056 ( .A(n2254), .B(n2308), .C(n2393), .Y(n799) );
  NAND2X1 U2057 ( .A(\mem<22><5> ), .B(n635), .Y(n2394) );
  OAI21X1 U2058 ( .A(n2254), .B(n2310), .C(n2394), .Y(n800) );
  NAND2X1 U2059 ( .A(\mem<22><6> ), .B(n635), .Y(n2395) );
  OAI21X1 U2060 ( .A(n2254), .B(n2312), .C(n2395), .Y(n801) );
  NAND2X1 U2061 ( .A(\mem<22><7> ), .B(n635), .Y(n2396) );
  OAI21X1 U2062 ( .A(n2254), .B(n2314), .C(n2396), .Y(n802) );
  OAI21X1 U2063 ( .A(n2255), .B(n2316), .C(n225), .Y(n803) );
  OAI21X1 U2064 ( .A(n2255), .B(n2318), .C(n227), .Y(n804) );
  OAI21X1 U2065 ( .A(n2255), .B(n2319), .C(n229), .Y(n805) );
  OAI21X1 U2066 ( .A(n2255), .B(n6), .C(n231), .Y(n806) );
  OAI21X1 U2067 ( .A(n2255), .B(n2324), .C(n233), .Y(n807) );
  OAI21X1 U2068 ( .A(n2255), .B(n2327), .C(n235), .Y(n808) );
  OAI21X1 U2069 ( .A(n2255), .B(n2329), .C(n237), .Y(n809) );
  OAI21X1 U2070 ( .A(n2255), .B(n2331), .C(n239), .Y(n810) );
  NAND2X1 U2071 ( .A(\mem<21><0> ), .B(n638), .Y(n2397) );
  OAI21X1 U2072 ( .A(n2256), .B(n2299), .C(n2397), .Y(n811) );
  NAND2X1 U2073 ( .A(\mem<21><1> ), .B(n638), .Y(n2398) );
  OAI21X1 U2074 ( .A(n2256), .B(n2302), .C(n2398), .Y(n812) );
  NAND2X1 U2075 ( .A(\mem<21><2> ), .B(n638), .Y(n2399) );
  OAI21X1 U2076 ( .A(n2256), .B(n2304), .C(n2399), .Y(n813) );
  NAND2X1 U2077 ( .A(\mem<21><3> ), .B(n638), .Y(n2400) );
  OAI21X1 U2078 ( .A(n2256), .B(n2306), .C(n2400), .Y(n814) );
  NAND2X1 U2079 ( .A(\mem<21><4> ), .B(n638), .Y(n2401) );
  OAI21X1 U2080 ( .A(n2256), .B(n2308), .C(n2401), .Y(n815) );
  NAND2X1 U2081 ( .A(\mem<21><5> ), .B(n638), .Y(n2402) );
  OAI21X1 U2082 ( .A(n2256), .B(n2310), .C(n2402), .Y(n816) );
  NAND2X1 U2083 ( .A(\mem<21><6> ), .B(n638), .Y(n2403) );
  OAI21X1 U2084 ( .A(n2256), .B(n2312), .C(n2403), .Y(n817) );
  NAND2X1 U2085 ( .A(\mem<21><7> ), .B(n638), .Y(n2404) );
  OAI21X1 U2086 ( .A(n2256), .B(n2314), .C(n2404), .Y(n818) );
  OAI21X1 U2087 ( .A(n2257), .B(n2316), .C(n241), .Y(n819) );
  OAI21X1 U2088 ( .A(n2257), .B(n2317), .C(n243), .Y(n820) );
  OAI21X1 U2089 ( .A(n2257), .B(n2320), .C(n245), .Y(n821) );
  OAI21X1 U2090 ( .A(n2257), .B(n6), .C(n247), .Y(n822) );
  OAI21X1 U2091 ( .A(n2257), .B(n2325), .C(n249), .Y(n823) );
  OAI21X1 U2092 ( .A(n2257), .B(n2326), .C(n251), .Y(n824) );
  OAI21X1 U2093 ( .A(n2257), .B(n2329), .C(n253), .Y(n825) );
  OAI21X1 U2094 ( .A(n2257), .B(n2330), .C(n255), .Y(n826) );
  NAND2X1 U2095 ( .A(\mem<20><0> ), .B(n641), .Y(n2405) );
  OAI21X1 U2096 ( .A(n2258), .B(n2299), .C(n2405), .Y(n827) );
  NAND2X1 U2097 ( .A(\mem<20><1> ), .B(n641), .Y(n2406) );
  OAI21X1 U2098 ( .A(n2258), .B(n2302), .C(n2406), .Y(n828) );
  NAND2X1 U2099 ( .A(\mem<20><2> ), .B(n641), .Y(n2407) );
  OAI21X1 U2100 ( .A(n2258), .B(n2304), .C(n2407), .Y(n829) );
  NAND2X1 U2101 ( .A(\mem<20><3> ), .B(n641), .Y(n2408) );
  OAI21X1 U2102 ( .A(n2258), .B(n2306), .C(n2408), .Y(n830) );
  NAND2X1 U2103 ( .A(\mem<20><4> ), .B(n641), .Y(n2409) );
  OAI21X1 U2104 ( .A(n2258), .B(n2308), .C(n2409), .Y(n831) );
  NAND2X1 U2105 ( .A(\mem<20><5> ), .B(n641), .Y(n2410) );
  OAI21X1 U2106 ( .A(n2258), .B(n2310), .C(n2410), .Y(n832) );
  NAND2X1 U2107 ( .A(\mem<20><6> ), .B(n641), .Y(n2411) );
  OAI21X1 U2108 ( .A(n2258), .B(n2312), .C(n2411), .Y(n833) );
  NAND2X1 U2109 ( .A(\mem<20><7> ), .B(n641), .Y(n2412) );
  OAI21X1 U2110 ( .A(n2258), .B(n2314), .C(n2412), .Y(n834) );
  OAI21X1 U2111 ( .A(n2259), .B(n2316), .C(n257), .Y(n835) );
  OAI21X1 U2112 ( .A(n2259), .B(n2317), .C(n259), .Y(n836) );
  OAI21X1 U2113 ( .A(n2259), .B(n2319), .C(n261), .Y(n837) );
  OAI21X1 U2114 ( .A(n2259), .B(n6), .C(n263), .Y(n838) );
  OAI21X1 U2115 ( .A(n2259), .B(n2324), .C(n265), .Y(n839) );
  OAI21X1 U2116 ( .A(n2259), .B(n2326), .C(n267), .Y(n840) );
  OAI21X1 U2117 ( .A(n2259), .B(n2329), .C(n269), .Y(n841) );
  OAI21X1 U2118 ( .A(n2259), .B(n2330), .C(n271), .Y(n842) );
  OAI21X1 U2119 ( .A(n2260), .B(n2299), .C(n353), .Y(n843) );
  OAI21X1 U2120 ( .A(n2260), .B(n2302), .C(n355), .Y(n844) );
  OAI21X1 U2121 ( .A(n2260), .B(n2304), .C(n357), .Y(n845) );
  OAI21X1 U2122 ( .A(n2260), .B(n2306), .C(n359), .Y(n846) );
  OAI21X1 U2123 ( .A(n2260), .B(n2308), .C(n361), .Y(n847) );
  OAI21X1 U2124 ( .A(n2260), .B(n2310), .C(n363), .Y(n848) );
  OAI21X1 U2125 ( .A(n2260), .B(n2312), .C(n365), .Y(n849) );
  OAI21X1 U2126 ( .A(n2260), .B(n2314), .C(n367), .Y(n850) );
  OAI21X1 U2127 ( .A(n2261), .B(n2316), .C(n369), .Y(n851) );
  OAI21X1 U2128 ( .A(n2261), .B(n2317), .C(n371), .Y(n852) );
  OAI21X1 U2129 ( .A(n2261), .B(n2319), .C(n373), .Y(n853) );
  OAI21X1 U2130 ( .A(n2261), .B(n2321), .C(n1207), .Y(n854) );
  OAI21X1 U2131 ( .A(n2261), .B(n2324), .C(n1209), .Y(n855) );
  OAI21X1 U2132 ( .A(n2261), .B(n2326), .C(n1211), .Y(n856) );
  OAI21X1 U2133 ( .A(n2261), .B(n2329), .C(n1213), .Y(n857) );
  OAI21X1 U2134 ( .A(n2261), .B(n7), .C(n1215), .Y(n858) );
  OAI21X1 U2135 ( .A(n2262), .B(n2300), .C(n375), .Y(n859) );
  OAI21X1 U2136 ( .A(n2262), .B(n2302), .C(n377), .Y(n860) );
  OAI21X1 U2137 ( .A(n2262), .B(n2304), .C(n379), .Y(n861) );
  OAI21X1 U2138 ( .A(n2262), .B(n2306), .C(n381), .Y(n862) );
  OAI21X1 U2139 ( .A(n2262), .B(n2308), .C(n383), .Y(n863) );
  OAI21X1 U2140 ( .A(n2262), .B(n2310), .C(n385), .Y(n864) );
  OAI21X1 U2141 ( .A(n2262), .B(n2312), .C(n387), .Y(n865) );
  OAI21X1 U2142 ( .A(n2262), .B(n2314), .C(n389), .Y(n866) );
  OAI21X1 U2143 ( .A(n2263), .B(n2316), .C(n391), .Y(n867) );
  OAI21X1 U2144 ( .A(n2263), .B(n2318), .C(n393), .Y(n868) );
  OAI21X1 U2145 ( .A(n2263), .B(n2320), .C(n395), .Y(n869) );
  OAI21X1 U2146 ( .A(n2263), .B(n6), .C(n1217), .Y(n870) );
  OAI21X1 U2147 ( .A(n2263), .B(n2325), .C(n1219), .Y(n871) );
  OAI21X1 U2148 ( .A(n2263), .B(n2327), .C(n1221), .Y(n872) );
  OAI21X1 U2149 ( .A(n2263), .B(n2329), .C(n1223), .Y(n873) );
  OAI21X1 U2150 ( .A(n2263), .B(n7), .C(n1225), .Y(n874) );
  OAI21X1 U2151 ( .A(n2264), .B(n2299), .C(n397), .Y(n875) );
  OAI21X1 U2152 ( .A(n2264), .B(n2302), .C(n399), .Y(n876) );
  OAI21X1 U2153 ( .A(n2264), .B(n2304), .C(n401), .Y(n877) );
  OAI21X1 U2154 ( .A(n2264), .B(n2306), .C(n403), .Y(n878) );
  OAI21X1 U2155 ( .A(n2264), .B(n2308), .C(n405), .Y(n879) );
  OAI21X1 U2156 ( .A(n2264), .B(n2310), .C(n407), .Y(n880) );
  OAI21X1 U2157 ( .A(n2264), .B(n2312), .C(n409), .Y(n881) );
  OAI21X1 U2158 ( .A(n2264), .B(n2314), .C(n411), .Y(n882) );
  OAI21X1 U2159 ( .A(n2265), .B(n2316), .C(n413), .Y(n883) );
  OAI21X1 U2160 ( .A(n2265), .B(n2318), .C(n415), .Y(n884) );
  OAI21X1 U2161 ( .A(n2265), .B(n2320), .C(n417), .Y(n885) );
  OAI21X1 U2162 ( .A(n2265), .B(n6), .C(n1227), .Y(n886) );
  OAI21X1 U2163 ( .A(n2265), .B(n2324), .C(n1229), .Y(n887) );
  OAI21X1 U2164 ( .A(n2265), .B(n2327), .C(n1231), .Y(n888) );
  OAI21X1 U2165 ( .A(n2265), .B(n2329), .C(n1233), .Y(n889) );
  OAI21X1 U2166 ( .A(n2265), .B(n2331), .C(n1235), .Y(n890) );
  OAI21X1 U2167 ( .A(n2267), .B(n2300), .C(n419), .Y(n891) );
  OAI21X1 U2168 ( .A(n2267), .B(n2302), .C(n421), .Y(n892) );
  OAI21X1 U2169 ( .A(n2267), .B(n2304), .C(n423), .Y(n893) );
  OAI21X1 U2170 ( .A(n2267), .B(n2306), .C(n425), .Y(n894) );
  OAI21X1 U2171 ( .A(n2267), .B(n2308), .C(n427), .Y(n895) );
  OAI21X1 U2172 ( .A(n2267), .B(n2310), .C(n429), .Y(n896) );
  OAI21X1 U2173 ( .A(n2267), .B(n2312), .C(n431), .Y(n897) );
  OAI21X1 U2174 ( .A(n2267), .B(n2314), .C(n433), .Y(n898) );
  OAI21X1 U2175 ( .A(n2267), .B(n2316), .C(n435), .Y(n899) );
  OAI21X1 U2176 ( .A(n2267), .B(n2318), .C(n437), .Y(n900) );
  OAI21X1 U2177 ( .A(n2267), .B(n2320), .C(n439), .Y(n901) );
  OAI21X1 U2178 ( .A(n2267), .B(n5), .C(n1237), .Y(n902) );
  OAI21X1 U2179 ( .A(n2267), .B(n2325), .C(n1239), .Y(n903) );
  OAI21X1 U2180 ( .A(n2267), .B(n2327), .C(n1241), .Y(n904) );
  OAI21X1 U2181 ( .A(n2267), .B(n2329), .C(n1243), .Y(n905) );
  OAI21X1 U2182 ( .A(n2267), .B(n2331), .C(n1245), .Y(n906) );
  NAND3X1 U2183 ( .A(n2339), .B(n214), .C(n2342), .Y(n2413) );
  OAI21X1 U2184 ( .A(n2268), .B(n2300), .C(n441), .Y(n907) );
  OAI21X1 U2185 ( .A(n2268), .B(n2302), .C(n443), .Y(n908) );
  OAI21X1 U2186 ( .A(n2268), .B(n2304), .C(n445), .Y(n909) );
  OAI21X1 U2187 ( .A(n2268), .B(n2306), .C(n447), .Y(n910) );
  OAI21X1 U2188 ( .A(n2268), .B(n2308), .C(n449), .Y(n911) );
  OAI21X1 U2189 ( .A(n2268), .B(n2310), .C(n451), .Y(n912) );
  OAI21X1 U2190 ( .A(n2268), .B(n2312), .C(n453), .Y(n913) );
  OAI21X1 U2191 ( .A(n2268), .B(n2314), .C(n455), .Y(n914) );
  OAI21X1 U2192 ( .A(n2269), .B(n2316), .C(n457), .Y(n915) );
  OAI21X1 U2193 ( .A(n2269), .B(n2318), .C(n459), .Y(n916) );
  OAI21X1 U2194 ( .A(n2269), .B(n2319), .C(n461), .Y(n917) );
  OAI21X1 U2195 ( .A(n2269), .B(n2321), .C(n1247), .Y(n918) );
  OAI21X1 U2196 ( .A(n2269), .B(n2324), .C(n1249), .Y(n919) );
  OAI21X1 U2197 ( .A(n2269), .B(n2327), .C(n1251), .Y(n920) );
  OAI21X1 U2198 ( .A(n2269), .B(n2329), .C(n1253), .Y(n921) );
  OAI21X1 U2199 ( .A(n2269), .B(n2331), .C(n1255), .Y(n922) );
  OAI21X1 U2200 ( .A(n2270), .B(n2299), .C(n463), .Y(n923) );
  OAI21X1 U2201 ( .A(n2270), .B(n2302), .C(n465), .Y(n924) );
  OAI21X1 U2202 ( .A(n2270), .B(n2304), .C(n467), .Y(n925) );
  OAI21X1 U2203 ( .A(n2270), .B(n2306), .C(n469), .Y(n926) );
  OAI21X1 U2204 ( .A(n2270), .B(n2308), .C(n471), .Y(n927) );
  OAI21X1 U2205 ( .A(n2270), .B(n2310), .C(n473), .Y(n928) );
  OAI21X1 U2206 ( .A(n2270), .B(n2312), .C(n475), .Y(n929) );
  OAI21X1 U2207 ( .A(n2270), .B(n2314), .C(n477), .Y(n930) );
  OAI21X1 U2208 ( .A(n2271), .B(n2316), .C(n479), .Y(n931) );
  OAI21X1 U2209 ( .A(n2271), .B(n2317), .C(n481), .Y(n932) );
  OAI21X1 U2210 ( .A(n2271), .B(n2320), .C(n483), .Y(n933) );
  OAI21X1 U2211 ( .A(n2271), .B(n6), .C(n1257), .Y(n934) );
  OAI21X1 U2212 ( .A(n2271), .B(n2325), .C(n1259), .Y(n935) );
  OAI21X1 U2213 ( .A(n2271), .B(n2326), .C(n1261), .Y(n936) );
  OAI21X1 U2214 ( .A(n2271), .B(n2329), .C(n1263), .Y(n937) );
  OAI21X1 U2215 ( .A(n2271), .B(n2330), .C(n1265), .Y(n938) );
  OAI21X1 U2216 ( .A(n2272), .B(n2300), .C(n485), .Y(n939) );
  OAI21X1 U2217 ( .A(n2272), .B(n2302), .C(n487), .Y(n940) );
  OAI21X1 U2218 ( .A(n2272), .B(n2304), .C(n489), .Y(n941) );
  OAI21X1 U2219 ( .A(n2272), .B(n2306), .C(n491), .Y(n942) );
  OAI21X1 U2220 ( .A(n2272), .B(n2308), .C(n493), .Y(n943) );
  OAI21X1 U2221 ( .A(n2272), .B(n2310), .C(n495), .Y(n944) );
  OAI21X1 U2222 ( .A(n2272), .B(n2312), .C(n497), .Y(n945) );
  OAI21X1 U2223 ( .A(n2272), .B(n2314), .C(n499), .Y(n946) );
  OAI21X1 U2224 ( .A(n2273), .B(n2316), .C(n501), .Y(n947) );
  OAI21X1 U2225 ( .A(n2273), .B(n2317), .C(n503), .Y(n948) );
  OAI21X1 U2226 ( .A(n2273), .B(n2320), .C(n505), .Y(n949) );
  OAI21X1 U2227 ( .A(n2273), .B(n2321), .C(n1267), .Y(n950) );
  OAI21X1 U2228 ( .A(n2273), .B(n2325), .C(n1269), .Y(n951) );
  OAI21X1 U2229 ( .A(n2273), .B(n2326), .C(n1271), .Y(n952) );
  OAI21X1 U2230 ( .A(n2273), .B(n2329), .C(n1273), .Y(n953) );
  OAI21X1 U2231 ( .A(n2273), .B(n2330), .C(n1275), .Y(n954) );
  OAI21X1 U2232 ( .A(n2274), .B(n2299), .C(n507), .Y(n955) );
  OAI21X1 U2233 ( .A(n2274), .B(n2302), .C(n509), .Y(n956) );
  OAI21X1 U2234 ( .A(n2274), .B(n2304), .C(n511), .Y(n957) );
  OAI21X1 U2235 ( .A(n2274), .B(n2306), .C(n513), .Y(n958) );
  OAI21X1 U2236 ( .A(n2274), .B(n2308), .C(n515), .Y(n959) );
  OAI21X1 U2237 ( .A(n2274), .B(n2310), .C(n517), .Y(n960) );
  OAI21X1 U2238 ( .A(n2274), .B(n2312), .C(n519), .Y(n961) );
  OAI21X1 U2239 ( .A(n2274), .B(n2314), .C(n521), .Y(n962) );
  OAI21X1 U2240 ( .A(n2275), .B(n2316), .C(n523), .Y(n963) );
  OAI21X1 U2241 ( .A(n2275), .B(n2318), .C(n525), .Y(n964) );
  OAI21X1 U2242 ( .A(n2275), .B(n2319), .C(n527), .Y(n965) );
  OAI21X1 U2243 ( .A(n2275), .B(n5), .C(n1277), .Y(n966) );
  OAI21X1 U2244 ( .A(n2275), .B(n2324), .C(n1279), .Y(n967) );
  OAI21X1 U2245 ( .A(n2275), .B(n2327), .C(n1281), .Y(n968) );
  OAI21X1 U2246 ( .A(n2275), .B(n2329), .C(n1283), .Y(n969) );
  OAI21X1 U2247 ( .A(n2275), .B(n7), .C(n1285), .Y(n970) );
  OAI21X1 U2248 ( .A(n2276), .B(n2300), .C(n529), .Y(n971) );
  OAI21X1 U2249 ( .A(n2276), .B(n2301), .C(n531), .Y(n972) );
  OAI21X1 U2250 ( .A(n2276), .B(n2303), .C(n533), .Y(n973) );
  OAI21X1 U2251 ( .A(n2276), .B(n2305), .C(n535), .Y(n974) );
  OAI21X1 U2252 ( .A(n2276), .B(n2307), .C(n537), .Y(n975) );
  OAI21X1 U2253 ( .A(n2276), .B(n2309), .C(n539), .Y(n976) );
  OAI21X1 U2254 ( .A(n2276), .B(n2311), .C(n541), .Y(n977) );
  OAI21X1 U2255 ( .A(n2276), .B(n2313), .C(n543), .Y(n978) );
  OAI21X1 U2256 ( .A(n2277), .B(n2315), .C(n545), .Y(n979) );
  OAI21X1 U2257 ( .A(n2277), .B(n2318), .C(n547), .Y(n980) );
  OAI21X1 U2258 ( .A(n2277), .B(n2320), .C(n549), .Y(n981) );
  OAI21X1 U2259 ( .A(n2277), .B(n2322), .C(n1287), .Y(n982) );
  OAI21X1 U2260 ( .A(n2277), .B(n2324), .C(n1289), .Y(n983) );
  OAI21X1 U2261 ( .A(n2277), .B(n2326), .C(n1291), .Y(n984) );
  OAI21X1 U2262 ( .A(n2277), .B(n2328), .C(n1293), .Y(n985) );
  OAI21X1 U2263 ( .A(n2277), .B(n7), .C(n1295), .Y(n986) );
  OAI21X1 U2264 ( .A(n2278), .B(n2300), .C(n551), .Y(n987) );
  OAI21X1 U2265 ( .A(n2278), .B(n2301), .C(n553), .Y(n988) );
  OAI21X1 U2266 ( .A(n2278), .B(n2303), .C(n555), .Y(n989) );
  OAI21X1 U2267 ( .A(n2278), .B(n2305), .C(n557), .Y(n990) );
  OAI21X1 U2268 ( .A(n2278), .B(n2307), .C(n559), .Y(n991) );
  OAI21X1 U2269 ( .A(n2278), .B(n2309), .C(n561), .Y(n992) );
  OAI21X1 U2270 ( .A(n2278), .B(n2311), .C(n563), .Y(n993) );
  OAI21X1 U2271 ( .A(n2278), .B(n2313), .C(n565), .Y(n994) );
  OAI21X1 U2272 ( .A(n2279), .B(n2315), .C(n567), .Y(n995) );
  OAI21X1 U2273 ( .A(n2279), .B(n2318), .C(n569), .Y(n996) );
  OAI21X1 U2274 ( .A(n2279), .B(n2320), .C(n571), .Y(n997) );
  OAI21X1 U2275 ( .A(n2279), .B(n2322), .C(n1297), .Y(n998) );
  OAI21X1 U2276 ( .A(n2279), .B(n2325), .C(n1299), .Y(n999) );
  OAI21X1 U2277 ( .A(n2279), .B(n2326), .C(n1301), .Y(n1000) );
  OAI21X1 U2278 ( .A(n2279), .B(n2328), .C(n1303), .Y(n1001) );
  OAI21X1 U2279 ( .A(n2279), .B(n7), .C(n1305), .Y(n1002) );
  OAI21X1 U2280 ( .A(n2280), .B(n2300), .C(n573), .Y(n1003) );
  OAI21X1 U2281 ( .A(n2280), .B(n2301), .C(n575), .Y(n1004) );
  OAI21X1 U2282 ( .A(n2280), .B(n2303), .C(n577), .Y(n1005) );
  OAI21X1 U2283 ( .A(n2280), .B(n2305), .C(n579), .Y(n1006) );
  OAI21X1 U2284 ( .A(n2280), .B(n2307), .C(n581), .Y(n1007) );
  OAI21X1 U2285 ( .A(n2280), .B(n2309), .C(n583), .Y(n1008) );
  OAI21X1 U2286 ( .A(n2280), .B(n2311), .C(n585), .Y(n1009) );
  OAI21X1 U2287 ( .A(n2280), .B(n2313), .C(n587), .Y(n1010) );
  OAI21X1 U2288 ( .A(n2281), .B(n2315), .C(n589), .Y(n1011) );
  OAI21X1 U2289 ( .A(n2281), .B(n2318), .C(n591), .Y(n1012) );
  OAI21X1 U2290 ( .A(n2281), .B(n2320), .C(n593), .Y(n1013) );
  OAI21X1 U2291 ( .A(n2281), .B(n2322), .C(n1307), .Y(n1014) );
  OAI21X1 U2292 ( .A(n2281), .B(n2325), .C(n1309), .Y(n1015) );
  OAI21X1 U2293 ( .A(n2281), .B(n2327), .C(n1311), .Y(n1016) );
  OAI21X1 U2294 ( .A(n2281), .B(n2328), .C(n1313), .Y(n1017) );
  OAI21X1 U2295 ( .A(n2281), .B(n2331), .C(n1315), .Y(n1018) );
  OAI21X1 U2296 ( .A(n2282), .B(n2300), .C(n1317), .Y(n1019) );
  OAI21X1 U2297 ( .A(n2282), .B(n2301), .C(n1319), .Y(n1020) );
  OAI21X1 U2298 ( .A(n2282), .B(n2303), .C(n1321), .Y(n1021) );
  OAI21X1 U2299 ( .A(n2282), .B(n2305), .C(n1323), .Y(n1022) );
  OAI21X1 U2300 ( .A(n2282), .B(n2307), .C(n1325), .Y(n1023) );
  OAI21X1 U2301 ( .A(n2282), .B(n2309), .C(n1327), .Y(n1024) );
  OAI21X1 U2302 ( .A(n2282), .B(n2311), .C(n1329), .Y(n1025) );
  OAI21X1 U2303 ( .A(n2282), .B(n2313), .C(n1331), .Y(n1026) );
  OAI21X1 U2304 ( .A(n2282), .B(n2315), .C(n1333), .Y(n1027) );
  OAI21X1 U2305 ( .A(n2282), .B(n2318), .C(n1335), .Y(n1028) );
  OAI21X1 U2306 ( .A(n2282), .B(n2319), .C(n1337), .Y(n1029) );
  OAI21X1 U2307 ( .A(n2282), .B(n2321), .C(n1505), .Y(n1030) );
  OAI21X1 U2308 ( .A(n2282), .B(n2324), .C(n1507), .Y(n1031) );
  OAI21X1 U2309 ( .A(n2282), .B(n2327), .C(n1509), .Y(n1032) );
  OAI21X1 U2310 ( .A(n2282), .B(n2328), .C(n1511), .Y(n1033) );
  OAI21X1 U2311 ( .A(n2282), .B(n2331), .C(n1513), .Y(n1034) );
  NAND3X1 U2312 ( .A(n2340), .B(n214), .C(n2342), .Y(n2415) );
  OAI21X1 U2313 ( .A(n2283), .B(n2300), .C(n1339), .Y(n1035) );
  OAI21X1 U2314 ( .A(n2283), .B(n2301), .C(n1341), .Y(n1036) );
  OAI21X1 U2315 ( .A(n2283), .B(n2303), .C(n1343), .Y(n1037) );
  OAI21X1 U2316 ( .A(n2283), .B(n2305), .C(n1345), .Y(n1038) );
  OAI21X1 U2317 ( .A(n2283), .B(n2307), .C(n1347), .Y(n1039) );
  OAI21X1 U2318 ( .A(n2283), .B(n2309), .C(n1349), .Y(n1040) );
  OAI21X1 U2319 ( .A(n2283), .B(n2311), .C(n1351), .Y(n1041) );
  OAI21X1 U2320 ( .A(n2283), .B(n2313), .C(n1353), .Y(n1042) );
  OAI21X1 U2321 ( .A(n2284), .B(n2315), .C(n1355), .Y(n1043) );
  OAI21X1 U2322 ( .A(n2284), .B(n2318), .C(n1357), .Y(n1044) );
  OAI21X1 U2323 ( .A(n2284), .B(n2320), .C(n1359), .Y(n1045) );
  OAI21X1 U2324 ( .A(n2284), .B(n2322), .C(n1515), .Y(n1046) );
  OAI21X1 U2325 ( .A(n2284), .B(n2325), .C(n1517), .Y(n1047) );
  OAI21X1 U2326 ( .A(n2284), .B(n2327), .C(n1519), .Y(n1048) );
  OAI21X1 U2327 ( .A(n2284), .B(n2328), .C(n1521), .Y(n1049) );
  OAI21X1 U2328 ( .A(n2284), .B(n2331), .C(n1523), .Y(n1050) );
  OAI21X1 U2329 ( .A(n2285), .B(n2300), .C(n1361), .Y(n1051) );
  OAI21X1 U2330 ( .A(n2285), .B(n2301), .C(n1363), .Y(n1052) );
  OAI21X1 U2331 ( .A(n2285), .B(n2303), .C(n1365), .Y(n1053) );
  OAI21X1 U2332 ( .A(n2285), .B(n2305), .C(n1367), .Y(n1054) );
  OAI21X1 U2333 ( .A(n2285), .B(n2307), .C(n1369), .Y(n1055) );
  OAI21X1 U2334 ( .A(n2285), .B(n2309), .C(n1371), .Y(n1056) );
  OAI21X1 U2335 ( .A(n2285), .B(n2311), .C(n1373), .Y(n1057) );
  OAI21X1 U2336 ( .A(n2285), .B(n2313), .C(n1375), .Y(n1058) );
  OAI21X1 U2337 ( .A(n2286), .B(n2315), .C(n1377), .Y(n1059) );
  OAI21X1 U2338 ( .A(n2286), .B(n2317), .C(n1379), .Y(n1060) );
  OAI21X1 U2339 ( .A(n2286), .B(n2319), .C(n1381), .Y(n1061) );
  OAI21X1 U2340 ( .A(n2286), .B(n2322), .C(n1525), .Y(n1062) );
  OAI21X1 U2341 ( .A(n2286), .B(n2324), .C(n1527), .Y(n1063) );
  OAI21X1 U2342 ( .A(n2286), .B(n2326), .C(n1529), .Y(n1064) );
  OAI21X1 U2343 ( .A(n2286), .B(n2328), .C(n1531), .Y(n1065) );
  OAI21X1 U2344 ( .A(n2286), .B(n2330), .C(n1533), .Y(n1066) );
  OAI21X1 U2345 ( .A(n2287), .B(n2300), .C(n1383), .Y(n1067) );
  OAI21X1 U2346 ( .A(n2287), .B(n2301), .C(n1385), .Y(n1068) );
  OAI21X1 U2347 ( .A(n2287), .B(n2303), .C(n1387), .Y(n1069) );
  OAI21X1 U2348 ( .A(n2287), .B(n2305), .C(n1389), .Y(n1070) );
  OAI21X1 U2349 ( .A(n2287), .B(n2307), .C(n1391), .Y(n1071) );
  OAI21X1 U2350 ( .A(n2287), .B(n2309), .C(n1393), .Y(n1072) );
  OAI21X1 U2351 ( .A(n2287), .B(n2311), .C(n1395), .Y(n1073) );
  OAI21X1 U2352 ( .A(n2287), .B(n2313), .C(n1397), .Y(n1074) );
  OAI21X1 U2353 ( .A(n2288), .B(n2315), .C(n1399), .Y(n1075) );
  OAI21X1 U2354 ( .A(n2288), .B(n2317), .C(n1401), .Y(n1076) );
  OAI21X1 U2355 ( .A(n2288), .B(n2319), .C(n1403), .Y(n1077) );
  OAI21X1 U2356 ( .A(n2288), .B(n2322), .C(n1535), .Y(n1078) );
  OAI21X1 U2357 ( .A(n2288), .B(n2324), .C(n1537), .Y(n1079) );
  OAI21X1 U2358 ( .A(n2288), .B(n2326), .C(n1539), .Y(n1080) );
  OAI21X1 U2359 ( .A(n2288), .B(n2328), .C(n1541), .Y(n1081) );
  OAI21X1 U2360 ( .A(n2288), .B(n2330), .C(n1543), .Y(n1082) );
  OAI21X1 U2361 ( .A(n2289), .B(n2300), .C(n1405), .Y(n1083) );
  OAI21X1 U2362 ( .A(n2289), .B(n2301), .C(n1407), .Y(n1084) );
  OAI21X1 U2363 ( .A(n2289), .B(n2303), .C(n1409), .Y(n1085) );
  OAI21X1 U2364 ( .A(n2289), .B(n2305), .C(n1411), .Y(n1086) );
  OAI21X1 U2365 ( .A(n2289), .B(n2307), .C(n1413), .Y(n1087) );
  OAI21X1 U2366 ( .A(n2289), .B(n2309), .C(n1415), .Y(n1088) );
  OAI21X1 U2367 ( .A(n2289), .B(n2311), .C(n1417), .Y(n1089) );
  OAI21X1 U2368 ( .A(n2289), .B(n2313), .C(n1419), .Y(n1090) );
  OAI21X1 U2369 ( .A(n2290), .B(n2315), .C(n1421), .Y(n1091) );
  OAI21X1 U2370 ( .A(n2290), .B(n2317), .C(n1423), .Y(n1092) );
  OAI21X1 U2371 ( .A(n2290), .B(n2319), .C(n1425), .Y(n1093) );
  OAI21X1 U2372 ( .A(n2290), .B(n6), .C(n1545), .Y(n1094) );
  OAI21X1 U2373 ( .A(n2290), .B(n2325), .C(n1547), .Y(n1095) );
  OAI21X1 U2374 ( .A(n2290), .B(n2327), .C(n1549), .Y(n1096) );
  OAI21X1 U2375 ( .A(n2290), .B(n2328), .C(n1551), .Y(n1097) );
  OAI21X1 U2376 ( .A(n2290), .B(n7), .C(n1553), .Y(n1098) );
  OAI21X1 U2377 ( .A(n2291), .B(n2300), .C(n1427), .Y(n1099) );
  OAI21X1 U2378 ( .A(n2291), .B(n2301), .C(n1429), .Y(n1100) );
  OAI21X1 U2379 ( .A(n2291), .B(n2303), .C(n1431), .Y(n1101) );
  OAI21X1 U2380 ( .A(n2291), .B(n2305), .C(n1433), .Y(n1102) );
  OAI21X1 U2381 ( .A(n2291), .B(n2307), .C(n1435), .Y(n1103) );
  OAI21X1 U2382 ( .A(n2291), .B(n2309), .C(n1437), .Y(n1104) );
  OAI21X1 U2383 ( .A(n2291), .B(n2311), .C(n1439), .Y(n1105) );
  OAI21X1 U2384 ( .A(n2291), .B(n2313), .C(n1441), .Y(n1106) );
  OAI21X1 U2385 ( .A(n2292), .B(n2315), .C(n1443), .Y(n1107) );
  OAI21X1 U2386 ( .A(n2292), .B(n2318), .C(n1445), .Y(n1108) );
  OAI21X1 U2387 ( .A(n2292), .B(n2319), .C(n1447), .Y(n1109) );
  OAI21X1 U2388 ( .A(n2292), .B(n2322), .C(n1555), .Y(n1110) );
  OAI21X1 U2389 ( .A(n2292), .B(n2324), .C(n1557), .Y(n1111) );
  OAI21X1 U2390 ( .A(n2292), .B(n2327), .C(n1559), .Y(n1112) );
  OAI21X1 U2391 ( .A(n2292), .B(n2328), .C(n1561), .Y(n1113) );
  OAI21X1 U2392 ( .A(n2292), .B(n7), .C(n1563), .Y(n1114) );
  OAI21X1 U2393 ( .A(n2293), .B(n2300), .C(n1449), .Y(n1115) );
  OAI21X1 U2394 ( .A(n2293), .B(n2301), .C(n1451), .Y(n1116) );
  OAI21X1 U2395 ( .A(n2293), .B(n2303), .C(n1453), .Y(n1117) );
  OAI21X1 U2396 ( .A(n2293), .B(n2305), .C(n1455), .Y(n1118) );
  OAI21X1 U2397 ( .A(n2293), .B(n2307), .C(n1457), .Y(n1119) );
  OAI21X1 U2398 ( .A(n2293), .B(n2309), .C(n1459), .Y(n1120) );
  OAI21X1 U2399 ( .A(n2293), .B(n2311), .C(n1461), .Y(n1121) );
  OAI21X1 U2400 ( .A(n2293), .B(n2313), .C(n1463), .Y(n1122) );
  OAI21X1 U2401 ( .A(n2294), .B(n2315), .C(n1465), .Y(n1123) );
  OAI21X1 U2402 ( .A(n2294), .B(n2318), .C(n1467), .Y(n1124) );
  OAI21X1 U2403 ( .A(n2294), .B(n2320), .C(n1469), .Y(n1125) );
  OAI21X1 U2404 ( .A(n2294), .B(n2321), .C(n1565), .Y(n1126) );
  OAI21X1 U2405 ( .A(n2294), .B(n2325), .C(n1567), .Y(n1127) );
  OAI21X1 U2406 ( .A(n2294), .B(n2327), .C(n1569), .Y(n1128) );
  OAI21X1 U2407 ( .A(n2294), .B(n2328), .C(n1571), .Y(n1129) );
  OAI21X1 U2408 ( .A(n2294), .B(n2331), .C(n1573), .Y(n1130) );
  OAI21X1 U2409 ( .A(n2295), .B(n2300), .C(n1471), .Y(n1131) );
  OAI21X1 U2410 ( .A(n2295), .B(n2301), .C(n1473), .Y(n1132) );
  OAI21X1 U2411 ( .A(n2295), .B(n2303), .C(n1475), .Y(n1133) );
  OAI21X1 U2412 ( .A(n2295), .B(n2305), .C(n1477), .Y(n1134) );
  OAI21X1 U2413 ( .A(n2295), .B(n2307), .C(n1479), .Y(n1135) );
  OAI21X1 U2414 ( .A(n2295), .B(n2309), .C(n1481), .Y(n1136) );
  OAI21X1 U2415 ( .A(n2295), .B(n2311), .C(n1483), .Y(n1137) );
  OAI21X1 U2416 ( .A(n2295), .B(n2313), .C(n1485), .Y(n1138) );
  OAI21X1 U2417 ( .A(n2296), .B(n2315), .C(n1487), .Y(n1139) );
  OAI21X1 U2418 ( .A(n2296), .B(n2318), .C(n1489), .Y(n1140) );
  OAI21X1 U2419 ( .A(n2296), .B(n2320), .C(n1491), .Y(n1141) );
  OAI21X1 U2420 ( .A(n2296), .B(n2322), .C(n1575), .Y(n1142) );
  OAI21X1 U2421 ( .A(n2296), .B(n2325), .C(n1577), .Y(n1143) );
  OAI21X1 U2422 ( .A(n2296), .B(n2327), .C(n1579), .Y(n1144) );
  OAI21X1 U2423 ( .A(n2296), .B(n2328), .C(n1581), .Y(n1145) );
  OAI21X1 U2424 ( .A(n2296), .B(n2331), .C(n1583), .Y(n1146) );
  OAI21X1 U2425 ( .A(n2297), .B(n2300), .C(n595), .Y(n1147) );
  OAI21X1 U2426 ( .A(n2297), .B(n2301), .C(n597), .Y(n1148) );
  OAI21X1 U2427 ( .A(n2297), .B(n2303), .C(n599), .Y(n1149) );
  OAI21X1 U2428 ( .A(n2297), .B(n2305), .C(n601), .Y(n1150) );
  OAI21X1 U2429 ( .A(n2297), .B(n2307), .C(n603), .Y(n1151) );
  OAI21X1 U2430 ( .A(n2297), .B(n2309), .C(n605), .Y(n1152) );
  OAI21X1 U2431 ( .A(n2297), .B(n2311), .C(n607), .Y(n1153) );
  OAI21X1 U2432 ( .A(n2297), .B(n2313), .C(n609), .Y(n1154) );
  OAI21X1 U2433 ( .A(n2297), .B(n2315), .C(n611), .Y(n1155) );
  OAI21X1 U2434 ( .A(n2297), .B(n2317), .C(n613), .Y(n1156) );
  OAI21X1 U2435 ( .A(n2297), .B(n2320), .C(n615), .Y(n1157) );
  OAI21X1 U2436 ( .A(n2297), .B(n6), .C(n1493), .Y(n1158) );
  OAI21X1 U2437 ( .A(n2297), .B(n2325), .C(n1495), .Y(n1159) );
  OAI21X1 U2438 ( .A(n2297), .B(n2326), .C(n1497), .Y(n1160) );
  OAI21X1 U2439 ( .A(n2297), .B(n2328), .C(n1499), .Y(n1161) );
  OAI21X1 U2440 ( .A(n2297), .B(n7), .C(n1501), .Y(n1162) );
endmodule


module memc_Size16_6 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n13,
         n14, n16, n18, n20, n22, n24, n26, n28, n30, n32, n34, n36, n38, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2462), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2463), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2464), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2465), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2466), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2467), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2468), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2469), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2470), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2471), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2472), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2473), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2474), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2475), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2476), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2477), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2478), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2479), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2480), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2481), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2482), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2483), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2484), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2485), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2486), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2487), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2488), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2489), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2490), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2491), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2492), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2493), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2494), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2495), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2496), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2497), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2498), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2499), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2500), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2501), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2502), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2503), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2504), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2505), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2506), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2507), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2508), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2509), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2510), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2511), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2512), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2513), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2514), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2515), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2516), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2517), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2518), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2519), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2520), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2521), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2522), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2523), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2524), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2525), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2526), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2527), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2528), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2529), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2530), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2531), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2532), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2533), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2534), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2535), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2536), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2537), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2538), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2539), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2540), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2541), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2542), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2543), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2544), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2545), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2546), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2547), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2548), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2549), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2550), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2551), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2552), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2553), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2554), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2555), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2556), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2557), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2558), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2559), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2560), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2561), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2562), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2563), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2564), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2565), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2566), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2567), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2568), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2569), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2570), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2571), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2572), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2573), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2574), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2575), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2576), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2577), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2578), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2579), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2580), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2581), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2582), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2583), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2584), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2585), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2586), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2587), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2588), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2589), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2590), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2591), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2592), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2593), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2594), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2595), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2596), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2597), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2598), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2599), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2600), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2601), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2602), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2603), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2604), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2605), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2606), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2607), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2608), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2609), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2610), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2611), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2612), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2613), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2614), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2615), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2616), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2617), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2618), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2619), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2620), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2621), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2622), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2623), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2624), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2625), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2626), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2627), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2628), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2629), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2630), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2631), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2632), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2633), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2634), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2635), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2636), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2637), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2638), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2639), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2640), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2641), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2642), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2643), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2644), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2645), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2646), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2647), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2648), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2649), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2650), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2651), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2652), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2653), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2654), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2655), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2656), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2657), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2658), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2659), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2660), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2661), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2662), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2663), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2664), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2665), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2666), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2667), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2668), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2669), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2670), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2671), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2672), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2673), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2674), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2675), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2676), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2677), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2678), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2679), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2680), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2681), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2682), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2683), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2684), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2685), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2686), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2687), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2688), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2689), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2690), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2691), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2692), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2693), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2694), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2695), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2696), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2697), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2698), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2699), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2700), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2701), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2702), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2703), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2704), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2705), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2706), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2707), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2708), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2709), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2710), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2711), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2712), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2713), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2714), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2715), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2716), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2717), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2718), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2719), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2720), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2721), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2722), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2723), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2724), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2725), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2726), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2727), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2728), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2729), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2730), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2731), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2732), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2733), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2734), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2735), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2736), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2737), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2738), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2739), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2740), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2741), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2742), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2743), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2744), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2745), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2746), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2747), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2748), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2749), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2750), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2751), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2752), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2753), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2754), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2755), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2756), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2757), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2758), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2759), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2760), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2761), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2762), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2763), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2764), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2765), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2766), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2767), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2768), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2769), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2770), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2771), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2772), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2773), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2774), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2775), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2776), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2777), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2778), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2779), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2780), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2781), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2782), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2783), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2784), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2785), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2786), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2787), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2788), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2789), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2790), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2791), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2792), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2793), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2794), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2795), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2796), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2797), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2798), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2799), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2800), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2801), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2802), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2803), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2804), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2805), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2806), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2807), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2808), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2809), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2810), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2811), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2812), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2813), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2814), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2815), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2816), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2817), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2818), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2819), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2820), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2821), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2822), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2823), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2824), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2825), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2826), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2827), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2828), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2829), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2830), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2831), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2832), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2833), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2834), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2835), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2836), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2837), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2838), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2839), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2840), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2841), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2842), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2843), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2844), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2845), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2846), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2847), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2848), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2849), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2850), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2851), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2852), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2853), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2854), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2855), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2856), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2857), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2858), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2859), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2860), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2861), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2862), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2863), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2864), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2865), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2866), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2867), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2868), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2869), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2870), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2871), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2872), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2873), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2874), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2875), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2876), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2877), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2878), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2879), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2880), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2881), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2882), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2883), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2884), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2885), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2886), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2887), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2888), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2889), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2890), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2891), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2892), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2893), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2894), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2895), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2896), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2897), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2898), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2899), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2900), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2901), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2902), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2903), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2904), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2905), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2906), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2907), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2908), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2909), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2910), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2911), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2912), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2913), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2914), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2915), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2916), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2917), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2918), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2919), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2920), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2921), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2922), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2923), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2924), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2925), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2926), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2927), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2928), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2929), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2930), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2931), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2932), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2933), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2934), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2935), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2936), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2937), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2938), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2939), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2940), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2941), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2942), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2943), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2944), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2945), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2946), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2947), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2948), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2949), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2950), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2951), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2952), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2953), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2954), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2955), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2956), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2957), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2958), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2959), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2960), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2961), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2962), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2963), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2964), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2965), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2966), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2967), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2968), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2969), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2970), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2971), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2972), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2973), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2974) );
  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n1418), .Y(n2) );
  INVX4 U4 ( .A(n42), .Y(n43) );
  INVX4 U5 ( .A(n40), .Y(n41) );
  INVX1 U6 ( .A(n2426), .Y(n2280) );
  INVX1 U7 ( .A(n2428), .Y(n2277) );
  INVX1 U8 ( .A(n2428), .Y(n2276) );
  INVX2 U9 ( .A(n2284), .Y(n2288) );
  INVX2 U10 ( .A(n2284), .Y(n2289) );
  INVX1 U11 ( .A(n2425), .Y(n2278) );
  INVX2 U12 ( .A(n2284), .Y(n2290) );
  INVX2 U13 ( .A(n2284), .Y(n2293) );
  INVX2 U14 ( .A(n2284), .Y(n2295) );
  INVX1 U15 ( .A(n2284), .Y(n2285) );
  INVX2 U16 ( .A(n2284), .Y(n2287) );
  INVX2 U17 ( .A(n2284), .Y(n2286) );
  INVX2 U18 ( .A(n2278), .Y(n2283) );
  INVX2 U19 ( .A(n2278), .Y(n2282) );
  INVX2 U20 ( .A(n2278), .Y(n2281) );
  INVX2 U21 ( .A(n2284), .Y(n2291) );
  INVX2 U22 ( .A(n2284), .Y(n2294) );
  INVX1 U23 ( .A(n2259), .Y(N32) );
  INVX1 U24 ( .A(n2260), .Y(N31) );
  INVX1 U25 ( .A(n2261), .Y(N30) );
  INVX1 U26 ( .A(n2262), .Y(N29) );
  INVX1 U27 ( .A(n2263), .Y(N28) );
  INVX1 U28 ( .A(n2264), .Y(N27) );
  INVX1 U29 ( .A(n2265), .Y(N26) );
  INVX1 U30 ( .A(n2266), .Y(N25) );
  INVX1 U31 ( .A(n2267), .Y(N24) );
  INVX1 U32 ( .A(n2268), .Y(N23) );
  INVX1 U33 ( .A(n2269), .Y(N22) );
  INVX1 U34 ( .A(n2270), .Y(N21) );
  INVX1 U35 ( .A(n2271), .Y(N20) );
  INVX1 U36 ( .A(n2272), .Y(N19) );
  INVX1 U37 ( .A(n2273), .Y(N18) );
  INVX1 U38 ( .A(n2274), .Y(N17) );
  BUFX2 U39 ( .A(n1724), .Y(n2329) );
  BUFX2 U40 ( .A(n1726), .Y(n2331) );
  BUFX2 U41 ( .A(n1728), .Y(n2333) );
  BUFX2 U42 ( .A(n1730), .Y(n2335) );
  BUFX2 U43 ( .A(n1732), .Y(n2337) );
  BUFX2 U44 ( .A(n1734), .Y(n2339) );
  BUFX2 U45 ( .A(n1736), .Y(n2341) );
  BUFX2 U46 ( .A(n1738), .Y(n2344) );
  BUFX2 U47 ( .A(n1740), .Y(n2346) );
  BUFX2 U48 ( .A(n1742), .Y(n2348) );
  BUFX2 U49 ( .A(n1744), .Y(n2350) );
  BUFX2 U50 ( .A(n1746), .Y(n2352) );
  BUFX2 U51 ( .A(n1748), .Y(n2354) );
  BUFX2 U52 ( .A(n1750), .Y(n2356) );
  BUFX2 U53 ( .A(n1752), .Y(n2359) );
  BUFX2 U54 ( .A(n1754), .Y(n2361) );
  BUFX2 U55 ( .A(n1756), .Y(n2363) );
  BUFX2 U56 ( .A(n1758), .Y(n2365) );
  BUFX2 U57 ( .A(n1760), .Y(n2367) );
  BUFX2 U58 ( .A(n1762), .Y(n2369) );
  BUFX2 U59 ( .A(n1764), .Y(n2371) );
  BUFX2 U60 ( .A(n1766), .Y(n2374) );
  BUFX2 U61 ( .A(n1768), .Y(n2376) );
  BUFX2 U62 ( .A(n1770), .Y(n2378) );
  BUFX2 U63 ( .A(n1772), .Y(n2380) );
  BUFX2 U64 ( .A(n1774), .Y(n2382) );
  BUFX2 U65 ( .A(n1776), .Y(n2384) );
  BUFX2 U66 ( .A(n1778), .Y(n2386) );
  INVX1 U67 ( .A(n2424), .Y(n2296) );
  INVX2 U68 ( .A(n2284), .Y(n2292) );
  INVX4 U69 ( .A(n2422), .Y(n2326) );
  INVX2 U70 ( .A(n2327), .Y(n2297) );
  INVX1 U71 ( .A(n2430), .Y(n2429) );
  INVX1 U72 ( .A(N14), .Y(n2430) );
  INVX1 U73 ( .A(N12), .Y(n2426) );
  INVX2 U74 ( .A(n2426), .Y(n2279) );
  INVX1 U75 ( .A(n2428), .Y(n2427) );
  INVX1 U76 ( .A(N13), .Y(n2428) );
  INVX1 U77 ( .A(n1721), .Y(n2373) );
  INVX1 U78 ( .A(n1722), .Y(n2388) );
  BUFX2 U79 ( .A(n1774), .Y(n2383) );
  BUFX2 U80 ( .A(n1778), .Y(n2387) );
  INVX1 U81 ( .A(n2430), .Y(n2275) );
  INVX1 U82 ( .A(rst), .Y(n2421) );
  INVX1 U83 ( .A(n1720), .Y(n2358) );
  BUFX2 U84 ( .A(n1724), .Y(n2330) );
  BUFX2 U85 ( .A(n1748), .Y(n2355) );
  BUFX2 U86 ( .A(n1752), .Y(n2360) );
  BUFX2 U87 ( .A(n1754), .Y(n2362) );
  BUFX2 U88 ( .A(n1758), .Y(n2366) );
  BUFX2 U89 ( .A(n1760), .Y(n2368) );
  BUFX2 U90 ( .A(n1762), .Y(n2370) );
  BUFX2 U91 ( .A(n1764), .Y(n2372) );
  BUFX2 U92 ( .A(n1766), .Y(n2375) );
  BUFX2 U93 ( .A(n1768), .Y(n2377) );
  BUFX2 U94 ( .A(n1770), .Y(n2379) );
  BUFX2 U95 ( .A(n1772), .Y(n2381) );
  BUFX2 U96 ( .A(n1776), .Y(n2385) );
  BUFX2 U97 ( .A(n1756), .Y(n2364) );
  BUFX2 U98 ( .A(n1750), .Y(n2357) );
  BUFX2 U99 ( .A(n1746), .Y(n2353) );
  BUFX2 U100 ( .A(n1744), .Y(n2351) );
  BUFX2 U101 ( .A(n1742), .Y(n2349) );
  BUFX2 U102 ( .A(n1740), .Y(n2347) );
  BUFX2 U103 ( .A(n1738), .Y(n2345) );
  BUFX2 U104 ( .A(n1736), .Y(n2342) );
  BUFX2 U105 ( .A(n1734), .Y(n2340) );
  BUFX2 U106 ( .A(n1732), .Y(n2338) );
  BUFX2 U107 ( .A(n1730), .Y(n2336) );
  BUFX2 U108 ( .A(n1728), .Y(n2334) );
  BUFX2 U109 ( .A(n1726), .Y(n2332) );
  INVX1 U110 ( .A(n1719), .Y(n2343) );
  INVX1 U111 ( .A(n1418), .Y(n3) );
  INVX1 U112 ( .A(n1418), .Y(n4) );
  INVX1 U113 ( .A(write), .Y(n5) );
  INVX1 U114 ( .A(write), .Y(n6) );
  INVX1 U115 ( .A(write), .Y(n1418) );
  INVX1 U116 ( .A(n6), .Y(n7) );
  INVX1 U117 ( .A(n5), .Y(n8) );
  INVX1 U118 ( .A(n5), .Y(n9) );
  INVX1 U119 ( .A(n136), .Y(n10) );
  AND2X2 U120 ( .A(n1679), .B(n10), .Y(\data_out<1> ) );
  AND2X2 U121 ( .A(n5), .B(n1696), .Y(\data_out<10> ) );
  OR2X2 U122 ( .A(n8), .B(n1678), .Y(n13) );
  OR2X2 U123 ( .A(n3), .B(n1681), .Y(n14) );
  INVX1 U124 ( .A(n14), .Y(\data_out<2> ) );
  OR2X2 U125 ( .A(n4), .B(n1683), .Y(n16) );
  INVX1 U126 ( .A(n16), .Y(\data_out<3> ) );
  OR2X2 U127 ( .A(n9), .B(n1685), .Y(n18) );
  INVX1 U128 ( .A(n18), .Y(\data_out<4> ) );
  OR2X2 U129 ( .A(n4), .B(n1687), .Y(n20) );
  INVX1 U130 ( .A(n20), .Y(\data_out<5> ) );
  OR2X2 U131 ( .A(n9), .B(n1689), .Y(n22) );
  INVX1 U132 ( .A(n22), .Y(\data_out<6> ) );
  OR2X2 U133 ( .A(n7), .B(n1691), .Y(n24) );
  INVX1 U134 ( .A(n24), .Y(\data_out<7> ) );
  OR2X2 U135 ( .A(n7), .B(n1693), .Y(n26) );
  INVX1 U136 ( .A(n26), .Y(\data_out<8> ) );
  OR2X2 U137 ( .A(n136), .B(n1695), .Y(n28) );
  INVX1 U138 ( .A(n28), .Y(\data_out<9> ) );
  OR2X2 U139 ( .A(n2), .B(n1698), .Y(n30) );
  INVX1 U140 ( .A(n30), .Y(\data_out<11> ) );
  OR2X2 U141 ( .A(n2), .B(n1700), .Y(n32) );
  INVX1 U142 ( .A(n32), .Y(\data_out<12> ) );
  OR2X2 U143 ( .A(n7), .B(n1702), .Y(n34) );
  INVX1 U144 ( .A(n34), .Y(\data_out<13> ) );
  OR2X2 U145 ( .A(n3), .B(n1704), .Y(n36) );
  INVX1 U146 ( .A(n36), .Y(\data_out<14> ) );
  OR2X2 U147 ( .A(n8), .B(n1706), .Y(n38) );
  INVX1 U148 ( .A(n38), .Y(\data_out<15> ) );
  AND2X2 U149 ( .A(n2461), .B(n1719), .Y(n40) );
  AND2X2 U150 ( .A(n2461), .B(n1747), .Y(n42) );
  AND2X2 U151 ( .A(n2461), .B(n1720), .Y(n44) );
  INVX1 U152 ( .A(n44), .Y(n45) );
  INVX1 U153 ( .A(n44), .Y(n46) );
  AND2X2 U154 ( .A(n2461), .B(n1751), .Y(n47) );
  INVX1 U155 ( .A(n47), .Y(n48) );
  INVX1 U156 ( .A(n47), .Y(n49) );
  AND2X2 U157 ( .A(n2461), .B(n1753), .Y(n50) );
  INVX1 U158 ( .A(n50), .Y(n51) );
  INVX1 U159 ( .A(n50), .Y(n52) );
  AND2X2 U160 ( .A(n2461), .B(n1757), .Y(n53) );
  INVX1 U161 ( .A(n53), .Y(n54) );
  INVX1 U162 ( .A(n53), .Y(n55) );
  AND2X2 U163 ( .A(n2461), .B(n1759), .Y(n56) );
  INVX1 U164 ( .A(n56), .Y(n57) );
  INVX1 U165 ( .A(n56), .Y(n58) );
  AND2X2 U166 ( .A(n2461), .B(n1761), .Y(n59) );
  INVX1 U167 ( .A(n59), .Y(n60) );
  INVX1 U168 ( .A(n59), .Y(n61) );
  AND2X2 U169 ( .A(n2461), .B(n1763), .Y(n62) );
  INVX1 U170 ( .A(n62), .Y(n63) );
  INVX1 U171 ( .A(n62), .Y(n64) );
  AND2X2 U172 ( .A(n2461), .B(n1721), .Y(n65) );
  INVX1 U173 ( .A(n65), .Y(n66) );
  INVX1 U174 ( .A(n65), .Y(n67) );
  AND2X2 U175 ( .A(n2461), .B(n1765), .Y(n68) );
  INVX1 U176 ( .A(n68), .Y(n69) );
  INVX1 U177 ( .A(n68), .Y(n70) );
  AND2X2 U178 ( .A(n2461), .B(n1767), .Y(n71) );
  INVX1 U179 ( .A(n71), .Y(n72) );
  INVX1 U180 ( .A(n71), .Y(n73) );
  AND2X2 U181 ( .A(n2461), .B(n1769), .Y(n74) );
  INVX1 U182 ( .A(n74), .Y(n75) );
  INVX1 U183 ( .A(n74), .Y(n76) );
  AND2X2 U184 ( .A(n2461), .B(n1771), .Y(n77) );
  INVX1 U185 ( .A(n77), .Y(n78) );
  INVX1 U186 ( .A(n77), .Y(n79) );
  AND2X2 U187 ( .A(n2461), .B(n1773), .Y(n80) );
  INVX1 U188 ( .A(n80), .Y(n81) );
  INVX1 U189 ( .A(n80), .Y(n82) );
  AND2X2 U190 ( .A(n2461), .B(n1775), .Y(n83) );
  INVX1 U191 ( .A(n83), .Y(n84) );
  INVX1 U192 ( .A(n83), .Y(n85) );
  AND2X2 U193 ( .A(n2461), .B(n1777), .Y(n86) );
  INVX1 U194 ( .A(n86), .Y(n87) );
  INVX1 U195 ( .A(n86), .Y(n88) );
  AND2X2 U196 ( .A(n2461), .B(n1722), .Y(n89) );
  INVX1 U197 ( .A(n89), .Y(n90) );
  INVX1 U198 ( .A(n89), .Y(n91) );
  AND2X2 U199 ( .A(\data_in<0> ), .B(n2461), .Y(n92) );
  AND2X2 U200 ( .A(\data_in<1> ), .B(n2461), .Y(n93) );
  AND2X2 U201 ( .A(\data_in<2> ), .B(n2461), .Y(n94) );
  AND2X2 U202 ( .A(\data_in<3> ), .B(n2461), .Y(n95) );
  AND2X2 U203 ( .A(\data_in<4> ), .B(n2461), .Y(n96) );
  AND2X2 U204 ( .A(\data_in<5> ), .B(n2461), .Y(n97) );
  AND2X2 U205 ( .A(\data_in<6> ), .B(n2461), .Y(n98) );
  AND2X2 U206 ( .A(\data_in<7> ), .B(n2461), .Y(n99) );
  AND2X2 U207 ( .A(\data_in<8> ), .B(n2461), .Y(n100) );
  AND2X2 U208 ( .A(\data_in<9> ), .B(n2461), .Y(n101) );
  AND2X2 U209 ( .A(\data_in<10> ), .B(n2461), .Y(n102) );
  AND2X2 U210 ( .A(\data_in<11> ), .B(n2461), .Y(n103) );
  AND2X2 U211 ( .A(\data_in<12> ), .B(n2461), .Y(n104) );
  AND2X2 U212 ( .A(\data_in<13> ), .B(n2461), .Y(n105) );
  AND2X2 U213 ( .A(\data_in<14> ), .B(n2461), .Y(n106) );
  AND2X2 U214 ( .A(\data_in<15> ), .B(n2461), .Y(n107) );
  INVX1 U215 ( .A(n122), .Y(n108) );
  INVX1 U216 ( .A(n123), .Y(n109) );
  INVX1 U217 ( .A(n124), .Y(n110) );
  INVX1 U218 ( .A(n125), .Y(n111) );
  INVX1 U219 ( .A(n126), .Y(n112) );
  INVX1 U220 ( .A(n127), .Y(n113) );
  INVX1 U221 ( .A(n128), .Y(n114) );
  INVX1 U222 ( .A(n129), .Y(n115) );
  INVX1 U223 ( .A(n130), .Y(n116) );
  INVX1 U224 ( .A(n131), .Y(n117) );
  INVX1 U225 ( .A(n132), .Y(n118) );
  INVX1 U226 ( .A(n133), .Y(n119) );
  INVX1 U227 ( .A(n134), .Y(n120) );
  INVX2 U228 ( .A(n135), .Y(n121) );
  INVX2 U229 ( .A(n135), .Y(n2432) );
  AND2X2 U230 ( .A(n2461), .B(n1755), .Y(n122) );
  INVX4 U231 ( .A(n122), .Y(n2451) );
  AND2X2 U232 ( .A(n2461), .B(n1749), .Y(n123) );
  INVX4 U233 ( .A(n123), .Y(n2449) );
  AND2X2 U234 ( .A(n2461), .B(n1745), .Y(n124) );
  INVX4 U235 ( .A(n124), .Y(n2448) );
  AND2X2 U236 ( .A(n2461), .B(n1743), .Y(n125) );
  INVX4 U237 ( .A(n125), .Y(n2447) );
  AND2X2 U238 ( .A(n2461), .B(n1741), .Y(n126) );
  INVX4 U239 ( .A(n126), .Y(n2446) );
  AND2X2 U240 ( .A(n2461), .B(n1739), .Y(n127) );
  INVX4 U241 ( .A(n127), .Y(n2445) );
  AND2X2 U242 ( .A(n2461), .B(n1737), .Y(n128) );
  INVX4 U243 ( .A(n128), .Y(n2444) );
  AND2X2 U244 ( .A(n2461), .B(n1735), .Y(n129) );
  INVX4 U245 ( .A(n129), .Y(n2443) );
  AND2X2 U246 ( .A(n2461), .B(n1733), .Y(n130) );
  INVX4 U247 ( .A(n130), .Y(n2441) );
  AND2X2 U248 ( .A(n2461), .B(n1731), .Y(n131) );
  INVX4 U249 ( .A(n131), .Y(n2439) );
  AND2X2 U250 ( .A(n2461), .B(n1729), .Y(n132) );
  INVX4 U251 ( .A(n132), .Y(n2437) );
  AND2X2 U252 ( .A(n2461), .B(n1727), .Y(n133) );
  INVX4 U253 ( .A(n133), .Y(n2435) );
  AND2X2 U254 ( .A(n2461), .B(n1725), .Y(n134) );
  INVX4 U255 ( .A(n134), .Y(n2433) );
  AND2X2 U256 ( .A(n2461), .B(n1723), .Y(n135) );
  INVX1 U257 ( .A(n6), .Y(n136) );
  OR2X2 U258 ( .A(n1), .B(rst), .Y(n2431) );
  AND2X2 U259 ( .A(\mem<31><0> ), .B(n2432), .Y(n137) );
  INVX1 U260 ( .A(n137), .Y(n138) );
  AND2X2 U261 ( .A(\mem<30><0> ), .B(n2433), .Y(n139) );
  INVX1 U262 ( .A(n139), .Y(n140) );
  AND2X2 U263 ( .A(\mem<29><0> ), .B(n2435), .Y(n141) );
  INVX1 U264 ( .A(n141), .Y(n142) );
  AND2X2 U265 ( .A(\mem<28><0> ), .B(n2437), .Y(n143) );
  INVX1 U266 ( .A(n143), .Y(n144) );
  AND2X2 U267 ( .A(\mem<27><0> ), .B(n2439), .Y(n145) );
  INVX1 U268 ( .A(n145), .Y(n146) );
  AND2X2 U269 ( .A(n116), .B(\mem<26><0> ), .Y(n147) );
  INVX1 U270 ( .A(n147), .Y(n148) );
  AND2X2 U271 ( .A(n115), .B(\mem<25><0> ), .Y(n149) );
  INVX1 U272 ( .A(n149), .Y(n150) );
  AND2X2 U273 ( .A(n41), .B(\mem<24><0> ), .Y(n151) );
  INVX1 U274 ( .A(n151), .Y(n152) );
  AND2X2 U275 ( .A(n114), .B(\mem<23><0> ), .Y(n153) );
  INVX1 U276 ( .A(n153), .Y(n154) );
  AND2X2 U277 ( .A(n114), .B(\mem<23><1> ), .Y(n155) );
  INVX1 U278 ( .A(n155), .Y(n156) );
  AND2X2 U279 ( .A(\mem<23><2> ), .B(n2444), .Y(n157) );
  INVX1 U280 ( .A(n157), .Y(n158) );
  AND2X2 U281 ( .A(\mem<23><3> ), .B(n2444), .Y(n159) );
  INVX1 U282 ( .A(n159), .Y(n160) );
  AND2X2 U283 ( .A(\mem<23><4> ), .B(n2444), .Y(n161) );
  INVX1 U284 ( .A(n161), .Y(n162) );
  AND2X2 U285 ( .A(n114), .B(\mem<23><5> ), .Y(n163) );
  INVX1 U286 ( .A(n163), .Y(n164) );
  AND2X2 U287 ( .A(\mem<23><6> ), .B(n2444), .Y(n165) );
  INVX1 U288 ( .A(n165), .Y(n166) );
  AND2X2 U289 ( .A(\mem<23><7> ), .B(n2444), .Y(n167) );
  INVX1 U290 ( .A(n167), .Y(n168) );
  AND2X2 U291 ( .A(n2444), .B(\mem<23><8> ), .Y(n169) );
  INVX1 U292 ( .A(n169), .Y(n170) );
  AND2X2 U293 ( .A(n114), .B(\mem<23><9> ), .Y(n171) );
  INVX1 U294 ( .A(n171), .Y(n172) );
  AND2X2 U295 ( .A(\mem<23><10> ), .B(n2444), .Y(n173) );
  INVX1 U296 ( .A(n173), .Y(n174) );
  AND2X2 U297 ( .A(\mem<23><11> ), .B(n2444), .Y(n175) );
  INVX1 U298 ( .A(n175), .Y(n176) );
  AND2X2 U299 ( .A(\mem<23><12> ), .B(n2444), .Y(n177) );
  INVX1 U300 ( .A(n177), .Y(n178) );
  AND2X2 U301 ( .A(n2444), .B(\mem<23><13> ), .Y(n179) );
  INVX1 U302 ( .A(n179), .Y(n180) );
  AND2X2 U303 ( .A(\mem<23><14> ), .B(n2444), .Y(n181) );
  INVX1 U304 ( .A(n181), .Y(n182) );
  AND2X2 U305 ( .A(\mem<23><15> ), .B(n2444), .Y(n183) );
  INVX1 U306 ( .A(n183), .Y(n184) );
  AND2X2 U307 ( .A(n113), .B(\mem<22><0> ), .Y(n185) );
  INVX1 U308 ( .A(n185), .Y(n186) );
  AND2X2 U309 ( .A(n113), .B(\mem<22><1> ), .Y(n187) );
  INVX1 U310 ( .A(n187), .Y(n188) );
  AND2X2 U311 ( .A(\mem<22><2> ), .B(n2445), .Y(n189) );
  INVX1 U312 ( .A(n189), .Y(n190) );
  AND2X2 U313 ( .A(\mem<22><3> ), .B(n2445), .Y(n191) );
  INVX1 U314 ( .A(n191), .Y(n192) );
  AND2X2 U315 ( .A(\mem<22><4> ), .B(n2445), .Y(n193) );
  INVX1 U316 ( .A(n193), .Y(n194) );
  AND2X2 U317 ( .A(n113), .B(\mem<22><5> ), .Y(n195) );
  INVX1 U318 ( .A(n195), .Y(n196) );
  AND2X2 U319 ( .A(\mem<22><6> ), .B(n2445), .Y(n197) );
  INVX1 U320 ( .A(n197), .Y(n198) );
  AND2X2 U321 ( .A(\mem<22><7> ), .B(n2445), .Y(n199) );
  INVX1 U322 ( .A(n199), .Y(n200) );
  AND2X2 U323 ( .A(n2445), .B(\mem<22><8> ), .Y(n201) );
  INVX1 U324 ( .A(n201), .Y(n202) );
  AND2X2 U325 ( .A(n113), .B(\mem<22><9> ), .Y(n203) );
  INVX1 U326 ( .A(n203), .Y(n204) );
  AND2X2 U327 ( .A(\mem<22><10> ), .B(n2445), .Y(n205) );
  INVX1 U328 ( .A(n205), .Y(n206) );
  AND2X2 U329 ( .A(\mem<22><11> ), .B(n2445), .Y(n207) );
  INVX1 U330 ( .A(n207), .Y(n208) );
  AND2X2 U331 ( .A(\mem<22><12> ), .B(n2445), .Y(n209) );
  INVX1 U332 ( .A(n209), .Y(n210) );
  AND2X2 U333 ( .A(n2445), .B(\mem<22><13> ), .Y(n211) );
  INVX1 U334 ( .A(n211), .Y(n212) );
  AND2X2 U335 ( .A(\mem<22><14> ), .B(n2445), .Y(n213) );
  INVX1 U336 ( .A(n213), .Y(n215) );
  AND2X2 U337 ( .A(\mem<22><15> ), .B(n2445), .Y(n216) );
  INVX1 U338 ( .A(n216), .Y(n217) );
  AND2X2 U339 ( .A(n112), .B(\mem<21><0> ), .Y(n218) );
  INVX1 U340 ( .A(n218), .Y(n219) );
  AND2X2 U341 ( .A(n112), .B(\mem<21><1> ), .Y(n220) );
  INVX1 U342 ( .A(n220), .Y(n221) );
  AND2X2 U343 ( .A(\mem<21><2> ), .B(n2446), .Y(n222) );
  INVX1 U344 ( .A(n222), .Y(n223) );
  AND2X2 U345 ( .A(\mem<21><3> ), .B(n2446), .Y(n224) );
  INVX1 U346 ( .A(n224), .Y(n225) );
  AND2X2 U347 ( .A(\mem<21><4> ), .B(n2446), .Y(n226) );
  INVX1 U348 ( .A(n226), .Y(n227) );
  AND2X2 U349 ( .A(n112), .B(\mem<21><5> ), .Y(n228) );
  INVX1 U350 ( .A(n228), .Y(n229) );
  AND2X2 U351 ( .A(\mem<21><6> ), .B(n2446), .Y(n230) );
  INVX1 U352 ( .A(n230), .Y(n231) );
  AND2X2 U353 ( .A(\mem<21><7> ), .B(n2446), .Y(n232) );
  INVX1 U354 ( .A(n232), .Y(n233) );
  AND2X2 U355 ( .A(n2446), .B(\mem<21><8> ), .Y(n234) );
  INVX1 U356 ( .A(n234), .Y(n235) );
  AND2X2 U357 ( .A(n112), .B(\mem<21><9> ), .Y(n236) );
  INVX1 U358 ( .A(n236), .Y(n237) );
  AND2X2 U359 ( .A(\mem<21><10> ), .B(n2446), .Y(n238) );
  INVX1 U360 ( .A(n238), .Y(n239) );
  AND2X2 U361 ( .A(\mem<21><11> ), .B(n2446), .Y(n240) );
  INVX1 U362 ( .A(n240), .Y(n241) );
  AND2X2 U363 ( .A(\mem<21><12> ), .B(n2446), .Y(n242) );
  INVX1 U364 ( .A(n242), .Y(n243) );
  AND2X2 U365 ( .A(n2446), .B(\mem<21><13> ), .Y(n244) );
  INVX1 U366 ( .A(n244), .Y(n245) );
  AND2X2 U367 ( .A(\mem<21><14> ), .B(n2446), .Y(n246) );
  INVX1 U368 ( .A(n246), .Y(n247) );
  AND2X2 U369 ( .A(\mem<21><15> ), .B(n2446), .Y(n248) );
  INVX1 U370 ( .A(n248), .Y(n249) );
  AND2X2 U371 ( .A(n111), .B(\mem<20><0> ), .Y(n250) );
  INVX1 U372 ( .A(n250), .Y(n251) );
  AND2X2 U373 ( .A(n111), .B(\mem<20><1> ), .Y(n252) );
  INVX1 U374 ( .A(n252), .Y(n253) );
  AND2X2 U375 ( .A(\mem<20><2> ), .B(n2447), .Y(n254) );
  INVX1 U376 ( .A(n254), .Y(n255) );
  AND2X2 U377 ( .A(\mem<20><3> ), .B(n2447), .Y(n256) );
  INVX1 U378 ( .A(n256), .Y(n257) );
  AND2X2 U379 ( .A(\mem<20><4> ), .B(n2447), .Y(n258) );
  INVX1 U380 ( .A(n258), .Y(n259) );
  AND2X2 U381 ( .A(n111), .B(\mem<20><5> ), .Y(n260) );
  INVX1 U382 ( .A(n260), .Y(n261) );
  AND2X2 U383 ( .A(\mem<20><6> ), .B(n2447), .Y(n262) );
  INVX1 U384 ( .A(n262), .Y(n263) );
  AND2X2 U385 ( .A(\mem<20><7> ), .B(n2447), .Y(n264) );
  INVX1 U386 ( .A(n264), .Y(n265) );
  AND2X2 U387 ( .A(n2447), .B(\mem<20><8> ), .Y(n266) );
  INVX1 U388 ( .A(n266), .Y(n267) );
  AND2X2 U389 ( .A(n111), .B(\mem<20><9> ), .Y(n268) );
  INVX1 U390 ( .A(n268), .Y(n269) );
  AND2X2 U391 ( .A(\mem<20><10> ), .B(n2447), .Y(n270) );
  INVX1 U392 ( .A(n270), .Y(n271) );
  AND2X2 U393 ( .A(\mem<20><11> ), .B(n2447), .Y(n272) );
  INVX1 U394 ( .A(n272), .Y(n273) );
  AND2X2 U395 ( .A(\mem<20><12> ), .B(n2447), .Y(n274) );
  INVX1 U396 ( .A(n274), .Y(n275) );
  AND2X2 U397 ( .A(n2447), .B(\mem<20><13> ), .Y(n276) );
  INVX1 U398 ( .A(n276), .Y(n277) );
  AND2X2 U399 ( .A(\mem<20><14> ), .B(n2447), .Y(n278) );
  INVX1 U400 ( .A(n278), .Y(n279) );
  AND2X2 U401 ( .A(\mem<20><15> ), .B(n2447), .Y(n280) );
  INVX1 U402 ( .A(n280), .Y(n281) );
  AND2X2 U403 ( .A(n110), .B(\mem<19><0> ), .Y(n282) );
  INVX1 U404 ( .A(n282), .Y(n283) );
  AND2X2 U405 ( .A(n110), .B(\mem<19><1> ), .Y(n284) );
  INVX1 U406 ( .A(n284), .Y(n285) );
  AND2X2 U407 ( .A(\mem<19><2> ), .B(n2448), .Y(n286) );
  INVX1 U408 ( .A(n286), .Y(n287) );
  AND2X2 U409 ( .A(\mem<19><3> ), .B(n2448), .Y(n288) );
  INVX1 U410 ( .A(n288), .Y(n289) );
  AND2X2 U411 ( .A(\mem<19><4> ), .B(n2448), .Y(n290) );
  INVX1 U412 ( .A(n290), .Y(n291) );
  AND2X2 U413 ( .A(n110), .B(\mem<19><5> ), .Y(n292) );
  INVX1 U414 ( .A(n292), .Y(n293) );
  AND2X2 U415 ( .A(\mem<19><6> ), .B(n2448), .Y(n294) );
  INVX1 U416 ( .A(n294), .Y(n295) );
  AND2X2 U417 ( .A(\mem<19><7> ), .B(n2448), .Y(n296) );
  INVX1 U418 ( .A(n296), .Y(n297) );
  AND2X2 U419 ( .A(n2448), .B(\mem<19><8> ), .Y(n298) );
  INVX1 U420 ( .A(n298), .Y(n299) );
  AND2X2 U421 ( .A(n110), .B(\mem<19><9> ), .Y(n300) );
  INVX1 U422 ( .A(n300), .Y(n301) );
  AND2X2 U423 ( .A(\mem<19><10> ), .B(n2448), .Y(n302) );
  INVX1 U424 ( .A(n302), .Y(n303) );
  AND2X2 U425 ( .A(\mem<19><11> ), .B(n2448), .Y(n304) );
  INVX1 U426 ( .A(n304), .Y(n305) );
  AND2X2 U427 ( .A(\mem<19><12> ), .B(n2448), .Y(n306) );
  INVX1 U428 ( .A(n306), .Y(n307) );
  AND2X2 U429 ( .A(n2448), .B(\mem<19><13> ), .Y(n308) );
  INVX1 U430 ( .A(n308), .Y(n309) );
  AND2X2 U431 ( .A(\mem<19><14> ), .B(n2448), .Y(n310) );
  INVX1 U432 ( .A(n310), .Y(n311) );
  AND2X2 U433 ( .A(\mem<19><15> ), .B(n2448), .Y(n312) );
  INVX1 U434 ( .A(n312), .Y(n313) );
  AND2X2 U435 ( .A(n43), .B(\mem<18><0> ), .Y(n314) );
  INVX1 U436 ( .A(n314), .Y(n315) );
  AND2X2 U437 ( .A(n43), .B(\mem<18><1> ), .Y(n316) );
  INVX1 U438 ( .A(n316), .Y(n317) );
  AND2X2 U439 ( .A(n43), .B(\mem<18><2> ), .Y(n318) );
  INVX1 U440 ( .A(n318), .Y(n319) );
  AND2X2 U441 ( .A(n43), .B(\mem<18><3> ), .Y(n320) );
  INVX1 U442 ( .A(n320), .Y(n321) );
  AND2X2 U443 ( .A(n43), .B(\mem<18><4> ), .Y(n322) );
  INVX1 U444 ( .A(n322), .Y(n323) );
  AND2X2 U445 ( .A(n43), .B(\mem<18><5> ), .Y(n324) );
  INVX1 U446 ( .A(n324), .Y(n325) );
  AND2X2 U447 ( .A(n43), .B(\mem<18><6> ), .Y(n326) );
  INVX1 U448 ( .A(n326), .Y(n327) );
  AND2X2 U449 ( .A(n43), .B(\mem<18><7> ), .Y(n328) );
  INVX1 U450 ( .A(n328), .Y(n329) );
  AND2X2 U451 ( .A(n43), .B(\mem<18><8> ), .Y(n330) );
  INVX1 U452 ( .A(n330), .Y(n331) );
  AND2X2 U453 ( .A(n43), .B(\mem<18><9> ), .Y(n332) );
  INVX1 U454 ( .A(n332), .Y(n333) );
  AND2X2 U455 ( .A(n43), .B(\mem<18><10> ), .Y(n334) );
  INVX1 U456 ( .A(n334), .Y(n335) );
  AND2X2 U457 ( .A(n43), .B(\mem<18><11> ), .Y(n336) );
  INVX1 U458 ( .A(n336), .Y(n337) );
  AND2X2 U459 ( .A(n43), .B(\mem<18><12> ), .Y(n338) );
  INVX1 U460 ( .A(n338), .Y(n339) );
  AND2X2 U461 ( .A(n43), .B(\mem<18><13> ), .Y(n340) );
  INVX1 U462 ( .A(n340), .Y(n341) );
  AND2X2 U463 ( .A(n43), .B(\mem<18><14> ), .Y(n342) );
  INVX1 U464 ( .A(n342), .Y(n343) );
  AND2X2 U465 ( .A(n43), .B(\mem<18><15> ), .Y(n344) );
  INVX1 U466 ( .A(n344), .Y(n345) );
  AND2X2 U467 ( .A(n109), .B(\mem<17><0> ), .Y(n346) );
  INVX1 U468 ( .A(n346), .Y(n347) );
  AND2X2 U469 ( .A(n109), .B(\mem<17><1> ), .Y(n348) );
  INVX1 U470 ( .A(n348), .Y(n349) );
  AND2X2 U471 ( .A(\mem<17><2> ), .B(n2449), .Y(n350) );
  INVX1 U472 ( .A(n350), .Y(n351) );
  AND2X2 U473 ( .A(\mem<17><3> ), .B(n2449), .Y(n352) );
  INVX1 U474 ( .A(n352), .Y(n353) );
  AND2X2 U475 ( .A(\mem<17><4> ), .B(n2449), .Y(n354) );
  INVX1 U476 ( .A(n354), .Y(n355) );
  AND2X2 U477 ( .A(n109), .B(\mem<17><5> ), .Y(n356) );
  INVX1 U478 ( .A(n356), .Y(n357) );
  AND2X2 U479 ( .A(\mem<17><6> ), .B(n2449), .Y(n358) );
  INVX1 U480 ( .A(n358), .Y(n359) );
  AND2X2 U481 ( .A(\mem<17><7> ), .B(n2449), .Y(n360) );
  INVX1 U482 ( .A(n360), .Y(n361) );
  AND2X2 U483 ( .A(n2449), .B(\mem<17><8> ), .Y(n362) );
  INVX1 U484 ( .A(n362), .Y(n363) );
  AND2X2 U485 ( .A(n2449), .B(\mem<17><9> ), .Y(n364) );
  INVX1 U486 ( .A(n364), .Y(n365) );
  AND2X2 U487 ( .A(\mem<17><10> ), .B(n2449), .Y(n366) );
  INVX1 U488 ( .A(n366), .Y(n367) );
  AND2X2 U489 ( .A(\mem<17><11> ), .B(n2449), .Y(n368) );
  INVX1 U490 ( .A(n368), .Y(n369) );
  AND2X2 U491 ( .A(\mem<17><12> ), .B(n2449), .Y(n370) );
  INVX1 U492 ( .A(n370), .Y(n371) );
  AND2X2 U493 ( .A(n109), .B(\mem<17><13> ), .Y(n372) );
  INVX1 U494 ( .A(n372), .Y(n373) );
  AND2X2 U495 ( .A(\mem<17><14> ), .B(n2449), .Y(n374) );
  INVX1 U496 ( .A(n374), .Y(n375) );
  AND2X2 U497 ( .A(\mem<17><15> ), .B(n2449), .Y(n376) );
  INVX1 U498 ( .A(n376), .Y(n377) );
  AND2X2 U499 ( .A(n46), .B(\mem<16><0> ), .Y(n378) );
  INVX1 U500 ( .A(n378), .Y(n379) );
  AND2X2 U501 ( .A(n45), .B(\mem<16><1> ), .Y(n380) );
  INVX1 U502 ( .A(n380), .Y(n381) );
  AND2X2 U503 ( .A(\mem<16><2> ), .B(n46), .Y(n382) );
  INVX1 U504 ( .A(n382), .Y(n383) );
  AND2X2 U505 ( .A(n45), .B(\mem<16><3> ), .Y(n384) );
  INVX1 U506 ( .A(n384), .Y(n385) );
  AND2X2 U507 ( .A(\mem<16><4> ), .B(n46), .Y(n386) );
  INVX1 U508 ( .A(n386), .Y(n387) );
  AND2X2 U509 ( .A(n45), .B(\mem<16><5> ), .Y(n388) );
  INVX1 U510 ( .A(n388), .Y(n389) );
  AND2X2 U511 ( .A(\mem<16><6> ), .B(n46), .Y(n390) );
  INVX1 U512 ( .A(n390), .Y(n391) );
  AND2X2 U513 ( .A(n45), .B(\mem<16><7> ), .Y(n392) );
  INVX1 U514 ( .A(n392), .Y(n393) );
  AND2X2 U515 ( .A(n45), .B(\mem<16><8> ), .Y(n394) );
  INVX1 U516 ( .A(n394), .Y(n395) );
  AND2X2 U517 ( .A(n45), .B(\mem<16><9> ), .Y(n396) );
  INVX1 U518 ( .A(n396), .Y(n397) );
  AND2X2 U519 ( .A(\mem<16><10> ), .B(n46), .Y(n398) );
  INVX1 U520 ( .A(n398), .Y(n399) );
  AND2X2 U521 ( .A(n45), .B(\mem<16><11> ), .Y(n400) );
  INVX1 U522 ( .A(n400), .Y(n401) );
  AND2X2 U523 ( .A(\mem<16><12> ), .B(n46), .Y(n402) );
  INVX1 U524 ( .A(n402), .Y(n403) );
  AND2X2 U525 ( .A(n45), .B(\mem<16><13> ), .Y(n404) );
  INVX1 U526 ( .A(n404), .Y(n405) );
  AND2X2 U527 ( .A(\mem<16><14> ), .B(n46), .Y(n406) );
  INVX1 U528 ( .A(n406), .Y(n407) );
  AND2X2 U529 ( .A(n45), .B(\mem<16><15> ), .Y(n408) );
  INVX1 U530 ( .A(n408), .Y(n409) );
  AND2X2 U531 ( .A(n49), .B(\mem<15><0> ), .Y(n410) );
  INVX1 U532 ( .A(n410), .Y(n411) );
  AND2X2 U533 ( .A(n49), .B(\mem<15><1> ), .Y(n412) );
  INVX1 U534 ( .A(n412), .Y(n413) );
  AND2X2 U535 ( .A(n49), .B(\mem<15><2> ), .Y(n414) );
  INVX1 U536 ( .A(n414), .Y(n415) );
  AND2X2 U537 ( .A(n49), .B(\mem<15><3> ), .Y(n416) );
  INVX1 U538 ( .A(n416), .Y(n417) );
  AND2X2 U539 ( .A(n49), .B(\mem<15><4> ), .Y(n418) );
  INVX1 U540 ( .A(n418), .Y(n419) );
  AND2X2 U541 ( .A(n49), .B(\mem<15><5> ), .Y(n420) );
  INVX1 U542 ( .A(n420), .Y(n421) );
  AND2X2 U543 ( .A(n49), .B(\mem<15><6> ), .Y(n422) );
  INVX1 U544 ( .A(n422), .Y(n423) );
  AND2X2 U545 ( .A(n49), .B(\mem<15><7> ), .Y(n424) );
  INVX1 U546 ( .A(n424), .Y(n425) );
  AND2X2 U547 ( .A(n48), .B(\mem<15><8> ), .Y(n426) );
  INVX1 U548 ( .A(n426), .Y(n427) );
  AND2X2 U549 ( .A(n48), .B(\mem<15><9> ), .Y(n428) );
  INVX1 U550 ( .A(n428), .Y(n429) );
  AND2X2 U551 ( .A(n48), .B(\mem<15><10> ), .Y(n430) );
  INVX1 U552 ( .A(n430), .Y(n431) );
  AND2X2 U553 ( .A(n48), .B(\mem<15><11> ), .Y(n432) );
  INVX1 U554 ( .A(n432), .Y(n433) );
  AND2X2 U555 ( .A(n48), .B(\mem<15><12> ), .Y(n434) );
  INVX1 U556 ( .A(n434), .Y(n435) );
  AND2X2 U557 ( .A(n48), .B(\mem<15><13> ), .Y(n436) );
  INVX1 U558 ( .A(n436), .Y(n437) );
  AND2X2 U559 ( .A(n48), .B(\mem<15><14> ), .Y(n438) );
  INVX1 U560 ( .A(n438), .Y(n439) );
  AND2X2 U561 ( .A(n48), .B(\mem<15><15> ), .Y(n440) );
  INVX1 U562 ( .A(n440), .Y(n441) );
  AND2X2 U563 ( .A(n52), .B(\mem<14><0> ), .Y(n442) );
  INVX1 U564 ( .A(n442), .Y(n443) );
  AND2X2 U565 ( .A(n52), .B(\mem<14><1> ), .Y(n444) );
  INVX1 U566 ( .A(n444), .Y(n445) );
  AND2X2 U567 ( .A(n52), .B(\mem<14><2> ), .Y(n446) );
  INVX1 U568 ( .A(n446), .Y(n447) );
  AND2X2 U569 ( .A(n52), .B(\mem<14><3> ), .Y(n448) );
  INVX1 U570 ( .A(n448), .Y(n449) );
  AND2X2 U571 ( .A(n52), .B(\mem<14><4> ), .Y(n450) );
  INVX1 U572 ( .A(n450), .Y(n451) );
  AND2X2 U573 ( .A(n52), .B(\mem<14><5> ), .Y(n452) );
  INVX1 U574 ( .A(n452), .Y(n453) );
  AND2X2 U575 ( .A(n52), .B(\mem<14><6> ), .Y(n454) );
  INVX1 U576 ( .A(n454), .Y(n455) );
  AND2X2 U577 ( .A(n52), .B(\mem<14><7> ), .Y(n456) );
  INVX1 U578 ( .A(n456), .Y(n457) );
  AND2X2 U579 ( .A(n51), .B(\mem<14><8> ), .Y(n458) );
  INVX1 U580 ( .A(n458), .Y(n459) );
  AND2X2 U581 ( .A(n51), .B(\mem<14><9> ), .Y(n460) );
  INVX1 U582 ( .A(n460), .Y(n461) );
  AND2X2 U583 ( .A(n51), .B(\mem<14><10> ), .Y(n462) );
  INVX1 U584 ( .A(n462), .Y(n463) );
  AND2X2 U585 ( .A(n51), .B(\mem<14><11> ), .Y(n464) );
  INVX1 U586 ( .A(n464), .Y(n465) );
  AND2X2 U587 ( .A(n51), .B(\mem<14><12> ), .Y(n466) );
  INVX1 U588 ( .A(n466), .Y(n467) );
  AND2X2 U589 ( .A(n51), .B(\mem<14><13> ), .Y(n468) );
  INVX1 U590 ( .A(n468), .Y(n469) );
  AND2X2 U591 ( .A(n51), .B(\mem<14><14> ), .Y(n470) );
  INVX1 U592 ( .A(n470), .Y(n471) );
  AND2X2 U593 ( .A(n51), .B(\mem<14><15> ), .Y(n472) );
  INVX1 U594 ( .A(n472), .Y(n473) );
  AND2X2 U595 ( .A(n108), .B(\mem<13><0> ), .Y(n474) );
  INVX1 U596 ( .A(n474), .Y(n475) );
  AND2X2 U597 ( .A(n108), .B(\mem<13><1> ), .Y(n476) );
  INVX1 U598 ( .A(n476), .Y(n477) );
  AND2X2 U599 ( .A(\mem<13><2> ), .B(n2451), .Y(n478) );
  INVX1 U600 ( .A(n478), .Y(n479) );
  AND2X2 U601 ( .A(\mem<13><3> ), .B(n2451), .Y(n480) );
  INVX1 U602 ( .A(n480), .Y(n481) );
  AND2X2 U603 ( .A(\mem<13><4> ), .B(n2451), .Y(n482) );
  INVX1 U604 ( .A(n482), .Y(n483) );
  AND2X2 U605 ( .A(n108), .B(\mem<13><5> ), .Y(n484) );
  INVX1 U606 ( .A(n484), .Y(n485) );
  AND2X2 U607 ( .A(\mem<13><6> ), .B(n2451), .Y(n486) );
  INVX1 U608 ( .A(n486), .Y(n487) );
  AND2X2 U609 ( .A(\mem<13><7> ), .B(n2451), .Y(n488) );
  INVX1 U610 ( .A(n488), .Y(n489) );
  AND2X2 U611 ( .A(n2451), .B(\mem<13><8> ), .Y(n490) );
  INVX1 U612 ( .A(n490), .Y(n491) );
  AND2X2 U613 ( .A(n108), .B(\mem<13><9> ), .Y(n492) );
  INVX1 U614 ( .A(n492), .Y(n493) );
  AND2X2 U615 ( .A(\mem<13><10> ), .B(n2451), .Y(n494) );
  INVX1 U616 ( .A(n494), .Y(n495) );
  AND2X2 U617 ( .A(\mem<13><11> ), .B(n2451), .Y(n496) );
  INVX1 U618 ( .A(n496), .Y(n497) );
  AND2X2 U619 ( .A(\mem<13><12> ), .B(n2451), .Y(n498) );
  INVX1 U620 ( .A(n498), .Y(n499) );
  AND2X2 U621 ( .A(n2451), .B(\mem<13><13> ), .Y(n500) );
  INVX1 U622 ( .A(n500), .Y(n501) );
  AND2X2 U623 ( .A(\mem<13><14> ), .B(n2451), .Y(n502) );
  INVX1 U624 ( .A(n502), .Y(n503) );
  AND2X2 U625 ( .A(\mem<13><15> ), .B(n2451), .Y(n504) );
  INVX1 U626 ( .A(n504), .Y(n505) );
  AND2X2 U627 ( .A(n55), .B(\mem<12><0> ), .Y(n506) );
  INVX1 U628 ( .A(n506), .Y(n507) );
  AND2X2 U629 ( .A(n55), .B(\mem<12><1> ), .Y(n508) );
  INVX1 U630 ( .A(n508), .Y(n509) );
  AND2X2 U631 ( .A(n55), .B(\mem<12><2> ), .Y(n510) );
  INVX1 U632 ( .A(n510), .Y(n511) );
  AND2X2 U633 ( .A(n55), .B(\mem<12><3> ), .Y(n512) );
  INVX1 U634 ( .A(n512), .Y(n513) );
  AND2X2 U635 ( .A(n55), .B(\mem<12><4> ), .Y(n514) );
  INVX1 U636 ( .A(n514), .Y(n515) );
  AND2X2 U637 ( .A(n55), .B(\mem<12><5> ), .Y(n516) );
  INVX1 U638 ( .A(n516), .Y(n517) );
  AND2X2 U639 ( .A(n55), .B(\mem<12><6> ), .Y(n518) );
  INVX1 U640 ( .A(n518), .Y(n519) );
  AND2X2 U641 ( .A(n55), .B(\mem<12><7> ), .Y(n520) );
  INVX1 U642 ( .A(n520), .Y(n521) );
  AND2X2 U643 ( .A(n54), .B(\mem<12><8> ), .Y(n522) );
  INVX1 U644 ( .A(n522), .Y(n523) );
  AND2X2 U645 ( .A(n54), .B(\mem<12><9> ), .Y(n524) );
  INVX1 U646 ( .A(n524), .Y(n525) );
  AND2X2 U647 ( .A(n54), .B(\mem<12><10> ), .Y(n526) );
  INVX1 U648 ( .A(n526), .Y(n527) );
  AND2X2 U649 ( .A(n54), .B(\mem<12><11> ), .Y(n528) );
  INVX1 U650 ( .A(n528), .Y(n529) );
  AND2X2 U651 ( .A(n54), .B(\mem<12><12> ), .Y(n530) );
  INVX1 U652 ( .A(n530), .Y(n531) );
  AND2X2 U653 ( .A(n54), .B(\mem<12><13> ), .Y(n532) );
  INVX1 U654 ( .A(n532), .Y(n533) );
  AND2X2 U655 ( .A(n54), .B(\mem<12><14> ), .Y(n534) );
  INVX1 U656 ( .A(n534), .Y(n535) );
  AND2X2 U657 ( .A(n54), .B(\mem<12><15> ), .Y(n536) );
  INVX1 U658 ( .A(n536), .Y(n537) );
  AND2X2 U659 ( .A(n58), .B(\mem<11><0> ), .Y(n538) );
  INVX1 U660 ( .A(n538), .Y(n539) );
  AND2X2 U661 ( .A(n58), .B(\mem<11><1> ), .Y(n540) );
  INVX1 U662 ( .A(n540), .Y(n541) );
  AND2X2 U663 ( .A(n58), .B(\mem<11><2> ), .Y(n542) );
  INVX1 U664 ( .A(n542), .Y(n543) );
  AND2X2 U665 ( .A(n58), .B(\mem<11><3> ), .Y(n544) );
  INVX1 U666 ( .A(n544), .Y(n545) );
  AND2X2 U667 ( .A(n58), .B(\mem<11><4> ), .Y(n546) );
  INVX1 U668 ( .A(n546), .Y(n547) );
  AND2X2 U669 ( .A(n58), .B(\mem<11><5> ), .Y(n548) );
  INVX1 U670 ( .A(n548), .Y(n549) );
  AND2X2 U671 ( .A(n58), .B(\mem<11><6> ), .Y(n550) );
  INVX1 U672 ( .A(n550), .Y(n551) );
  AND2X2 U673 ( .A(n58), .B(\mem<11><7> ), .Y(n552) );
  INVX1 U674 ( .A(n552), .Y(n553) );
  AND2X2 U675 ( .A(n57), .B(\mem<11><8> ), .Y(n554) );
  INVX1 U676 ( .A(n554), .Y(n555) );
  AND2X2 U677 ( .A(n57), .B(\mem<11><9> ), .Y(n556) );
  INVX1 U678 ( .A(n556), .Y(n557) );
  AND2X2 U679 ( .A(n57), .B(\mem<11><10> ), .Y(n558) );
  INVX1 U680 ( .A(n558), .Y(n559) );
  AND2X2 U681 ( .A(n57), .B(\mem<11><11> ), .Y(n560) );
  INVX1 U682 ( .A(n560), .Y(n561) );
  AND2X2 U683 ( .A(n57), .B(\mem<11><12> ), .Y(n562) );
  INVX1 U684 ( .A(n562), .Y(n563) );
  AND2X2 U685 ( .A(n57), .B(\mem<11><13> ), .Y(n564) );
  INVX1 U686 ( .A(n564), .Y(n565) );
  AND2X2 U687 ( .A(n57), .B(\mem<11><14> ), .Y(n566) );
  INVX1 U688 ( .A(n566), .Y(n567) );
  AND2X2 U689 ( .A(n57), .B(\mem<11><15> ), .Y(n568) );
  INVX1 U690 ( .A(n568), .Y(n569) );
  AND2X2 U691 ( .A(n61), .B(\mem<10><0> ), .Y(n570) );
  INVX1 U692 ( .A(n570), .Y(n571) );
  AND2X2 U693 ( .A(n61), .B(\mem<10><1> ), .Y(n572) );
  INVX1 U694 ( .A(n572), .Y(n573) );
  AND2X2 U695 ( .A(n61), .B(\mem<10><2> ), .Y(n574) );
  INVX1 U696 ( .A(n574), .Y(n575) );
  AND2X2 U697 ( .A(n61), .B(\mem<10><3> ), .Y(n576) );
  INVX1 U698 ( .A(n576), .Y(n577) );
  AND2X2 U699 ( .A(n61), .B(\mem<10><4> ), .Y(n578) );
  INVX1 U700 ( .A(n578), .Y(n579) );
  AND2X2 U701 ( .A(n61), .B(\mem<10><5> ), .Y(n580) );
  INVX1 U702 ( .A(n580), .Y(n581) );
  AND2X2 U703 ( .A(n61), .B(\mem<10><6> ), .Y(n582) );
  INVX1 U704 ( .A(n582), .Y(n583) );
  AND2X2 U705 ( .A(n61), .B(\mem<10><7> ), .Y(n584) );
  INVX1 U706 ( .A(n584), .Y(n585) );
  AND2X2 U707 ( .A(n60), .B(\mem<10><8> ), .Y(n586) );
  INVX1 U708 ( .A(n586), .Y(n587) );
  AND2X2 U709 ( .A(n60), .B(\mem<10><9> ), .Y(n588) );
  INVX1 U710 ( .A(n588), .Y(n589) );
  AND2X2 U711 ( .A(n60), .B(\mem<10><10> ), .Y(n590) );
  INVX1 U712 ( .A(n590), .Y(n591) );
  AND2X2 U713 ( .A(n60), .B(\mem<10><11> ), .Y(n592) );
  INVX1 U714 ( .A(n592), .Y(n593) );
  AND2X2 U715 ( .A(n60), .B(\mem<10><12> ), .Y(n594) );
  INVX1 U716 ( .A(n594), .Y(n595) );
  AND2X2 U717 ( .A(n60), .B(\mem<10><13> ), .Y(n596) );
  INVX1 U718 ( .A(n596), .Y(n597) );
  AND2X2 U719 ( .A(n60), .B(\mem<10><14> ), .Y(n598) );
  INVX1 U720 ( .A(n598), .Y(n599) );
  AND2X2 U721 ( .A(n60), .B(\mem<10><15> ), .Y(n600) );
  INVX1 U722 ( .A(n600), .Y(n601) );
  AND2X2 U723 ( .A(n64), .B(\mem<9><0> ), .Y(n602) );
  INVX1 U724 ( .A(n602), .Y(n603) );
  AND2X2 U725 ( .A(n64), .B(\mem<9><1> ), .Y(n604) );
  INVX1 U726 ( .A(n604), .Y(n605) );
  AND2X2 U727 ( .A(n64), .B(\mem<9><2> ), .Y(n606) );
  INVX1 U728 ( .A(n606), .Y(n607) );
  AND2X2 U729 ( .A(n64), .B(\mem<9><3> ), .Y(n608) );
  INVX1 U730 ( .A(n608), .Y(n609) );
  AND2X2 U731 ( .A(n64), .B(\mem<9><4> ), .Y(n610) );
  INVX1 U732 ( .A(n610), .Y(n611) );
  AND2X2 U733 ( .A(n64), .B(\mem<9><5> ), .Y(n612) );
  INVX1 U734 ( .A(n612), .Y(n613) );
  AND2X2 U735 ( .A(n64), .B(\mem<9><6> ), .Y(n614) );
  INVX1 U736 ( .A(n614), .Y(n615) );
  AND2X2 U737 ( .A(n64), .B(\mem<9><7> ), .Y(n616) );
  INVX1 U738 ( .A(n616), .Y(n617) );
  AND2X2 U739 ( .A(n63), .B(\mem<9><8> ), .Y(n618) );
  INVX1 U740 ( .A(n618), .Y(n619) );
  AND2X2 U741 ( .A(n63), .B(\mem<9><9> ), .Y(n620) );
  INVX1 U742 ( .A(n620), .Y(n621) );
  AND2X2 U743 ( .A(n63), .B(\mem<9><10> ), .Y(n622) );
  INVX1 U744 ( .A(n622), .Y(n623) );
  AND2X2 U745 ( .A(n63), .B(\mem<9><11> ), .Y(n624) );
  INVX1 U746 ( .A(n624), .Y(n625) );
  AND2X2 U747 ( .A(n63), .B(\mem<9><12> ), .Y(n626) );
  INVX1 U748 ( .A(n626), .Y(n627) );
  AND2X2 U749 ( .A(n63), .B(\mem<9><13> ), .Y(n628) );
  INVX1 U750 ( .A(n628), .Y(n629) );
  AND2X2 U751 ( .A(n63), .B(\mem<9><14> ), .Y(n630) );
  INVX1 U752 ( .A(n630), .Y(n631) );
  AND2X2 U753 ( .A(n63), .B(\mem<9><15> ), .Y(n632) );
  INVX1 U754 ( .A(n632), .Y(n633) );
  AND2X2 U755 ( .A(n67), .B(\mem<8><0> ), .Y(n634) );
  INVX1 U756 ( .A(n634), .Y(n635) );
  AND2X2 U757 ( .A(n66), .B(\mem<8><1> ), .Y(n636) );
  INVX1 U758 ( .A(n636), .Y(n637) );
  AND2X2 U759 ( .A(\mem<8><2> ), .B(n67), .Y(n638) );
  INVX1 U760 ( .A(n638), .Y(n639) );
  AND2X2 U761 ( .A(n66), .B(\mem<8><3> ), .Y(n640) );
  INVX1 U762 ( .A(n640), .Y(n641) );
  AND2X2 U763 ( .A(\mem<8><4> ), .B(n67), .Y(n642) );
  INVX1 U764 ( .A(n642), .Y(n643) );
  AND2X2 U765 ( .A(n66), .B(\mem<8><5> ), .Y(n644) );
  INVX1 U766 ( .A(n644), .Y(n645) );
  AND2X2 U767 ( .A(\mem<8><6> ), .B(n67), .Y(n646) );
  INVX1 U768 ( .A(n646), .Y(n647) );
  AND2X2 U769 ( .A(n66), .B(\mem<8><7> ), .Y(n648) );
  INVX1 U770 ( .A(n648), .Y(n649) );
  AND2X2 U771 ( .A(n66), .B(\mem<8><8> ), .Y(n650) );
  INVX1 U772 ( .A(n650), .Y(n1163) );
  AND2X2 U773 ( .A(n66), .B(\mem<8><9> ), .Y(n1164) );
  INVX1 U774 ( .A(n1164), .Y(n1165) );
  AND2X2 U775 ( .A(\mem<8><10> ), .B(n67), .Y(n1166) );
  INVX1 U776 ( .A(n1166), .Y(n1167) );
  AND2X2 U777 ( .A(n66), .B(\mem<8><11> ), .Y(n1168) );
  INVX1 U778 ( .A(n1168), .Y(n1169) );
  AND2X2 U779 ( .A(\mem<8><12> ), .B(n67), .Y(n1170) );
  INVX1 U780 ( .A(n1170), .Y(n1171) );
  AND2X2 U781 ( .A(n66), .B(\mem<8><13> ), .Y(n1172) );
  INVX1 U782 ( .A(n1172), .Y(n1173) );
  AND2X2 U783 ( .A(\mem<8><14> ), .B(n67), .Y(n1174) );
  INVX1 U784 ( .A(n1174), .Y(n1175) );
  AND2X2 U785 ( .A(n66), .B(\mem<8><15> ), .Y(n1176) );
  INVX1 U786 ( .A(n1176), .Y(n1177) );
  AND2X2 U787 ( .A(n70), .B(\mem<7><1> ), .Y(n1178) );
  INVX1 U788 ( .A(n1178), .Y(n1179) );
  AND2X2 U789 ( .A(n70), .B(\mem<7><2> ), .Y(n1180) );
  INVX1 U790 ( .A(n1180), .Y(n1181) );
  AND2X2 U791 ( .A(n70), .B(\mem<7><3> ), .Y(n1182) );
  INVX1 U792 ( .A(n1182), .Y(n1183) );
  AND2X2 U793 ( .A(n70), .B(\mem<7><4> ), .Y(n1184) );
  INVX1 U794 ( .A(n1184), .Y(n1185) );
  AND2X2 U795 ( .A(n70), .B(\mem<7><5> ), .Y(n1186) );
  INVX1 U796 ( .A(n1186), .Y(n1187) );
  AND2X2 U797 ( .A(n70), .B(\mem<7><6> ), .Y(n1188) );
  INVX1 U798 ( .A(n1188), .Y(n1189) );
  AND2X2 U799 ( .A(n70), .B(\mem<7><7> ), .Y(n1190) );
  INVX1 U800 ( .A(n1190), .Y(n1191) );
  AND2X2 U801 ( .A(n69), .B(\mem<7><8> ), .Y(n1192) );
  INVX1 U802 ( .A(n1192), .Y(n1193) );
  AND2X2 U803 ( .A(n69), .B(\mem<7><9> ), .Y(n1194) );
  INVX1 U804 ( .A(n1194), .Y(n1195) );
  AND2X2 U805 ( .A(n69), .B(\mem<7><10> ), .Y(n1196) );
  INVX1 U806 ( .A(n1196), .Y(n1197) );
  AND2X2 U807 ( .A(n69), .B(\mem<7><11> ), .Y(n1198) );
  INVX1 U808 ( .A(n1198), .Y(n1199) );
  AND2X2 U809 ( .A(n69), .B(\mem<7><12> ), .Y(n1200) );
  INVX1 U810 ( .A(n1200), .Y(n1201) );
  AND2X2 U811 ( .A(n69), .B(\mem<7><13> ), .Y(n1202) );
  INVX1 U812 ( .A(n1202), .Y(n1203) );
  AND2X2 U813 ( .A(n69), .B(\mem<7><14> ), .Y(n1204) );
  INVX1 U814 ( .A(n1204), .Y(n1205) );
  AND2X2 U815 ( .A(n69), .B(\mem<7><15> ), .Y(n1206) );
  INVX1 U816 ( .A(n1206), .Y(n1207) );
  AND2X2 U817 ( .A(n73), .B(\mem<6><1> ), .Y(n1208) );
  INVX1 U818 ( .A(n1208), .Y(n1209) );
  AND2X2 U819 ( .A(n73), .B(\mem<6><2> ), .Y(n1210) );
  INVX1 U820 ( .A(n1210), .Y(n1211) );
  AND2X2 U821 ( .A(n73), .B(\mem<6><3> ), .Y(n1212) );
  INVX1 U822 ( .A(n1212), .Y(n1213) );
  AND2X2 U823 ( .A(n73), .B(\mem<6><4> ), .Y(n1214) );
  INVX1 U824 ( .A(n1214), .Y(n1215) );
  AND2X2 U825 ( .A(n73), .B(\mem<6><5> ), .Y(n1216) );
  INVX1 U826 ( .A(n1216), .Y(n1217) );
  AND2X2 U827 ( .A(n73), .B(\mem<6><6> ), .Y(n1218) );
  INVX1 U828 ( .A(n1218), .Y(n1219) );
  AND2X2 U829 ( .A(n73), .B(\mem<6><7> ), .Y(n1220) );
  INVX1 U830 ( .A(n1220), .Y(n1221) );
  AND2X2 U831 ( .A(n72), .B(\mem<6><8> ), .Y(n1222) );
  INVX1 U832 ( .A(n1222), .Y(n1223) );
  AND2X2 U833 ( .A(n72), .B(\mem<6><9> ), .Y(n1224) );
  INVX1 U834 ( .A(n1224), .Y(n1225) );
  AND2X2 U835 ( .A(n72), .B(\mem<6><10> ), .Y(n1226) );
  INVX1 U836 ( .A(n1226), .Y(n1227) );
  AND2X2 U837 ( .A(n72), .B(\mem<6><11> ), .Y(n1228) );
  INVX1 U838 ( .A(n1228), .Y(n1229) );
  AND2X2 U839 ( .A(n72), .B(\mem<6><12> ), .Y(n1230) );
  INVX1 U840 ( .A(n1230), .Y(n1231) );
  AND2X2 U841 ( .A(n72), .B(\mem<6><13> ), .Y(n1232) );
  INVX1 U842 ( .A(n1232), .Y(n1233) );
  AND2X2 U843 ( .A(n72), .B(\mem<6><14> ), .Y(n1234) );
  INVX1 U844 ( .A(n1234), .Y(n1235) );
  AND2X2 U845 ( .A(n72), .B(\mem<6><15> ), .Y(n1236) );
  INVX1 U846 ( .A(n1236), .Y(n1237) );
  AND2X2 U847 ( .A(n76), .B(\mem<5><1> ), .Y(n1238) );
  INVX1 U848 ( .A(n1238), .Y(n1239) );
  AND2X2 U849 ( .A(n76), .B(\mem<5><2> ), .Y(n1240) );
  INVX1 U850 ( .A(n1240), .Y(n1241) );
  AND2X2 U851 ( .A(n76), .B(\mem<5><3> ), .Y(n1242) );
  INVX1 U852 ( .A(n1242), .Y(n1243) );
  AND2X2 U853 ( .A(n76), .B(\mem<5><4> ), .Y(n1244) );
  INVX1 U854 ( .A(n1244), .Y(n1245) );
  AND2X2 U855 ( .A(n76), .B(\mem<5><5> ), .Y(n1246) );
  INVX1 U856 ( .A(n1246), .Y(n1247) );
  AND2X2 U857 ( .A(n76), .B(\mem<5><6> ), .Y(n1248) );
  INVX1 U858 ( .A(n1248), .Y(n1249) );
  AND2X2 U859 ( .A(n76), .B(\mem<5><7> ), .Y(n1250) );
  INVX1 U860 ( .A(n1250), .Y(n1251) );
  AND2X2 U861 ( .A(n75), .B(\mem<5><8> ), .Y(n1252) );
  INVX1 U862 ( .A(n1252), .Y(n1253) );
  AND2X2 U863 ( .A(n75), .B(\mem<5><9> ), .Y(n1254) );
  INVX1 U864 ( .A(n1254), .Y(n1255) );
  AND2X2 U865 ( .A(n75), .B(\mem<5><10> ), .Y(n1256) );
  INVX1 U866 ( .A(n1256), .Y(n1257) );
  AND2X2 U867 ( .A(n75), .B(\mem<5><11> ), .Y(n1258) );
  INVX1 U868 ( .A(n1258), .Y(n1259) );
  AND2X2 U869 ( .A(n75), .B(\mem<5><12> ), .Y(n1260) );
  INVX1 U870 ( .A(n1260), .Y(n1261) );
  AND2X2 U871 ( .A(n75), .B(\mem<5><13> ), .Y(n1262) );
  INVX1 U872 ( .A(n1262), .Y(n1263) );
  AND2X2 U873 ( .A(n75), .B(\mem<5><14> ), .Y(n1264) );
  INVX1 U874 ( .A(n1264), .Y(n1265) );
  AND2X2 U875 ( .A(n75), .B(\mem<5><15> ), .Y(n1266) );
  INVX1 U876 ( .A(n1266), .Y(n1267) );
  AND2X2 U877 ( .A(n79), .B(\mem<4><1> ), .Y(n1268) );
  INVX1 U878 ( .A(n1268), .Y(n1269) );
  AND2X2 U879 ( .A(n79), .B(\mem<4><2> ), .Y(n1270) );
  INVX1 U880 ( .A(n1270), .Y(n1271) );
  AND2X2 U881 ( .A(n79), .B(\mem<4><3> ), .Y(n1272) );
  INVX1 U882 ( .A(n1272), .Y(n1273) );
  AND2X2 U883 ( .A(n79), .B(\mem<4><4> ), .Y(n1274) );
  INVX1 U884 ( .A(n1274), .Y(n1275) );
  AND2X2 U885 ( .A(n79), .B(\mem<4><5> ), .Y(n1276) );
  INVX1 U886 ( .A(n1276), .Y(n1277) );
  AND2X2 U887 ( .A(n79), .B(\mem<4><6> ), .Y(n1278) );
  INVX1 U888 ( .A(n1278), .Y(n1279) );
  AND2X2 U889 ( .A(n79), .B(\mem<4><7> ), .Y(n1280) );
  INVX1 U890 ( .A(n1280), .Y(n1281) );
  AND2X2 U891 ( .A(n78), .B(\mem<4><8> ), .Y(n1282) );
  INVX1 U892 ( .A(n1282), .Y(n1283) );
  AND2X2 U893 ( .A(n78), .B(\mem<4><9> ), .Y(n1284) );
  INVX1 U894 ( .A(n1284), .Y(n1285) );
  AND2X2 U895 ( .A(n78), .B(\mem<4><10> ), .Y(n1286) );
  INVX1 U896 ( .A(n1286), .Y(n1287) );
  AND2X2 U897 ( .A(n78), .B(\mem<4><11> ), .Y(n1288) );
  INVX1 U898 ( .A(n1288), .Y(n1289) );
  AND2X2 U899 ( .A(n78), .B(\mem<4><12> ), .Y(n1290) );
  INVX1 U900 ( .A(n1290), .Y(n1291) );
  AND2X2 U901 ( .A(n78), .B(\mem<4><13> ), .Y(n1292) );
  INVX1 U902 ( .A(n1292), .Y(n1293) );
  AND2X2 U903 ( .A(n78), .B(\mem<4><14> ), .Y(n1294) );
  INVX1 U904 ( .A(n1294), .Y(n1295) );
  AND2X2 U905 ( .A(n78), .B(\mem<4><15> ), .Y(n1296) );
  INVX1 U906 ( .A(n1296), .Y(n1297) );
  AND2X2 U907 ( .A(n81), .B(\mem<3><1> ), .Y(n1298) );
  INVX1 U908 ( .A(n1298), .Y(n1299) );
  AND2X2 U909 ( .A(n81), .B(\mem<3><2> ), .Y(n1300) );
  INVX1 U910 ( .A(n1300), .Y(n1301) );
  AND2X2 U911 ( .A(n81), .B(\mem<3><3> ), .Y(n1302) );
  INVX1 U912 ( .A(n1302), .Y(n1303) );
  AND2X2 U913 ( .A(n81), .B(\mem<3><4> ), .Y(n1304) );
  INVX1 U914 ( .A(n1304), .Y(n1305) );
  AND2X2 U915 ( .A(\mem<3><5> ), .B(n82), .Y(n1306) );
  INVX1 U916 ( .A(n1306), .Y(n1307) );
  AND2X2 U917 ( .A(n81), .B(\mem<3><6> ), .Y(n1308) );
  INVX1 U918 ( .A(n1308), .Y(n1309) );
  AND2X2 U919 ( .A(\mem<3><7> ), .B(n82), .Y(n1310) );
  INVX1 U920 ( .A(n1310), .Y(n1311) );
  AND2X2 U921 ( .A(n81), .B(\mem<3><8> ), .Y(n1312) );
  INVX1 U922 ( .A(n1312), .Y(n1313) );
  AND2X2 U923 ( .A(n81), .B(\mem<3><9> ), .Y(n1314) );
  INVX1 U924 ( .A(n1314), .Y(n1315) );
  AND2X2 U925 ( .A(n82), .B(\mem<3><10> ), .Y(n1316) );
  INVX1 U926 ( .A(n1316), .Y(n1317) );
  AND2X2 U927 ( .A(n82), .B(\mem<3><11> ), .Y(n1318) );
  INVX1 U928 ( .A(n1318), .Y(n1319) );
  AND2X2 U929 ( .A(\mem<3><12> ), .B(n82), .Y(n1320) );
  INVX1 U930 ( .A(n1320), .Y(n1321) );
  AND2X2 U931 ( .A(n81), .B(\mem<3><13> ), .Y(n1322) );
  INVX1 U932 ( .A(n1322), .Y(n1323) );
  AND2X2 U933 ( .A(n81), .B(\mem<3><14> ), .Y(n1324) );
  INVX1 U934 ( .A(n1324), .Y(n1325) );
  AND2X2 U935 ( .A(\mem<3><15> ), .B(n82), .Y(n1326) );
  INVX1 U936 ( .A(n1326), .Y(n1327) );
  AND2X2 U937 ( .A(n84), .B(\mem<2><1> ), .Y(n1328) );
  INVX1 U938 ( .A(n1328), .Y(n1329) );
  AND2X2 U939 ( .A(n84), .B(\mem<2><2> ), .Y(n1330) );
  INVX1 U940 ( .A(n1330), .Y(n1331) );
  AND2X2 U941 ( .A(n84), .B(\mem<2><3> ), .Y(n1332) );
  INVX1 U942 ( .A(n1332), .Y(n1333) );
  AND2X2 U943 ( .A(n84), .B(\mem<2><4> ), .Y(n1334) );
  INVX1 U944 ( .A(n1334), .Y(n1335) );
  AND2X2 U945 ( .A(\mem<2><5> ), .B(n85), .Y(n1336) );
  INVX1 U946 ( .A(n1336), .Y(n1337) );
  AND2X2 U947 ( .A(n84), .B(\mem<2><6> ), .Y(n1338) );
  INVX1 U948 ( .A(n1338), .Y(n1339) );
  AND2X2 U949 ( .A(\mem<2><7> ), .B(n85), .Y(n1340) );
  INVX1 U950 ( .A(n1340), .Y(n1341) );
  AND2X2 U951 ( .A(n84), .B(\mem<2><8> ), .Y(n1342) );
  INVX1 U952 ( .A(n1342), .Y(n1343) );
  AND2X2 U953 ( .A(n84), .B(\mem<2><9> ), .Y(n1344) );
  INVX1 U954 ( .A(n1344), .Y(n1345) );
  AND2X2 U955 ( .A(n85), .B(\mem<2><10> ), .Y(n1346) );
  INVX1 U956 ( .A(n1346), .Y(n1347) );
  AND2X2 U957 ( .A(\mem<2><11> ), .B(n85), .Y(n1348) );
  INVX1 U958 ( .A(n1348), .Y(n1349) );
  AND2X2 U959 ( .A(\mem<2><12> ), .B(n85), .Y(n1350) );
  INVX1 U960 ( .A(n1350), .Y(n1351) );
  AND2X2 U961 ( .A(n84), .B(\mem<2><13> ), .Y(n1352) );
  INVX1 U962 ( .A(n1352), .Y(n1353) );
  AND2X2 U963 ( .A(n84), .B(\mem<2><14> ), .Y(n1354) );
  INVX1 U964 ( .A(n1354), .Y(n1355) );
  AND2X2 U965 ( .A(\mem<2><15> ), .B(n85), .Y(n1356) );
  INVX1 U966 ( .A(n1356), .Y(n1357) );
  AND2X2 U967 ( .A(n87), .B(\mem<1><1> ), .Y(n1358) );
  INVX1 U968 ( .A(n1358), .Y(n1359) );
  AND2X2 U969 ( .A(n87), .B(\mem<1><2> ), .Y(n1360) );
  INVX1 U970 ( .A(n1360), .Y(n1361) );
  AND2X2 U971 ( .A(n87), .B(\mem<1><3> ), .Y(n1362) );
  INVX1 U972 ( .A(n1362), .Y(n1363) );
  AND2X2 U973 ( .A(\mem<1><4> ), .B(n88), .Y(n1364) );
  INVX1 U974 ( .A(n1364), .Y(n1365) );
  AND2X2 U975 ( .A(\mem<1><5> ), .B(n88), .Y(n1366) );
  INVX1 U976 ( .A(n1366), .Y(n1367) );
  AND2X2 U977 ( .A(n87), .B(\mem<1><6> ), .Y(n1368) );
  INVX1 U978 ( .A(n1368), .Y(n1369) );
  AND2X2 U979 ( .A(\mem<1><7> ), .B(n88), .Y(n1370) );
  INVX1 U980 ( .A(n1370), .Y(n1371) );
  AND2X2 U981 ( .A(n87), .B(\mem<1><8> ), .Y(n1372) );
  INVX1 U982 ( .A(n1372), .Y(n1373) );
  AND2X2 U983 ( .A(n87), .B(\mem<1><9> ), .Y(n1374) );
  INVX1 U984 ( .A(n1374), .Y(n1375) );
  AND2X2 U985 ( .A(n87), .B(\mem<1><10> ), .Y(n1376) );
  INVX1 U986 ( .A(n1376), .Y(n1377) );
  AND2X2 U987 ( .A(\mem<1><11> ), .B(n88), .Y(n1378) );
  INVX1 U988 ( .A(n1378), .Y(n1379) );
  AND2X2 U989 ( .A(\mem<1><12> ), .B(n88), .Y(n1380) );
  INVX1 U990 ( .A(n1380), .Y(n1381) );
  AND2X2 U991 ( .A(n87), .B(\mem<1><13> ), .Y(n1382) );
  INVX1 U992 ( .A(n1382), .Y(n1383) );
  AND2X2 U993 ( .A(n87), .B(\mem<1><14> ), .Y(n1384) );
  INVX1 U994 ( .A(n1384), .Y(n1385) );
  AND2X2 U995 ( .A(\mem<1><15> ), .B(n88), .Y(n1386) );
  INVX1 U996 ( .A(n1386), .Y(n1387) );
  AND2X2 U997 ( .A(n90), .B(\mem<0><1> ), .Y(n1388) );
  INVX1 U998 ( .A(n1388), .Y(n1389) );
  AND2X2 U999 ( .A(n91), .B(\mem<0><2> ), .Y(n1390) );
  INVX1 U1000 ( .A(n1390), .Y(n1391) );
  AND2X2 U1001 ( .A(n90), .B(\mem<0><3> ), .Y(n1392) );
  INVX1 U1002 ( .A(n1392), .Y(n1393) );
  AND2X2 U1003 ( .A(\mem<0><4> ), .B(n91), .Y(n1394) );
  INVX1 U1004 ( .A(n1394), .Y(n1395) );
  AND2X2 U1005 ( .A(n90), .B(\mem<0><5> ), .Y(n1396) );
  INVX1 U1006 ( .A(n1396), .Y(n1397) );
  AND2X2 U1007 ( .A(\mem<0><6> ), .B(n91), .Y(n1398) );
  INVX1 U1008 ( .A(n1398), .Y(n1399) );
  AND2X2 U1009 ( .A(n90), .B(\mem<0><7> ), .Y(n1400) );
  INVX1 U1010 ( .A(n1400), .Y(n1401) );
  AND2X2 U1011 ( .A(n90), .B(\mem<0><8> ), .Y(n1402) );
  INVX1 U1012 ( .A(n1402), .Y(n1403) );
  AND2X2 U1013 ( .A(n90), .B(\mem<0><9> ), .Y(n1404) );
  INVX1 U1014 ( .A(n1404), .Y(n1405) );
  AND2X2 U1015 ( .A(\mem<0><10> ), .B(n91), .Y(n1406) );
  INVX1 U1016 ( .A(n1406), .Y(n1407) );
  AND2X2 U1017 ( .A(n90), .B(\mem<0><11> ), .Y(n1408) );
  INVX1 U1018 ( .A(n1408), .Y(n1409) );
  AND2X2 U1019 ( .A(\mem<0><12> ), .B(n91), .Y(n1410) );
  INVX1 U1020 ( .A(n1410), .Y(n1411) );
  AND2X2 U1021 ( .A(n90), .B(\mem<0><13> ), .Y(n1412) );
  INVX1 U1022 ( .A(n1412), .Y(n1413) );
  AND2X2 U1023 ( .A(\mem<0><14> ), .B(n91), .Y(n1414) );
  INVX1 U1024 ( .A(n1414), .Y(n1415) );
  AND2X2 U1025 ( .A(n90), .B(\mem<0><15> ), .Y(n1416) );
  INVX1 U1026 ( .A(n1416), .Y(n1417) );
  INVX1 U1027 ( .A(n2426), .Y(n2425) );
  INVX1 U1028 ( .A(n2423), .Y(n2422) );
  AND2X1 U1029 ( .A(n2425), .B(n2292), .Y(n1419) );
  AND2X1 U1030 ( .A(n2974), .B(n2429), .Y(n1420) );
  AND2X2 U1031 ( .A(\mem<31><1> ), .B(n121), .Y(n1421) );
  INVX1 U1032 ( .A(n1421), .Y(n1422) );
  AND2X2 U1033 ( .A(\mem<31><2> ), .B(n121), .Y(n1423) );
  INVX1 U1034 ( .A(n1423), .Y(n1424) );
  AND2X2 U1035 ( .A(\mem<31><3> ), .B(n121), .Y(n1425) );
  INVX1 U1036 ( .A(n1425), .Y(n1426) );
  AND2X2 U1037 ( .A(\mem<31><4> ), .B(n2432), .Y(n1427) );
  INVX1 U1038 ( .A(n1427), .Y(n1428) );
  AND2X2 U1039 ( .A(\mem<31><5> ), .B(n121), .Y(n1429) );
  INVX1 U1040 ( .A(n1429), .Y(n1430) );
  AND2X2 U1041 ( .A(\mem<31><6> ), .B(n2432), .Y(n1431) );
  INVX1 U1042 ( .A(n1431), .Y(n1432) );
  AND2X2 U1043 ( .A(\mem<31><7> ), .B(n121), .Y(n1433) );
  INVX1 U1044 ( .A(n1433), .Y(n1434) );
  AND2X2 U1045 ( .A(\mem<31><8> ), .B(n121), .Y(n1435) );
  INVX1 U1046 ( .A(n1435), .Y(n1436) );
  AND2X2 U1047 ( .A(\mem<31><9> ), .B(n121), .Y(n1437) );
  INVX1 U1048 ( .A(n1437), .Y(n1438) );
  AND2X2 U1049 ( .A(\mem<31><10> ), .B(n2432), .Y(n1439) );
  INVX1 U1050 ( .A(n1439), .Y(n1440) );
  AND2X2 U1051 ( .A(\mem<31><11> ), .B(n2432), .Y(n1441) );
  INVX1 U1052 ( .A(n1441), .Y(n1442) );
  AND2X2 U1053 ( .A(\mem<31><12> ), .B(n121), .Y(n1443) );
  INVX1 U1054 ( .A(n1443), .Y(n1444) );
  AND2X2 U1055 ( .A(\mem<31><13> ), .B(n2432), .Y(n1445) );
  INVX1 U1056 ( .A(n1445), .Y(n1446) );
  AND2X2 U1057 ( .A(\mem<31><14> ), .B(n2432), .Y(n1447) );
  INVX1 U1058 ( .A(n1447), .Y(n1448) );
  AND2X2 U1059 ( .A(\mem<31><15> ), .B(n2432), .Y(n1449) );
  INVX1 U1060 ( .A(n1449), .Y(n1450) );
  AND2X2 U1061 ( .A(n120), .B(\mem<30><1> ), .Y(n1451) );
  INVX1 U1062 ( .A(n1451), .Y(n1452) );
  AND2X2 U1063 ( .A(\mem<30><2> ), .B(n2433), .Y(n1453) );
  INVX1 U1064 ( .A(n1453), .Y(n1454) );
  AND2X2 U1065 ( .A(n120), .B(\mem<30><3> ), .Y(n1455) );
  INVX1 U1066 ( .A(n1455), .Y(n1456) );
  AND2X2 U1067 ( .A(\mem<30><4> ), .B(n2433), .Y(n1457) );
  INVX1 U1068 ( .A(n1457), .Y(n1458) );
  AND2X2 U1069 ( .A(n120), .B(\mem<30><5> ), .Y(n1459) );
  INVX1 U1070 ( .A(n1459), .Y(n1460) );
  AND2X2 U1071 ( .A(\mem<30><6> ), .B(n2433), .Y(n1461) );
  INVX1 U1072 ( .A(n1461), .Y(n1462) );
  AND2X2 U1073 ( .A(n120), .B(\mem<30><7> ), .Y(n1463) );
  INVX1 U1074 ( .A(n1463), .Y(n1464) );
  AND2X2 U1075 ( .A(\mem<30><8> ), .B(n2433), .Y(n1465) );
  INVX1 U1076 ( .A(n1465), .Y(n1466) );
  AND2X2 U1077 ( .A(\mem<30><9> ), .B(n2433), .Y(n1467) );
  INVX1 U1078 ( .A(n1467), .Y(n1468) );
  AND2X2 U1079 ( .A(\mem<30><10> ), .B(n2433), .Y(n1469) );
  INVX1 U1080 ( .A(n1469), .Y(n1470) );
  AND2X2 U1081 ( .A(\mem<30><11> ), .B(n2433), .Y(n1471) );
  INVX1 U1082 ( .A(n1471), .Y(n1472) );
  AND2X2 U1083 ( .A(\mem<30><12> ), .B(n2433), .Y(n1473) );
  INVX1 U1084 ( .A(n1473), .Y(n1474) );
  AND2X2 U1085 ( .A(\mem<30><13> ), .B(n2433), .Y(n1475) );
  INVX1 U1086 ( .A(n1475), .Y(n1476) );
  AND2X2 U1087 ( .A(\mem<30><14> ), .B(n2433), .Y(n1477) );
  INVX1 U1088 ( .A(n1477), .Y(n1478) );
  AND2X2 U1089 ( .A(\mem<30><15> ), .B(n2433), .Y(n1479) );
  INVX1 U1090 ( .A(n1479), .Y(n1480) );
  AND2X2 U1091 ( .A(n119), .B(\mem<29><1> ), .Y(n1481) );
  INVX1 U1092 ( .A(n1481), .Y(n1482) );
  AND2X2 U1093 ( .A(\mem<29><2> ), .B(n2435), .Y(n1483) );
  INVX1 U1094 ( .A(n1483), .Y(n1484) );
  AND2X2 U1095 ( .A(n119), .B(\mem<29><3> ), .Y(n1485) );
  INVX1 U1096 ( .A(n1485), .Y(n1486) );
  AND2X2 U1097 ( .A(\mem<29><4> ), .B(n2435), .Y(n1487) );
  INVX1 U1098 ( .A(n1487), .Y(n1488) );
  AND2X2 U1099 ( .A(n119), .B(\mem<29><5> ), .Y(n1489) );
  INVX1 U1100 ( .A(n1489), .Y(n1490) );
  AND2X2 U1101 ( .A(\mem<29><6> ), .B(n2435), .Y(n1491) );
  INVX1 U1102 ( .A(n1491), .Y(n1492) );
  AND2X2 U1103 ( .A(n119), .B(\mem<29><7> ), .Y(n1493) );
  INVX1 U1104 ( .A(n1493), .Y(n1494) );
  AND2X2 U1105 ( .A(\mem<29><8> ), .B(n2435), .Y(n1495) );
  INVX1 U1106 ( .A(n1495), .Y(n1496) );
  AND2X2 U1107 ( .A(\mem<29><9> ), .B(n2435), .Y(n1497) );
  INVX1 U1108 ( .A(n1497), .Y(n1498) );
  AND2X2 U1109 ( .A(\mem<29><10> ), .B(n2435), .Y(n1499) );
  INVX1 U1110 ( .A(n1499), .Y(n1500) );
  AND2X2 U1111 ( .A(\mem<29><11> ), .B(n2435), .Y(n1501) );
  INVX1 U1112 ( .A(n1501), .Y(n1502) );
  AND2X2 U1113 ( .A(\mem<29><12> ), .B(n2435), .Y(n1503) );
  INVX1 U1114 ( .A(n1503), .Y(n1504) );
  AND2X2 U1115 ( .A(\mem<29><13> ), .B(n2435), .Y(n1505) );
  INVX1 U1116 ( .A(n1505), .Y(n1506) );
  AND2X2 U1117 ( .A(\mem<29><14> ), .B(n2435), .Y(n1507) );
  INVX1 U1118 ( .A(n1507), .Y(n1508) );
  AND2X2 U1119 ( .A(\mem<29><15> ), .B(n2435), .Y(n1509) );
  INVX1 U1120 ( .A(n1509), .Y(n1510) );
  AND2X2 U1121 ( .A(\mem<28><1> ), .B(n2437), .Y(n1511) );
  INVX1 U1122 ( .A(n1511), .Y(n1512) );
  AND2X2 U1123 ( .A(\mem<28><2> ), .B(n2437), .Y(n1513) );
  INVX1 U1124 ( .A(n1513), .Y(n1514) );
  AND2X2 U1125 ( .A(\mem<28><3> ), .B(n2437), .Y(n1515) );
  INVX1 U1126 ( .A(n1515), .Y(n1516) );
  AND2X2 U1127 ( .A(n118), .B(\mem<28><4> ), .Y(n1517) );
  INVX1 U1128 ( .A(n1517), .Y(n1518) );
  AND2X2 U1129 ( .A(n118), .B(\mem<28><5> ), .Y(n1519) );
  INVX1 U1130 ( .A(n1519), .Y(n1520) );
  AND2X2 U1131 ( .A(n118), .B(\mem<28><6> ), .Y(n1521) );
  INVX1 U1132 ( .A(n1521), .Y(n1522) );
  AND2X2 U1133 ( .A(n118), .B(\mem<28><7> ), .Y(n1523) );
  INVX1 U1134 ( .A(n1523), .Y(n1524) );
  AND2X2 U1135 ( .A(\mem<28><8> ), .B(n2437), .Y(n1525) );
  INVX1 U1136 ( .A(n1525), .Y(n1526) );
  AND2X2 U1137 ( .A(\mem<28><9> ), .B(n2437), .Y(n1527) );
  INVX1 U1138 ( .A(n1527), .Y(n1528) );
  AND2X2 U1139 ( .A(\mem<28><10> ), .B(n2437), .Y(n1529) );
  INVX1 U1140 ( .A(n1529), .Y(n1530) );
  AND2X2 U1141 ( .A(\mem<28><11> ), .B(n2437), .Y(n1531) );
  INVX1 U1142 ( .A(n1531), .Y(n1532) );
  AND2X2 U1143 ( .A(\mem<28><12> ), .B(n2437), .Y(n1533) );
  INVX1 U1144 ( .A(n1533), .Y(n1534) );
  AND2X2 U1145 ( .A(\mem<28><13> ), .B(n2437), .Y(n1535) );
  INVX1 U1146 ( .A(n1535), .Y(n1536) );
  AND2X2 U1147 ( .A(\mem<28><14> ), .B(n2437), .Y(n1537) );
  INVX1 U1148 ( .A(n1537), .Y(n1538) );
  AND2X2 U1149 ( .A(\mem<28><15> ), .B(n2437), .Y(n1539) );
  INVX1 U1150 ( .A(n1539), .Y(n1540) );
  AND2X2 U1151 ( .A(\mem<27><1> ), .B(n2439), .Y(n1541) );
  INVX1 U1152 ( .A(n1541), .Y(n1542) );
  AND2X2 U1153 ( .A(\mem<27><2> ), .B(n2439), .Y(n1543) );
  INVX1 U1154 ( .A(n1543), .Y(n1544) );
  AND2X2 U1155 ( .A(\mem<27><3> ), .B(n2439), .Y(n1545) );
  INVX1 U1156 ( .A(n1545), .Y(n1546) );
  AND2X2 U1157 ( .A(n117), .B(\mem<27><4> ), .Y(n1547) );
  INVX1 U1158 ( .A(n1547), .Y(n1548) );
  AND2X2 U1159 ( .A(\mem<27><5> ), .B(n2439), .Y(n1549) );
  INVX1 U1160 ( .A(n1549), .Y(n1550) );
  AND2X2 U1161 ( .A(\mem<27><6> ), .B(n2439), .Y(n1551) );
  INVX1 U1162 ( .A(n1551), .Y(n1552) );
  AND2X2 U1163 ( .A(n117), .B(\mem<27><7> ), .Y(n1553) );
  INVX1 U1164 ( .A(n1553), .Y(n1554) );
  AND2X2 U1165 ( .A(\mem<27><8> ), .B(n2439), .Y(n1555) );
  INVX1 U1166 ( .A(n1555), .Y(n1556) );
  AND2X2 U1167 ( .A(\mem<27><9> ), .B(n2439), .Y(n1557) );
  INVX1 U1168 ( .A(n1557), .Y(n1558) );
  AND2X2 U1169 ( .A(\mem<27><10> ), .B(n2439), .Y(n1559) );
  INVX1 U1170 ( .A(n1559), .Y(n1560) );
  AND2X2 U1171 ( .A(n117), .B(\mem<27><11> ), .Y(n1561) );
  INVX1 U1172 ( .A(n1561), .Y(n1562) );
  AND2X2 U1173 ( .A(\mem<27><12> ), .B(n2439), .Y(n1563) );
  INVX1 U1174 ( .A(n1563), .Y(n1564) );
  AND2X2 U1175 ( .A(\mem<27><13> ), .B(n2439), .Y(n1565) );
  INVX1 U1177 ( .A(n1565), .Y(n1566) );
  AND2X2 U1178 ( .A(\mem<27><14> ), .B(n2439), .Y(n1567) );
  INVX1 U1179 ( .A(n1567), .Y(n1568) );
  AND2X2 U1180 ( .A(n117), .B(\mem<27><15> ), .Y(n1569) );
  INVX1 U1181 ( .A(n1569), .Y(n1570) );
  AND2X2 U1182 ( .A(n116), .B(\mem<26><1> ), .Y(n1571) );
  INVX1 U1183 ( .A(n1571), .Y(n1572) );
  AND2X2 U1184 ( .A(\mem<26><2> ), .B(n2441), .Y(n1573) );
  INVX1 U1185 ( .A(n1573), .Y(n1574) );
  AND2X2 U1186 ( .A(\mem<26><3> ), .B(n2441), .Y(n1575) );
  INVX1 U1187 ( .A(n1575), .Y(n1576) );
  AND2X2 U1188 ( .A(\mem<26><4> ), .B(n2441), .Y(n1577) );
  INVX1 U1189 ( .A(n1577), .Y(n1578) );
  AND2X2 U1190 ( .A(n116), .B(\mem<26><5> ), .Y(n1579) );
  INVX1 U1191 ( .A(n1579), .Y(n1580) );
  AND2X2 U1192 ( .A(\mem<26><6> ), .B(n2441), .Y(n1581) );
  INVX1 U1193 ( .A(n1581), .Y(n1582) );
  AND2X2 U1194 ( .A(\mem<26><7> ), .B(n2441), .Y(n1583) );
  INVX1 U1195 ( .A(n1583), .Y(n1584) );
  AND2X2 U1196 ( .A(n2441), .B(\mem<26><8> ), .Y(n1585) );
  INVX1 U1197 ( .A(n1585), .Y(n1586) );
  AND2X2 U1198 ( .A(n116), .B(\mem<26><9> ), .Y(n1587) );
  INVX1 U1199 ( .A(n1587), .Y(n1588) );
  AND2X2 U1200 ( .A(\mem<26><10> ), .B(n2441), .Y(n1589) );
  INVX1 U1201 ( .A(n1589), .Y(n1590) );
  AND2X2 U1202 ( .A(\mem<26><11> ), .B(n2441), .Y(n1591) );
  INVX1 U1203 ( .A(n1591), .Y(n1592) );
  AND2X2 U1204 ( .A(\mem<26><12> ), .B(n2441), .Y(n1593) );
  INVX1 U1205 ( .A(n1593), .Y(n1594) );
  AND2X2 U1206 ( .A(n2441), .B(\mem<26><13> ), .Y(n1595) );
  INVX1 U1207 ( .A(n1595), .Y(n1596) );
  AND2X2 U1208 ( .A(\mem<26><14> ), .B(n2441), .Y(n1597) );
  INVX1 U1209 ( .A(n1597), .Y(n1598) );
  AND2X2 U1210 ( .A(\mem<26><15> ), .B(n2441), .Y(n1599) );
  INVX1 U1211 ( .A(n1599), .Y(n1600) );
  AND2X2 U1212 ( .A(n115), .B(\mem<25><1> ), .Y(n1601) );
  INVX1 U1213 ( .A(n1601), .Y(n1602) );
  AND2X2 U1214 ( .A(\mem<25><2> ), .B(n2443), .Y(n1603) );
  INVX1 U1215 ( .A(n1603), .Y(n1604) );
  AND2X2 U1216 ( .A(\mem<25><3> ), .B(n2443), .Y(n1605) );
  INVX1 U1217 ( .A(n1605), .Y(n1606) );
  AND2X2 U1218 ( .A(\mem<25><4> ), .B(n2443), .Y(n1607) );
  INVX1 U1219 ( .A(n1607), .Y(n1608) );
  AND2X2 U1220 ( .A(n115), .B(\mem<25><5> ), .Y(n1609) );
  INVX1 U1221 ( .A(n1609), .Y(n1610) );
  AND2X2 U1222 ( .A(\mem<25><6> ), .B(n2443), .Y(n1611) );
  INVX1 U1223 ( .A(n1611), .Y(n1612) );
  AND2X2 U1224 ( .A(\mem<25><7> ), .B(n2443), .Y(n1613) );
  INVX1 U1225 ( .A(n1613), .Y(n1614) );
  AND2X2 U1226 ( .A(n2443), .B(\mem<25><8> ), .Y(n1615) );
  INVX1 U1227 ( .A(n1615), .Y(n1616) );
  AND2X2 U1228 ( .A(n115), .B(\mem<25><9> ), .Y(n1617) );
  INVX1 U1229 ( .A(n1617), .Y(n1618) );
  AND2X2 U1230 ( .A(\mem<25><10> ), .B(n2443), .Y(n1619) );
  INVX1 U1231 ( .A(n1619), .Y(n1620) );
  AND2X2 U1232 ( .A(\mem<25><11> ), .B(n2443), .Y(n1621) );
  INVX1 U1233 ( .A(n1621), .Y(n1622) );
  AND2X2 U1234 ( .A(\mem<25><12> ), .B(n2443), .Y(n1623) );
  INVX1 U1235 ( .A(n1623), .Y(n1624) );
  AND2X2 U1236 ( .A(n2443), .B(\mem<25><13> ), .Y(n1625) );
  INVX1 U1237 ( .A(n1625), .Y(n1626) );
  AND2X2 U1238 ( .A(\mem<25><14> ), .B(n2443), .Y(n1627) );
  INVX1 U1239 ( .A(n1627), .Y(n1628) );
  AND2X2 U1240 ( .A(\mem<25><15> ), .B(n2443), .Y(n1629) );
  INVX1 U1241 ( .A(n1629), .Y(n1630) );
  AND2X2 U1242 ( .A(n41), .B(\mem<24><1> ), .Y(n1631) );
  INVX1 U1243 ( .A(n1631), .Y(n1632) );
  AND2X2 U1244 ( .A(\mem<24><2> ), .B(n41), .Y(n1633) );
  INVX1 U1245 ( .A(n1633), .Y(n1634) );
  AND2X2 U1246 ( .A(n41), .B(\mem<24><3> ), .Y(n1635) );
  INVX1 U1247 ( .A(n1635), .Y(n1636) );
  AND2X2 U1248 ( .A(\mem<24><4> ), .B(n41), .Y(n1637) );
  INVX1 U1249 ( .A(n1637), .Y(n1638) );
  AND2X2 U1250 ( .A(n41), .B(\mem<24><5> ), .Y(n1639) );
  INVX1 U1251 ( .A(n1639), .Y(n1640) );
  AND2X2 U1252 ( .A(\mem<24><6> ), .B(n41), .Y(n1641) );
  INVX1 U1253 ( .A(n1641), .Y(n1642) );
  AND2X2 U1254 ( .A(n41), .B(\mem<24><7> ), .Y(n1643) );
  INVX1 U1255 ( .A(n1643), .Y(n1644) );
  AND2X2 U1256 ( .A(n41), .B(\mem<24><8> ), .Y(n1645) );
  INVX1 U1257 ( .A(n1645), .Y(n1646) );
  AND2X2 U1258 ( .A(n41), .B(\mem<24><9> ), .Y(n1647) );
  INVX1 U1259 ( .A(n1647), .Y(n1648) );
  AND2X2 U1260 ( .A(\mem<24><10> ), .B(n41), .Y(n1649) );
  INVX1 U1261 ( .A(n1649), .Y(n1650) );
  AND2X2 U1262 ( .A(n41), .B(\mem<24><11> ), .Y(n1651) );
  INVX1 U1263 ( .A(n1651), .Y(n1652) );
  AND2X2 U1264 ( .A(\mem<24><12> ), .B(n41), .Y(n1653) );
  INVX1 U1265 ( .A(n1653), .Y(n1654) );
  AND2X2 U1266 ( .A(n41), .B(\mem<24><13> ), .Y(n1655) );
  INVX1 U1267 ( .A(n1655), .Y(n1656) );
  AND2X2 U1268 ( .A(\mem<24><14> ), .B(n41), .Y(n1657) );
  INVX1 U1269 ( .A(n1657), .Y(n1658) );
  AND2X2 U1270 ( .A(n41), .B(\mem<24><15> ), .Y(n1659) );
  INVX1 U1271 ( .A(n1659), .Y(n1660) );
  AND2X2 U1272 ( .A(n70), .B(\mem<7><0> ), .Y(n1661) );
  INVX1 U1273 ( .A(n1661), .Y(n1662) );
  AND2X2 U1274 ( .A(n73), .B(\mem<6><0> ), .Y(n1663) );
  INVX1 U1275 ( .A(n1663), .Y(n1664) );
  AND2X2 U1276 ( .A(n76), .B(\mem<5><0> ), .Y(n1665) );
  INVX1 U1277 ( .A(n1665), .Y(n1666) );
  AND2X2 U1278 ( .A(n79), .B(\mem<4><0> ), .Y(n1667) );
  INVX1 U1279 ( .A(n1667), .Y(n1668) );
  AND2X2 U1280 ( .A(\mem<3><0> ), .B(n82), .Y(n1669) );
  INVX1 U1281 ( .A(n1669), .Y(n1670) );
  AND2X2 U1282 ( .A(\mem<2><0> ), .B(n85), .Y(n1671) );
  INVX1 U1283 ( .A(n1671), .Y(n1672) );
  AND2X2 U1284 ( .A(\mem<1><0> ), .B(n88), .Y(n1673) );
  INVX1 U1285 ( .A(n1673), .Y(n1674) );
  AND2X2 U1286 ( .A(\mem<0><0> ), .B(n91), .Y(n1675) );
  INVX1 U1287 ( .A(n1675), .Y(n1676) );
  AND2X1 U1288 ( .A(N32), .B(n2421), .Y(n1677) );
  INVX1 U1289 ( .A(n1677), .Y(n1678) );
  AND2X1 U1290 ( .A(N31), .B(n2421), .Y(n1679) );
  AND2X1 U1291 ( .A(N30), .B(n2421), .Y(n1680) );
  INVX1 U1292 ( .A(n1680), .Y(n1681) );
  AND2X1 U1293 ( .A(N29), .B(n2421), .Y(n1682) );
  INVX1 U1294 ( .A(n1682), .Y(n1683) );
  AND2X1 U1295 ( .A(N28), .B(n2421), .Y(n1684) );
  INVX1 U1296 ( .A(n1684), .Y(n1685) );
  AND2X1 U1297 ( .A(N27), .B(n2421), .Y(n1686) );
  INVX1 U1298 ( .A(n1686), .Y(n1687) );
  AND2X1 U1299 ( .A(N26), .B(n2421), .Y(n1688) );
  INVX1 U1300 ( .A(n1688), .Y(n1689) );
  AND2X1 U1301 ( .A(N25), .B(n2421), .Y(n1690) );
  INVX1 U1302 ( .A(n1690), .Y(n1691) );
  AND2X1 U1303 ( .A(N24), .B(n2421), .Y(n1692) );
  INVX1 U1304 ( .A(n1692), .Y(n1693) );
  AND2X1 U1305 ( .A(N23), .B(n2421), .Y(n1694) );
  INVX1 U1306 ( .A(n1694), .Y(n1695) );
  AND2X1 U1307 ( .A(N22), .B(n2421), .Y(n1696) );
  AND2X1 U1308 ( .A(N21), .B(n2421), .Y(n1697) );
  INVX1 U1309 ( .A(n1697), .Y(n1698) );
  AND2X1 U1310 ( .A(N20), .B(n2421), .Y(n1699) );
  INVX1 U1311 ( .A(n1699), .Y(n1700) );
  AND2X1 U1312 ( .A(N19), .B(n2421), .Y(n1701) );
  INVX1 U1313 ( .A(n1701), .Y(n1702) );
  AND2X1 U1314 ( .A(N18), .B(n2421), .Y(n1703) );
  INVX1 U1315 ( .A(n1703), .Y(n1704) );
  AND2X1 U1316 ( .A(N17), .B(n2421), .Y(n1705) );
  INVX1 U1317 ( .A(n1705), .Y(n1706) );
  BUFX2 U1318 ( .A(n2434), .Y(n1707) );
  INVX1 U1319 ( .A(n1707), .Y(n2454) );
  BUFX2 U1320 ( .A(n2436), .Y(n1708) );
  INVX1 U1321 ( .A(n1708), .Y(n2455) );
  BUFX2 U1322 ( .A(n2438), .Y(n1709) );
  INVX1 U1323 ( .A(n1709), .Y(n2456) );
  BUFX2 U1324 ( .A(n2440), .Y(n1710) );
  INVX1 U1325 ( .A(n1710), .Y(n2457) );
  BUFX2 U1326 ( .A(n2442), .Y(n1711) );
  INVX1 U1327 ( .A(n1711), .Y(n2458) );
  BUFX2 U1328 ( .A(n2450), .Y(n1712) );
  INVX1 U1329 ( .A(n1712), .Y(n2452) );
  BUFX2 U1330 ( .A(n2453), .Y(n1713) );
  INVX1 U1331 ( .A(n1713), .Y(n2459) );
  AND2X1 U1332 ( .A(n2422), .B(n1419), .Y(n1714) );
  AND2X1 U1333 ( .A(n2427), .B(n1420), .Y(n1715) );
  AND2X1 U1334 ( .A(n2423), .B(n1419), .Y(n1716) );
  AND2X1 U1335 ( .A(n2428), .B(n1420), .Y(n1717) );
  INVX1 U1336 ( .A(n13), .Y(\data_out<0> ) );
  AND2X1 U1337 ( .A(n1715), .B(n2460), .Y(n1719) );
  AND2X1 U1338 ( .A(n2460), .B(n1717), .Y(n1720) );
  AND2X1 U1339 ( .A(n2460), .B(n2452), .Y(n1721) );
  AND2X1 U1340 ( .A(n2460), .B(n2459), .Y(n1722) );
  AND2X1 U1341 ( .A(n1714), .B(n1715), .Y(n1723) );
  INVX1 U1342 ( .A(n1723), .Y(n1724) );
  AND2X1 U1343 ( .A(n1715), .B(n1716), .Y(n1725) );
  INVX1 U1344 ( .A(n1725), .Y(n1726) );
  AND2X1 U1345 ( .A(n1715), .B(n2454), .Y(n1727) );
  INVX1 U1346 ( .A(n1727), .Y(n1728) );
  AND2X1 U1347 ( .A(n1715), .B(n2455), .Y(n1729) );
  INVX1 U1348 ( .A(n1729), .Y(n1730) );
  AND2X1 U1349 ( .A(n1715), .B(n2456), .Y(n1731) );
  INVX1 U1350 ( .A(n1731), .Y(n1732) );
  AND2X1 U1351 ( .A(n1715), .B(n2457), .Y(n1733) );
  INVX1 U1352 ( .A(n1733), .Y(n1734) );
  AND2X1 U1353 ( .A(n1715), .B(n2458), .Y(n1735) );
  INVX1 U1354 ( .A(n1735), .Y(n1736) );
  AND2X1 U1355 ( .A(n1714), .B(n1717), .Y(n1737) );
  INVX1 U1356 ( .A(n1737), .Y(n1738) );
  AND2X1 U1357 ( .A(n1716), .B(n1717), .Y(n1739) );
  INVX1 U1358 ( .A(n1739), .Y(n1740) );
  AND2X1 U1359 ( .A(n2454), .B(n1717), .Y(n1741) );
  INVX1 U1360 ( .A(n1741), .Y(n1742) );
  AND2X1 U1361 ( .A(n2455), .B(n1717), .Y(n1743) );
  INVX1 U1362 ( .A(n1743), .Y(n1744) );
  AND2X1 U1363 ( .A(n2456), .B(n1717), .Y(n1745) );
  INVX1 U1364 ( .A(n1745), .Y(n1746) );
  AND2X1 U1365 ( .A(n2457), .B(n1717), .Y(n1747) );
  INVX1 U1366 ( .A(n1747), .Y(n1748) );
  AND2X1 U1367 ( .A(n2458), .B(n1717), .Y(n1749) );
  INVX1 U1368 ( .A(n1749), .Y(n1750) );
  AND2X1 U1369 ( .A(n1714), .B(n2452), .Y(n1751) );
  INVX1 U1370 ( .A(n1751), .Y(n1752) );
  AND2X1 U1371 ( .A(n1716), .B(n2452), .Y(n1753) );
  INVX1 U1372 ( .A(n1753), .Y(n1754) );
  AND2X1 U1373 ( .A(n2454), .B(n2452), .Y(n1755) );
  INVX1 U1374 ( .A(n1755), .Y(n1756) );
  AND2X1 U1375 ( .A(n2455), .B(n2452), .Y(n1757) );
  INVX1 U1376 ( .A(n1757), .Y(n1758) );
  AND2X1 U1377 ( .A(n2456), .B(n2452), .Y(n1759) );
  INVX1 U1378 ( .A(n1759), .Y(n1760) );
  AND2X1 U1379 ( .A(n2457), .B(n2452), .Y(n1761) );
  INVX1 U1380 ( .A(n1761), .Y(n1762) );
  AND2X1 U1381 ( .A(n2458), .B(n2452), .Y(n1763) );
  INVX1 U1382 ( .A(n1763), .Y(n1764) );
  AND2X1 U1383 ( .A(n1714), .B(n2459), .Y(n1765) );
  INVX1 U1384 ( .A(n1765), .Y(n1766) );
  AND2X1 U1385 ( .A(n1716), .B(n2459), .Y(n1767) );
  INVX1 U1386 ( .A(n1767), .Y(n1768) );
  AND2X1 U1387 ( .A(n2454), .B(n2459), .Y(n1769) );
  INVX1 U1388 ( .A(n1769), .Y(n1770) );
  AND2X1 U1389 ( .A(n2455), .B(n2459), .Y(n1771) );
  INVX1 U1390 ( .A(n1771), .Y(n1772) );
  AND2X1 U1391 ( .A(n2456), .B(n2459), .Y(n1773) );
  INVX1 U1392 ( .A(n1773), .Y(n1774) );
  AND2X1 U1393 ( .A(n2457), .B(n2459), .Y(n1775) );
  INVX1 U1394 ( .A(n1775), .Y(n1776) );
  AND2X1 U1395 ( .A(n2458), .B(n2459), .Y(n1777) );
  INVX1 U1396 ( .A(n1777), .Y(n1778) );
  INVX1 U1397 ( .A(N11), .Y(n2424) );
  MUX2X1 U1398 ( .B(n1780), .A(n1781), .S(n2285), .Y(n1779) );
  MUX2X1 U1399 ( .B(n1783), .A(n1784), .S(n2285), .Y(n1782) );
  MUX2X1 U1400 ( .B(n1786), .A(n1787), .S(n2285), .Y(n1785) );
  MUX2X1 U1401 ( .B(n1789), .A(n1790), .S(n2285), .Y(n1788) );
  MUX2X1 U1402 ( .B(n1792), .A(n1793), .S(n2277), .Y(n1791) );
  MUX2X1 U1403 ( .B(n1795), .A(n1796), .S(n2285), .Y(n1794) );
  MUX2X1 U1404 ( .B(n1798), .A(n1799), .S(n2285), .Y(n1797) );
  MUX2X1 U1405 ( .B(n1801), .A(n1802), .S(n2285), .Y(n1800) );
  MUX2X1 U1406 ( .B(n1804), .A(n1805), .S(n2285), .Y(n1803) );
  MUX2X1 U1407 ( .B(n1807), .A(n1808), .S(n2277), .Y(n1806) );
  MUX2X1 U1408 ( .B(n1810), .A(n1811), .S(n2286), .Y(n1809) );
  MUX2X1 U1409 ( .B(n1813), .A(n1814), .S(n2286), .Y(n1812) );
  MUX2X1 U1410 ( .B(n1816), .A(n1817), .S(n2286), .Y(n1815) );
  MUX2X1 U1411 ( .B(n1819), .A(n1820), .S(n2286), .Y(n1818) );
  MUX2X1 U1412 ( .B(n1822), .A(n1823), .S(n2277), .Y(n1821) );
  MUX2X1 U1413 ( .B(n1825), .A(n1826), .S(n2286), .Y(n1824) );
  MUX2X1 U1414 ( .B(n1828), .A(n1829), .S(n2286), .Y(n1827) );
  MUX2X1 U1415 ( .B(n1831), .A(n1832), .S(n2286), .Y(n1830) );
  MUX2X1 U1416 ( .B(n1834), .A(n1835), .S(n2286), .Y(n1833) );
  MUX2X1 U1417 ( .B(n1837), .A(n1838), .S(n2277), .Y(n1836) );
  MUX2X1 U1418 ( .B(n1840), .A(n1841), .S(n2286), .Y(n1839) );
  MUX2X1 U1419 ( .B(n1843), .A(n1844), .S(n2286), .Y(n1842) );
  MUX2X1 U1420 ( .B(n1846), .A(n1847), .S(n2286), .Y(n1845) );
  MUX2X1 U1421 ( .B(n1849), .A(n1850), .S(n2286), .Y(n1848) );
  MUX2X1 U1422 ( .B(n1852), .A(n1853), .S(n2277), .Y(n1851) );
  MUX2X1 U1423 ( .B(n1855), .A(n1856), .S(n2287), .Y(n1854) );
  MUX2X1 U1424 ( .B(n1858), .A(n1859), .S(n2287), .Y(n1857) );
  MUX2X1 U1425 ( .B(n1861), .A(n1862), .S(n2287), .Y(n1860) );
  MUX2X1 U1426 ( .B(n1864), .A(n1865), .S(n2287), .Y(n1863) );
  MUX2X1 U1427 ( .B(n1867), .A(n1868), .S(n2277), .Y(n1866) );
  MUX2X1 U1428 ( .B(n1870), .A(n1871), .S(n2287), .Y(n1869) );
  MUX2X1 U1429 ( .B(n1873), .A(n1874), .S(n2287), .Y(n1872) );
  MUX2X1 U1430 ( .B(n1876), .A(n1877), .S(n2287), .Y(n1875) );
  MUX2X1 U1431 ( .B(n1879), .A(n1880), .S(n2287), .Y(n1878) );
  MUX2X1 U1432 ( .B(n1882), .A(n1883), .S(n2277), .Y(n1881) );
  MUX2X1 U1433 ( .B(n1885), .A(n1886), .S(n2287), .Y(n1884) );
  MUX2X1 U1434 ( .B(n1888), .A(n1889), .S(n2287), .Y(n1887) );
  MUX2X1 U1435 ( .B(n1891), .A(n1892), .S(n2287), .Y(n1890) );
  MUX2X1 U1436 ( .B(n1894), .A(n1895), .S(n2287), .Y(n1893) );
  MUX2X1 U1437 ( .B(n1897), .A(n1898), .S(n2277), .Y(n1896) );
  MUX2X1 U1438 ( .B(n1900), .A(n1901), .S(n2288), .Y(n1899) );
  MUX2X1 U1439 ( .B(n1903), .A(n1904), .S(n2288), .Y(n1902) );
  MUX2X1 U1440 ( .B(n1906), .A(n1907), .S(n2288), .Y(n1905) );
  MUX2X1 U1441 ( .B(n1909), .A(n1910), .S(n2288), .Y(n1908) );
  MUX2X1 U1442 ( .B(n1912), .A(n1913), .S(n2277), .Y(n1911) );
  MUX2X1 U1443 ( .B(n1915), .A(n1916), .S(n2288), .Y(n1914) );
  MUX2X1 U1444 ( .B(n1918), .A(n1919), .S(n2288), .Y(n1917) );
  MUX2X1 U1445 ( .B(n1921), .A(n1922), .S(n2288), .Y(n1920) );
  MUX2X1 U1446 ( .B(n1924), .A(n1925), .S(n2288), .Y(n1923) );
  MUX2X1 U1447 ( .B(n1927), .A(n1928), .S(n2277), .Y(n1926) );
  MUX2X1 U1448 ( .B(n1930), .A(n1931), .S(n2288), .Y(n1929) );
  MUX2X1 U1449 ( .B(n1933), .A(n1934), .S(n2288), .Y(n1932) );
  MUX2X1 U1450 ( .B(n1936), .A(n1937), .S(n2288), .Y(n1935) );
  MUX2X1 U1451 ( .B(n1939), .A(n1940), .S(n2288), .Y(n1938) );
  MUX2X1 U1452 ( .B(n1942), .A(n1943), .S(n2277), .Y(n1941) );
  MUX2X1 U1453 ( .B(n1945), .A(n1946), .S(n2289), .Y(n1944) );
  MUX2X1 U1454 ( .B(n1948), .A(n1949), .S(n2289), .Y(n1947) );
  MUX2X1 U1455 ( .B(n1951), .A(n1952), .S(n2289), .Y(n1950) );
  MUX2X1 U1456 ( .B(n1954), .A(n1955), .S(n2289), .Y(n1953) );
  MUX2X1 U1457 ( .B(n1957), .A(n1958), .S(n2277), .Y(n1956) );
  MUX2X1 U1458 ( .B(n1960), .A(n1961), .S(n2289), .Y(n1959) );
  MUX2X1 U1459 ( .B(n1963), .A(n1964), .S(n2289), .Y(n1962) );
  MUX2X1 U1460 ( .B(n1966), .A(n1967), .S(n2289), .Y(n1965) );
  MUX2X1 U1461 ( .B(n1969), .A(n1970), .S(n2289), .Y(n1968) );
  MUX2X1 U1462 ( .B(n1972), .A(n1973), .S(n2276), .Y(n1971) );
  MUX2X1 U1463 ( .B(n1975), .A(n1976), .S(n2289), .Y(n1974) );
  MUX2X1 U1464 ( .B(n1978), .A(n1979), .S(n2289), .Y(n1977) );
  MUX2X1 U1465 ( .B(n1981), .A(n1982), .S(n2289), .Y(n1980) );
  MUX2X1 U1466 ( .B(n1984), .A(n1985), .S(n2289), .Y(n1983) );
  MUX2X1 U1467 ( .B(n1987), .A(n1988), .S(n2276), .Y(n1986) );
  MUX2X1 U1468 ( .B(n1990), .A(n1991), .S(n2290), .Y(n1989) );
  MUX2X1 U1469 ( .B(n1993), .A(n1994), .S(n2290), .Y(n1992) );
  MUX2X1 U1470 ( .B(n1996), .A(n1997), .S(n2290), .Y(n1995) );
  MUX2X1 U1471 ( .B(n1999), .A(n2000), .S(n2290), .Y(n1998) );
  MUX2X1 U1472 ( .B(n2002), .A(n2003), .S(n2276), .Y(n2001) );
  MUX2X1 U1473 ( .B(n2005), .A(n2006), .S(n2290), .Y(n2004) );
  MUX2X1 U1474 ( .B(n2008), .A(n2009), .S(n2290), .Y(n2007) );
  MUX2X1 U1475 ( .B(n2011), .A(n2012), .S(n2290), .Y(n2010) );
  MUX2X1 U1476 ( .B(n2014), .A(n2015), .S(n2290), .Y(n2013) );
  MUX2X1 U1477 ( .B(n2017), .A(n2018), .S(n2276), .Y(n2016) );
  MUX2X1 U1478 ( .B(n2020), .A(n2021), .S(n2290), .Y(n2019) );
  MUX2X1 U1479 ( .B(n2023), .A(n2024), .S(n2290), .Y(n2022) );
  MUX2X1 U1480 ( .B(n2026), .A(n2027), .S(n2290), .Y(n2025) );
  MUX2X1 U1481 ( .B(n2029), .A(n2030), .S(n2290), .Y(n2028) );
  MUX2X1 U1482 ( .B(n2032), .A(n2033), .S(n2276), .Y(n2031) );
  MUX2X1 U1483 ( .B(n2035), .A(n2036), .S(n2291), .Y(n2034) );
  MUX2X1 U1484 ( .B(n2038), .A(n2039), .S(n2291), .Y(n2037) );
  MUX2X1 U1485 ( .B(n2041), .A(n2042), .S(n2291), .Y(n2040) );
  MUX2X1 U1486 ( .B(n2044), .A(n2045), .S(n2291), .Y(n2043) );
  MUX2X1 U1487 ( .B(n2047), .A(n2048), .S(n2276), .Y(n2046) );
  MUX2X1 U1488 ( .B(n2050), .A(n2051), .S(n2291), .Y(n2049) );
  MUX2X1 U1489 ( .B(n2053), .A(n2054), .S(n2291), .Y(n2052) );
  MUX2X1 U1490 ( .B(n2056), .A(n2057), .S(n2291), .Y(n2055) );
  MUX2X1 U1491 ( .B(n2059), .A(n2060), .S(n2291), .Y(n2058) );
  MUX2X1 U1492 ( .B(n2062), .A(n2063), .S(n2276), .Y(n2061) );
  MUX2X1 U1493 ( .B(n2065), .A(n2066), .S(n2291), .Y(n2064) );
  MUX2X1 U1494 ( .B(n2068), .A(n2069), .S(n2291), .Y(n2067) );
  MUX2X1 U1495 ( .B(n2071), .A(n2072), .S(n2291), .Y(n2070) );
  MUX2X1 U1496 ( .B(n2074), .A(n2075), .S(n2291), .Y(n2073) );
  MUX2X1 U1497 ( .B(n2077), .A(n2078), .S(n2276), .Y(n2076) );
  MUX2X1 U1498 ( .B(n2080), .A(n2081), .S(n2292), .Y(n2079) );
  MUX2X1 U1499 ( .B(n2083), .A(n2084), .S(n2292), .Y(n2082) );
  MUX2X1 U1500 ( .B(n2086), .A(n2087), .S(n2292), .Y(n2085) );
  MUX2X1 U1501 ( .B(n2089), .A(n2090), .S(n2292), .Y(n2088) );
  MUX2X1 U1502 ( .B(n2092), .A(n2093), .S(n2276), .Y(n2091) );
  MUX2X1 U1503 ( .B(n2095), .A(n2096), .S(n2292), .Y(n2094) );
  MUX2X1 U1504 ( .B(n2098), .A(n2099), .S(n2292), .Y(n2097) );
  MUX2X1 U1505 ( .B(n2101), .A(n2102), .S(n2292), .Y(n2100) );
  MUX2X1 U1506 ( .B(n2104), .A(n2105), .S(n2292), .Y(n2103) );
  MUX2X1 U1507 ( .B(n2107), .A(n2108), .S(n2276), .Y(n2106) );
  MUX2X1 U1508 ( .B(n2110), .A(n2111), .S(n2292), .Y(n2109) );
  MUX2X1 U1509 ( .B(n2113), .A(n2114), .S(n2292), .Y(n2112) );
  MUX2X1 U1510 ( .B(n2116), .A(n2117), .S(n2292), .Y(n2115) );
  MUX2X1 U1511 ( .B(n2119), .A(n2120), .S(n2292), .Y(n2118) );
  MUX2X1 U1512 ( .B(n2122), .A(n2123), .S(n2276), .Y(n2121) );
  MUX2X1 U1513 ( .B(n2125), .A(n2126), .S(n2293), .Y(n2124) );
  MUX2X1 U1514 ( .B(n2128), .A(n2129), .S(n2293), .Y(n2127) );
  MUX2X1 U1515 ( .B(n2131), .A(n2132), .S(n2293), .Y(n2130) );
  MUX2X1 U1516 ( .B(n2134), .A(n2135), .S(n2293), .Y(n2133) );
  MUX2X1 U1517 ( .B(n2137), .A(n2138), .S(n2276), .Y(n2136) );
  MUX2X1 U1518 ( .B(n2140), .A(n2141), .S(n2293), .Y(n2139) );
  MUX2X1 U1519 ( .B(n2143), .A(n2144), .S(n2293), .Y(n2142) );
  MUX2X1 U1520 ( .B(n2146), .A(n2147), .S(n2293), .Y(n2145) );
  MUX2X1 U1521 ( .B(n2149), .A(n2150), .S(n2293), .Y(n2148) );
  MUX2X1 U1522 ( .B(n2152), .A(n2153), .S(n2277), .Y(n2151) );
  MUX2X1 U1523 ( .B(n2155), .A(n2156), .S(n2293), .Y(n2154) );
  MUX2X1 U1524 ( .B(n2158), .A(n2159), .S(n2293), .Y(n2157) );
  MUX2X1 U1525 ( .B(n2161), .A(n2162), .S(n2293), .Y(n2160) );
  MUX2X1 U1526 ( .B(n2164), .A(n2165), .S(n2293), .Y(n2163) );
  MUX2X1 U1527 ( .B(n2167), .A(n2168), .S(n2427), .Y(n2166) );
  MUX2X1 U1528 ( .B(n2170), .A(n2171), .S(n2294), .Y(n2169) );
  MUX2X1 U1529 ( .B(n2173), .A(n2174), .S(n2294), .Y(n2172) );
  MUX2X1 U1530 ( .B(n2176), .A(n2177), .S(n2294), .Y(n2175) );
  MUX2X1 U1531 ( .B(n2179), .A(n2180), .S(n2294), .Y(n2178) );
  MUX2X1 U1532 ( .B(n2182), .A(n2183), .S(n2427), .Y(n2181) );
  MUX2X1 U1533 ( .B(n2185), .A(n2186), .S(n2294), .Y(n2184) );
  MUX2X1 U1534 ( .B(n2188), .A(n2189), .S(n2294), .Y(n2187) );
  MUX2X1 U1535 ( .B(n2191), .A(n2192), .S(n2294), .Y(n2190) );
  MUX2X1 U1536 ( .B(n2194), .A(n2195), .S(n2294), .Y(n2193) );
  MUX2X1 U1537 ( .B(n2197), .A(n2198), .S(n2277), .Y(n2196) );
  MUX2X1 U1538 ( .B(n2200), .A(n2201), .S(n2294), .Y(n2199) );
  MUX2X1 U1539 ( .B(n2203), .A(n2204), .S(n2294), .Y(n2202) );
  MUX2X1 U1540 ( .B(n2206), .A(n2207), .S(n2294), .Y(n2205) );
  MUX2X1 U1541 ( .B(n2209), .A(n2210), .S(n2294), .Y(n2208) );
  MUX2X1 U1542 ( .B(n2212), .A(n2213), .S(n2277), .Y(n2211) );
  MUX2X1 U1543 ( .B(n2215), .A(n2216), .S(n2295), .Y(n2214) );
  MUX2X1 U1544 ( .B(n2218), .A(n2219), .S(n2295), .Y(n2217) );
  MUX2X1 U1545 ( .B(n2221), .A(n2222), .S(n2295), .Y(n2220) );
  MUX2X1 U1546 ( .B(n2224), .A(n2225), .S(n2295), .Y(n2223) );
  MUX2X1 U1547 ( .B(n2227), .A(n2228), .S(n2277), .Y(n2226) );
  MUX2X1 U1548 ( .B(n2230), .A(n2231), .S(n2295), .Y(n2229) );
  MUX2X1 U1549 ( .B(n2233), .A(n2234), .S(n2295), .Y(n2232) );
  MUX2X1 U1550 ( .B(n2236), .A(n2237), .S(n2295), .Y(n2235) );
  MUX2X1 U1551 ( .B(n2239), .A(n2240), .S(n2295), .Y(n2238) );
  MUX2X1 U1552 ( .B(n2242), .A(n2243), .S(n2277), .Y(n2241) );
  MUX2X1 U1553 ( .B(n2245), .A(n2246), .S(n2295), .Y(n2244) );
  MUX2X1 U1554 ( .B(n2248), .A(n2249), .S(n2295), .Y(n2247) );
  MUX2X1 U1555 ( .B(n2251), .A(n2252), .S(n2295), .Y(n2250) );
  MUX2X1 U1556 ( .B(n2254), .A(n2255), .S(n2295), .Y(n2253) );
  MUX2X1 U1557 ( .B(n2257), .A(n2258), .S(n2277), .Y(n2256) );
  MUX2X1 U1558 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n2304), .Y(n1781) );
  MUX2X1 U1559 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n2304), .Y(n1780) );
  MUX2X1 U1560 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n2304), .Y(n1784) );
  MUX2X1 U1561 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n2304), .Y(n1783) );
  MUX2X1 U1562 ( .B(n1782), .A(n1779), .S(n2283), .Y(n1793) );
  MUX2X1 U1563 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n2305), .Y(n1787) );
  MUX2X1 U1564 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n2305), .Y(n1786) );
  MUX2X1 U1565 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n2305), .Y(n1790) );
  MUX2X1 U1566 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n2305), .Y(n1789) );
  MUX2X1 U1567 ( .B(n1788), .A(n1785), .S(n2283), .Y(n1792) );
  MUX2X1 U1568 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n2305), .Y(n1796) );
  MUX2X1 U1569 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n2305), .Y(n1795) );
  MUX2X1 U1570 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n2305), .Y(n1799) );
  MUX2X1 U1571 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n2305), .Y(n1798) );
  MUX2X1 U1572 ( .B(n1797), .A(n1794), .S(n2283), .Y(n1808) );
  MUX2X1 U1573 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n2305), .Y(n1802) );
  MUX2X1 U1574 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n2305), .Y(n1801) );
  MUX2X1 U1575 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n2305), .Y(n1805) );
  MUX2X1 U1576 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n2305), .Y(n1804) );
  MUX2X1 U1577 ( .B(n1803), .A(n1800), .S(n2283), .Y(n1807) );
  MUX2X1 U1578 ( .B(n1806), .A(n1791), .S(n2275), .Y(n2259) );
  MUX2X1 U1579 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n2306), .Y(n1811) );
  MUX2X1 U1580 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n2306), .Y(n1810) );
  MUX2X1 U1581 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n2306), .Y(n1814) );
  MUX2X1 U1582 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n2306), .Y(n1813) );
  MUX2X1 U1583 ( .B(n1812), .A(n1809), .S(n2283), .Y(n1823) );
  MUX2X1 U1584 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n2306), .Y(n1817) );
  MUX2X1 U1585 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n2306), .Y(n1816) );
  MUX2X1 U1586 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n2306), .Y(n1820) );
  MUX2X1 U1587 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n2306), .Y(n1819) );
  MUX2X1 U1588 ( .B(n1818), .A(n1815), .S(n2283), .Y(n1822) );
  MUX2X1 U1589 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n2306), .Y(n1826) );
  MUX2X1 U1590 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n2306), .Y(n1825) );
  MUX2X1 U1591 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n2306), .Y(n1829) );
  MUX2X1 U1592 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n2306), .Y(n1828) );
  MUX2X1 U1593 ( .B(n1827), .A(n1824), .S(n2283), .Y(n1838) );
  MUX2X1 U1594 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n2307), .Y(n1832) );
  MUX2X1 U1595 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n2307), .Y(n1831) );
  MUX2X1 U1596 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n2307), .Y(n1835) );
  MUX2X1 U1597 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n2307), .Y(n1834) );
  MUX2X1 U1598 ( .B(n1833), .A(n1830), .S(n2283), .Y(n1837) );
  MUX2X1 U1599 ( .B(n1836), .A(n1821), .S(n2275), .Y(n2260) );
  MUX2X1 U1600 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n2307), .Y(n1841) );
  MUX2X1 U1601 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n2307), .Y(n1840) );
  MUX2X1 U1602 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n2307), .Y(n1844) );
  MUX2X1 U1603 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n2307), .Y(n1843) );
  MUX2X1 U1604 ( .B(n1842), .A(n1839), .S(n2283), .Y(n1853) );
  MUX2X1 U1605 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n2307), .Y(n1847) );
  MUX2X1 U1606 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n2307), .Y(n1846) );
  MUX2X1 U1607 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n2307), .Y(n1850) );
  MUX2X1 U1608 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n2307), .Y(n1849) );
  MUX2X1 U1609 ( .B(n1848), .A(n1845), .S(n2283), .Y(n1852) );
  MUX2X1 U1610 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n2308), .Y(n1856) );
  MUX2X1 U1611 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n2308), .Y(n1855) );
  MUX2X1 U1612 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n2308), .Y(n1859) );
  MUX2X1 U1613 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n2308), .Y(n1858) );
  MUX2X1 U1614 ( .B(n1857), .A(n1854), .S(n2283), .Y(n1868) );
  MUX2X1 U1615 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n2308), .Y(n1862) );
  MUX2X1 U1616 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n2308), .Y(n1861) );
  MUX2X1 U1617 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n2308), .Y(n1865) );
  MUX2X1 U1618 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n2308), .Y(n1864) );
  MUX2X1 U1619 ( .B(n1863), .A(n1860), .S(n2283), .Y(n1867) );
  MUX2X1 U1620 ( .B(n1866), .A(n1851), .S(n2275), .Y(n2261) );
  MUX2X1 U1621 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n2308), .Y(n1871) );
  MUX2X1 U1622 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n2308), .Y(n1870) );
  MUX2X1 U1623 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n2308), .Y(n1874) );
  MUX2X1 U1624 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n2308), .Y(n1873) );
  MUX2X1 U1625 ( .B(n1872), .A(n1869), .S(n2282), .Y(n1883) );
  MUX2X1 U1626 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n2309), .Y(n1877) );
  MUX2X1 U1627 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n2309), .Y(n1876) );
  MUX2X1 U1628 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n2309), .Y(n1880) );
  MUX2X1 U1629 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n2309), .Y(n1879) );
  MUX2X1 U1630 ( .B(n1878), .A(n1875), .S(n2282), .Y(n1882) );
  MUX2X1 U1631 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n2309), .Y(n1886) );
  MUX2X1 U1632 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n2309), .Y(n1885) );
  MUX2X1 U1633 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n2309), .Y(n1889) );
  MUX2X1 U1634 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n2309), .Y(n1888) );
  MUX2X1 U1635 ( .B(n1887), .A(n1884), .S(n2282), .Y(n1898) );
  MUX2X1 U1636 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n2309), .Y(n1892) );
  MUX2X1 U1637 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n2309), .Y(n1891) );
  MUX2X1 U1638 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n2309), .Y(n1895) );
  MUX2X1 U1639 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n2309), .Y(n1894) );
  MUX2X1 U1640 ( .B(n1893), .A(n1890), .S(n2282), .Y(n1897) );
  MUX2X1 U1641 ( .B(n1896), .A(n1881), .S(n2275), .Y(n2262) );
  MUX2X1 U1642 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n2310), .Y(n1901) );
  MUX2X1 U1643 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n2310), .Y(n1900) );
  MUX2X1 U1644 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n2310), .Y(n1904) );
  MUX2X1 U1645 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n2310), .Y(n1903) );
  MUX2X1 U1646 ( .B(n1902), .A(n1899), .S(n2282), .Y(n1913) );
  MUX2X1 U1647 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n2310), .Y(n1907) );
  MUX2X1 U1648 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n2310), .Y(n1906) );
  MUX2X1 U1649 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n2310), .Y(n1910) );
  MUX2X1 U1650 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n2310), .Y(n1909) );
  MUX2X1 U1651 ( .B(n1908), .A(n1905), .S(n2282), .Y(n1912) );
  MUX2X1 U1652 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n2310), .Y(n1916) );
  MUX2X1 U1653 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n2310), .Y(n1915) );
  MUX2X1 U1654 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n2310), .Y(n1919) );
  MUX2X1 U1655 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n2310), .Y(n1918) );
  MUX2X1 U1656 ( .B(n1917), .A(n1914), .S(n2282), .Y(n1928) );
  MUX2X1 U1657 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n2311), .Y(n1922) );
  MUX2X1 U1658 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n2311), .Y(n1921) );
  MUX2X1 U1659 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n2311), .Y(n1925) );
  MUX2X1 U1660 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n2311), .Y(n1924) );
  MUX2X1 U1661 ( .B(n1923), .A(n1920), .S(n2282), .Y(n1927) );
  MUX2X1 U1662 ( .B(n1926), .A(n1911), .S(n2275), .Y(n2263) );
  MUX2X1 U1663 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n2311), .Y(n1931) );
  MUX2X1 U1664 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n2311), .Y(n1930) );
  MUX2X1 U1665 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n2311), .Y(n1934) );
  MUX2X1 U1666 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n2311), .Y(n1933) );
  MUX2X1 U1667 ( .B(n1932), .A(n1929), .S(n2282), .Y(n1943) );
  MUX2X1 U1668 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n2311), .Y(n1937) );
  MUX2X1 U1669 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n2311), .Y(n1936) );
  MUX2X1 U1670 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n2311), .Y(n1940) );
  MUX2X1 U1671 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n2311), .Y(n1939) );
  MUX2X1 U1672 ( .B(n1938), .A(n1935), .S(n2282), .Y(n1942) );
  MUX2X1 U1673 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n2312), .Y(n1946) );
  MUX2X1 U1674 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n2312), .Y(n1945) );
  MUX2X1 U1675 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n2312), .Y(n1949) );
  MUX2X1 U1676 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n2312), .Y(n1948) );
  MUX2X1 U1677 ( .B(n1947), .A(n1944), .S(n2282), .Y(n1958) );
  MUX2X1 U1678 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n2312), .Y(n1952) );
  MUX2X1 U1679 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n2312), .Y(n1951) );
  MUX2X1 U1680 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n2312), .Y(n1955) );
  MUX2X1 U1681 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n2312), .Y(n1954) );
  MUX2X1 U1682 ( .B(n1953), .A(n1950), .S(n2282), .Y(n1957) );
  MUX2X1 U1683 ( .B(n1956), .A(n1941), .S(n2275), .Y(n2264) );
  MUX2X1 U1684 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n2312), .Y(n1961) );
  MUX2X1 U1685 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n2312), .Y(n1960) );
  MUX2X1 U1686 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n2312), .Y(n1964) );
  MUX2X1 U1687 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n2312), .Y(n1963) );
  MUX2X1 U1688 ( .B(n1962), .A(n1959), .S(n2281), .Y(n1973) );
  MUX2X1 U1689 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n2313), .Y(n1967) );
  MUX2X1 U1690 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n2313), .Y(n1966) );
  MUX2X1 U1691 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n2313), .Y(n1970) );
  MUX2X1 U1692 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n2313), .Y(n1969) );
  MUX2X1 U1693 ( .B(n1968), .A(n1965), .S(n2281), .Y(n1972) );
  MUX2X1 U1694 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n2313), .Y(n1976) );
  MUX2X1 U1695 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n2313), .Y(n1975) );
  MUX2X1 U1696 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n2313), .Y(n1979) );
  MUX2X1 U1697 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n2313), .Y(n1978) );
  MUX2X1 U1698 ( .B(n1977), .A(n1974), .S(n2281), .Y(n1988) );
  MUX2X1 U1699 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n2313), .Y(n1982) );
  MUX2X1 U1700 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n2313), .Y(n1981) );
  MUX2X1 U1701 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n2313), .Y(n1985) );
  MUX2X1 U1702 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n2313), .Y(n1984) );
  MUX2X1 U1703 ( .B(n1983), .A(n1980), .S(n2281), .Y(n1987) );
  MUX2X1 U1704 ( .B(n1986), .A(n1971), .S(n2275), .Y(n2265) );
  MUX2X1 U1705 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n2314), .Y(n1991) );
  MUX2X1 U1706 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n2314), .Y(n1990) );
  MUX2X1 U1707 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n2314), .Y(n1994) );
  MUX2X1 U1708 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n2314), .Y(n1993) );
  MUX2X1 U1709 ( .B(n1992), .A(n1989), .S(n2281), .Y(n2003) );
  MUX2X1 U1710 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n2314), .Y(n1997) );
  MUX2X1 U1711 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n2314), .Y(n1996) );
  MUX2X1 U1712 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n2314), .Y(n2000) );
  MUX2X1 U1713 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n2314), .Y(n1999) );
  MUX2X1 U1714 ( .B(n1998), .A(n1995), .S(n2281), .Y(n2002) );
  MUX2X1 U1715 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n2314), .Y(n2006) );
  MUX2X1 U1716 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n2314), .Y(n2005) );
  MUX2X1 U1717 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n2314), .Y(n2009) );
  MUX2X1 U1718 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n2314), .Y(n2008) );
  MUX2X1 U1719 ( .B(n2007), .A(n2004), .S(n2281), .Y(n2018) );
  MUX2X1 U1720 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n2315), .Y(n2012) );
  MUX2X1 U1721 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n2315), .Y(n2011) );
  MUX2X1 U1722 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n2315), .Y(n2015) );
  MUX2X1 U1723 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n2315), .Y(n2014) );
  MUX2X1 U1724 ( .B(n2013), .A(n2010), .S(n2281), .Y(n2017) );
  MUX2X1 U1725 ( .B(n2016), .A(n2001), .S(n2275), .Y(n2266) );
  MUX2X1 U1726 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n2315), .Y(n2021) );
  MUX2X1 U1727 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n2315), .Y(n2020) );
  MUX2X1 U1728 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n2315), .Y(n2024) );
  MUX2X1 U1729 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n2315), .Y(n2023) );
  MUX2X1 U1730 ( .B(n2022), .A(n2019), .S(n2281), .Y(n2033) );
  MUX2X1 U1731 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n2315), .Y(n2027) );
  MUX2X1 U1732 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n2315), .Y(n2026) );
  MUX2X1 U1733 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n2315), .Y(n2030) );
  MUX2X1 U1734 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n2315), .Y(n2029) );
  MUX2X1 U1735 ( .B(n2028), .A(n2025), .S(n2281), .Y(n2032) );
  MUX2X1 U1736 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n2316), .Y(n2036) );
  MUX2X1 U1737 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n2316), .Y(n2035) );
  MUX2X1 U1738 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n2316), .Y(n2039) );
  MUX2X1 U1739 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n2316), .Y(n2038) );
  MUX2X1 U1740 ( .B(n2037), .A(n2034), .S(n2281), .Y(n2048) );
  MUX2X1 U1741 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n2316), .Y(n2042) );
  MUX2X1 U1742 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n2316), .Y(n2041) );
  MUX2X1 U1743 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n2316), .Y(n2045) );
  MUX2X1 U1744 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n2316), .Y(n2044) );
  MUX2X1 U1745 ( .B(n2043), .A(n2040), .S(n2281), .Y(n2047) );
  MUX2X1 U1746 ( .B(n2046), .A(n2031), .S(n2275), .Y(n2267) );
  MUX2X1 U1747 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n2316), .Y(n2051) );
  MUX2X1 U1748 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n2316), .Y(n2050) );
  MUX2X1 U1749 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n2316), .Y(n2054) );
  MUX2X1 U1750 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n2316), .Y(n2053) );
  MUX2X1 U1751 ( .B(n2052), .A(n2049), .S(n2280), .Y(n2063) );
  MUX2X1 U1752 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n2317), .Y(n2057) );
  MUX2X1 U1753 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n2317), .Y(n2056) );
  MUX2X1 U1754 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n2317), .Y(n2060) );
  MUX2X1 U1755 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n2317), .Y(n2059) );
  MUX2X1 U1756 ( .B(n2058), .A(n2055), .S(n2280), .Y(n2062) );
  MUX2X1 U1757 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n2317), .Y(n2066) );
  MUX2X1 U1758 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n2317), .Y(n2065) );
  MUX2X1 U1759 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n2317), .Y(n2069) );
  MUX2X1 U1760 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n2317), .Y(n2068) );
  MUX2X1 U1761 ( .B(n2067), .A(n2064), .S(n2280), .Y(n2078) );
  MUX2X1 U1762 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n2317), .Y(n2072) );
  MUX2X1 U1763 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n2317), .Y(n2071) );
  MUX2X1 U1764 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n2317), .Y(n2075) );
  MUX2X1 U1765 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n2317), .Y(n2074) );
  MUX2X1 U1766 ( .B(n2073), .A(n2070), .S(n2280), .Y(n2077) );
  MUX2X1 U1767 ( .B(n2076), .A(n2061), .S(n2275), .Y(n2268) );
  MUX2X1 U1768 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n2318), .Y(n2081) );
  MUX2X1 U1769 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n2318), .Y(n2080) );
  MUX2X1 U1770 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n2318), .Y(n2084) );
  MUX2X1 U1771 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n2318), .Y(n2083) );
  MUX2X1 U1772 ( .B(n2082), .A(n2079), .S(n2280), .Y(n2093) );
  MUX2X1 U1773 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n2318), .Y(n2087) );
  MUX2X1 U1774 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n2318), .Y(n2086) );
  MUX2X1 U1775 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n2318), .Y(n2090) );
  MUX2X1 U1776 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n2318), .Y(n2089) );
  MUX2X1 U1777 ( .B(n2088), .A(n2085), .S(n2280), .Y(n2092) );
  MUX2X1 U1778 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n2318), .Y(n2096) );
  MUX2X1 U1779 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n2318), .Y(n2095) );
  MUX2X1 U1780 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n2318), .Y(n2099) );
  MUX2X1 U1781 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n2318), .Y(n2098) );
  MUX2X1 U1782 ( .B(n2097), .A(n2094), .S(n2280), .Y(n2108) );
  MUX2X1 U1783 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n2319), .Y(n2102) );
  MUX2X1 U1784 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n2319), .Y(n2101) );
  MUX2X1 U1785 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n2319), .Y(n2105) );
  MUX2X1 U1786 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n2319), .Y(n2104) );
  MUX2X1 U1787 ( .B(n2103), .A(n2100), .S(n2280), .Y(n2107) );
  MUX2X1 U1788 ( .B(n2106), .A(n2091), .S(n2275), .Y(n2269) );
  MUX2X1 U1789 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n2319), .Y(n2111) );
  MUX2X1 U1790 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n2319), .Y(n2110) );
  MUX2X1 U1791 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n2319), .Y(n2114) );
  MUX2X1 U1792 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n2319), .Y(n2113) );
  MUX2X1 U1793 ( .B(n2112), .A(n2109), .S(n2280), .Y(n2123) );
  MUX2X1 U1794 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n2319), .Y(n2117) );
  MUX2X1 U1795 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n2319), .Y(n2116) );
  MUX2X1 U1796 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n2319), .Y(n2120) );
  MUX2X1 U1797 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n2319), .Y(n2119) );
  MUX2X1 U1798 ( .B(n2118), .A(n2115), .S(n2280), .Y(n2122) );
  MUX2X1 U1799 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n2320), .Y(n2126) );
  MUX2X1 U1800 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n2320), .Y(n2125) );
  MUX2X1 U1801 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n2320), .Y(n2129) );
  MUX2X1 U1802 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n2320), .Y(n2128) );
  MUX2X1 U1803 ( .B(n2127), .A(n2124), .S(n2280), .Y(n2138) );
  MUX2X1 U1804 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n2320), .Y(n2132) );
  MUX2X1 U1805 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n2320), .Y(n2131) );
  MUX2X1 U1806 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n2320), .Y(n2135) );
  MUX2X1 U1807 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n2320), .Y(n2134) );
  MUX2X1 U1808 ( .B(n2133), .A(n2130), .S(n2280), .Y(n2137) );
  MUX2X1 U1809 ( .B(n2136), .A(n2121), .S(n2275), .Y(n2270) );
  MUX2X1 U1810 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n2320), .Y(n2141) );
  MUX2X1 U1811 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n2320), .Y(n2140) );
  MUX2X1 U1812 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n2320), .Y(n2144) );
  MUX2X1 U1813 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n2320), .Y(n2143) );
  MUX2X1 U1814 ( .B(n2142), .A(n2139), .S(n2279), .Y(n2153) );
  MUX2X1 U1815 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n2321), .Y(n2147) );
  MUX2X1 U1816 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n2321), .Y(n2146) );
  MUX2X1 U1817 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n2321), .Y(n2150) );
  MUX2X1 U1818 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n2321), .Y(n2149) );
  MUX2X1 U1819 ( .B(n2148), .A(n2145), .S(n2279), .Y(n2152) );
  MUX2X1 U1820 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n2321), .Y(n2156) );
  MUX2X1 U1821 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n2321), .Y(n2155) );
  MUX2X1 U1822 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n2321), .Y(n2159) );
  MUX2X1 U1823 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n2321), .Y(n2158) );
  MUX2X1 U1824 ( .B(n2157), .A(n2154), .S(n2279), .Y(n2168) );
  MUX2X1 U1825 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n2321), .Y(n2162) );
  MUX2X1 U1826 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n2321), .Y(n2161) );
  MUX2X1 U1827 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n2321), .Y(n2165) );
  MUX2X1 U1828 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n2321), .Y(n2164) );
  MUX2X1 U1829 ( .B(n2163), .A(n2160), .S(n2279), .Y(n2167) );
  MUX2X1 U1830 ( .B(n2166), .A(n2151), .S(n2275), .Y(n2271) );
  MUX2X1 U1831 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n2322), .Y(n2171) );
  MUX2X1 U1832 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n2322), .Y(n2170) );
  MUX2X1 U1833 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n2322), .Y(n2174) );
  MUX2X1 U1834 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n2322), .Y(n2173) );
  MUX2X1 U1835 ( .B(n2172), .A(n2169), .S(n2279), .Y(n2183) );
  MUX2X1 U1836 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n2322), .Y(n2177) );
  MUX2X1 U1837 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n2322), .Y(n2176) );
  MUX2X1 U1838 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n2322), .Y(n2180) );
  MUX2X1 U1839 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n2322), .Y(n2179) );
  MUX2X1 U1840 ( .B(n2178), .A(n2175), .S(n2279), .Y(n2182) );
  MUX2X1 U1841 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n2322), .Y(n2186) );
  MUX2X1 U1842 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n2322), .Y(n2185) );
  MUX2X1 U1843 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n2322), .Y(n2189) );
  MUX2X1 U1844 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n2322), .Y(n2188) );
  MUX2X1 U1845 ( .B(n2187), .A(n2184), .S(n2279), .Y(n2198) );
  MUX2X1 U1846 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n2323), .Y(n2192) );
  MUX2X1 U1847 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n2323), .Y(n2191) );
  MUX2X1 U1848 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n2323), .Y(n2195) );
  MUX2X1 U1849 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n2323), .Y(n2194) );
  MUX2X1 U1850 ( .B(n2193), .A(n2190), .S(n2279), .Y(n2197) );
  MUX2X1 U1851 ( .B(n2196), .A(n2181), .S(n2275), .Y(n2272) );
  MUX2X1 U1852 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n2323), .Y(n2201) );
  MUX2X1 U1853 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n2323), .Y(n2200) );
  MUX2X1 U1854 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n2323), .Y(n2204) );
  MUX2X1 U1855 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n2323), .Y(n2203) );
  MUX2X1 U1856 ( .B(n2202), .A(n2199), .S(n2279), .Y(n2213) );
  MUX2X1 U1857 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n2323), .Y(n2207) );
  MUX2X1 U1858 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n2323), .Y(n2206) );
  MUX2X1 U1859 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n2323), .Y(n2210) );
  MUX2X1 U1860 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n2323), .Y(n2209) );
  MUX2X1 U1861 ( .B(n2208), .A(n2205), .S(n2279), .Y(n2212) );
  MUX2X1 U1862 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n2324), .Y(n2216) );
  MUX2X1 U1863 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n2324), .Y(n2215) );
  MUX2X1 U1864 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n2324), .Y(n2219) );
  MUX2X1 U1865 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n2324), .Y(n2218) );
  MUX2X1 U1866 ( .B(n2217), .A(n2214), .S(n2279), .Y(n2228) );
  MUX2X1 U1867 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n2324), .Y(n2222) );
  MUX2X1 U1868 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n2324), .Y(n2221) );
  MUX2X1 U1869 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n2324), .Y(n2225) );
  MUX2X1 U1870 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n2324), .Y(n2224) );
  MUX2X1 U1871 ( .B(n2223), .A(n2220), .S(n2279), .Y(n2227) );
  MUX2X1 U1872 ( .B(n2226), .A(n2211), .S(n2275), .Y(n2273) );
  MUX2X1 U1873 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n2324), .Y(n2231) );
  MUX2X1 U1874 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n2324), .Y(n2230) );
  MUX2X1 U1875 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n2324), .Y(n2234) );
  MUX2X1 U1876 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n2324), .Y(n2233) );
  MUX2X1 U1877 ( .B(n2232), .A(n2229), .S(n2280), .Y(n2243) );
  MUX2X1 U1878 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n2325), .Y(n2237) );
  MUX2X1 U1879 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n2325), .Y(n2236) );
  MUX2X1 U1880 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n2325), .Y(n2240) );
  MUX2X1 U1881 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n2325), .Y(n2239) );
  MUX2X1 U1882 ( .B(n2238), .A(n2235), .S(n2279), .Y(n2242) );
  MUX2X1 U1883 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n2325), .Y(n2246) );
  MUX2X1 U1884 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n2325), .Y(n2245) );
  MUX2X1 U1885 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n2325), .Y(n2249) );
  MUX2X1 U1886 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n2325), .Y(n2248) );
  MUX2X1 U1887 ( .B(n2247), .A(n2244), .S(n2279), .Y(n2258) );
  MUX2X1 U1888 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n2325), .Y(n2252) );
  MUX2X1 U1889 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n2325), .Y(n2251) );
  MUX2X1 U1890 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n2325), .Y(n2255) );
  MUX2X1 U1891 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n2325), .Y(n2254) );
  MUX2X1 U1892 ( .B(n2253), .A(n2250), .S(n2279), .Y(n2257) );
  MUX2X1 U1893 ( .B(n2256), .A(n2241), .S(n2275), .Y(n2274) );
  INVX8 U1894 ( .A(n2296), .Y(n2284) );
  INVX8 U1895 ( .A(n2328), .Y(n2298) );
  INVX8 U1896 ( .A(n2327), .Y(n2299) );
  INVX8 U1897 ( .A(n2327), .Y(n2300) );
  INVX8 U1898 ( .A(n2328), .Y(n2301) );
  INVX8 U1899 ( .A(n2328), .Y(n2302) );
  INVX8 U1900 ( .A(n2328), .Y(n2303) );
  INVX8 U1901 ( .A(n2303), .Y(n2304) );
  INVX8 U1902 ( .A(n2303), .Y(n2305) );
  INVX8 U1903 ( .A(n2303), .Y(n2306) );
  INVX8 U1904 ( .A(n2302), .Y(n2307) );
  INVX8 U1905 ( .A(n2302), .Y(n2308) );
  INVX8 U1906 ( .A(n2302), .Y(n2309) );
  INVX8 U1907 ( .A(n2301), .Y(n2310) );
  INVX8 U1908 ( .A(n2301), .Y(n2311) );
  INVX8 U1909 ( .A(n2301), .Y(n2312) );
  INVX8 U1910 ( .A(n2300), .Y(n2313) );
  INVX8 U1911 ( .A(n2300), .Y(n2314) );
  INVX8 U1912 ( .A(n2300), .Y(n2315) );
  INVX8 U1913 ( .A(n2326), .Y(n2316) );
  INVX8 U1914 ( .A(n2297), .Y(n2317) );
  INVX8 U1915 ( .A(n2301), .Y(n2318) );
  INVX8 U1916 ( .A(n2299), .Y(n2319) );
  INVX8 U1917 ( .A(n2299), .Y(n2320) );
  INVX8 U1918 ( .A(n2299), .Y(n2321) );
  INVX8 U1919 ( .A(n2298), .Y(n2322) );
  INVX8 U1920 ( .A(n2298), .Y(n2323) );
  INVX8 U1921 ( .A(n2298), .Y(n2324) );
  INVX8 U1922 ( .A(n2297), .Y(n2325) );
  INVX8 U1923 ( .A(n2326), .Y(n2327) );
  INVX8 U1924 ( .A(n2326), .Y(n2328) );
  INVX8 U1925 ( .A(n2431), .Y(n2461) );
  INVX1 U1926 ( .A(N10), .Y(n2423) );
  INVX8 U1927 ( .A(n92), .Y(n2389) );
  INVX8 U1928 ( .A(n92), .Y(n2390) );
  INVX8 U1929 ( .A(n93), .Y(n2391) );
  INVX8 U1930 ( .A(n93), .Y(n2392) );
  INVX8 U1931 ( .A(n94), .Y(n2393) );
  INVX8 U1932 ( .A(n94), .Y(n2394) );
  INVX8 U1933 ( .A(n95), .Y(n2395) );
  INVX8 U1934 ( .A(n95), .Y(n2396) );
  INVX8 U1935 ( .A(n96), .Y(n2397) );
  INVX8 U1936 ( .A(n96), .Y(n2398) );
  INVX8 U1937 ( .A(n97), .Y(n2399) );
  INVX8 U1938 ( .A(n97), .Y(n2400) );
  INVX8 U1939 ( .A(n98), .Y(n2401) );
  INVX8 U1940 ( .A(n98), .Y(n2402) );
  INVX8 U1941 ( .A(n99), .Y(n2403) );
  INVX8 U1942 ( .A(n99), .Y(n2404) );
  INVX8 U1943 ( .A(n100), .Y(n2405) );
  INVX8 U1944 ( .A(n100), .Y(n2406) );
  INVX8 U1945 ( .A(n101), .Y(n2407) );
  INVX8 U1946 ( .A(n101), .Y(n2408) );
  INVX8 U1947 ( .A(n102), .Y(n2409) );
  INVX8 U1948 ( .A(n102), .Y(n2410) );
  INVX8 U1949 ( .A(n103), .Y(n2411) );
  INVX8 U1950 ( .A(n103), .Y(n2412) );
  INVX8 U1951 ( .A(n104), .Y(n2413) );
  INVX8 U1952 ( .A(n104), .Y(n2414) );
  INVX8 U1953 ( .A(n105), .Y(n2415) );
  INVX8 U1954 ( .A(n105), .Y(n2416) );
  INVX8 U1955 ( .A(n106), .Y(n2417) );
  INVX8 U1956 ( .A(n106), .Y(n2418) );
  INVX8 U1957 ( .A(n107), .Y(n2419) );
  INVX8 U1958 ( .A(n107), .Y(n2420) );
  OAI21X1 U1959 ( .A(n2330), .B(n2389), .C(n138), .Y(n2973) );
  OAI21X1 U1960 ( .A(n2391), .B(n2329), .C(n1422), .Y(n2972) );
  OAI21X1 U1961 ( .A(n2393), .B(n2329), .C(n1424), .Y(n2971) );
  OAI21X1 U1962 ( .A(n2395), .B(n2329), .C(n1426), .Y(n2970) );
  OAI21X1 U1963 ( .A(n2397), .B(n2329), .C(n1428), .Y(n2969) );
  OAI21X1 U1964 ( .A(n2399), .B(n2329), .C(n1430), .Y(n2968) );
  OAI21X1 U1965 ( .A(n2401), .B(n2329), .C(n1432), .Y(n2967) );
  OAI21X1 U1966 ( .A(n2403), .B(n2329), .C(n1434), .Y(n2966) );
  OAI21X1 U1967 ( .A(n2406), .B(n2329), .C(n1436), .Y(n2965) );
  OAI21X1 U1968 ( .A(n2408), .B(n2330), .C(n1438), .Y(n2964) );
  OAI21X1 U1969 ( .A(n2410), .B(n2330), .C(n1440), .Y(n2963) );
  OAI21X1 U1970 ( .A(n2412), .B(n2330), .C(n1442), .Y(n2962) );
  OAI21X1 U1971 ( .A(n2414), .B(n2330), .C(n1444), .Y(n2961) );
  OAI21X1 U1972 ( .A(n2416), .B(n2330), .C(n1446), .Y(n2960) );
  OAI21X1 U1973 ( .A(n2418), .B(n2330), .C(n1448), .Y(n2959) );
  OAI21X1 U1974 ( .A(n2420), .B(n2330), .C(n1450), .Y(n2958) );
  OAI21X1 U1975 ( .A(n2331), .B(n2389), .C(n140), .Y(n2957) );
  OAI21X1 U1976 ( .A(n2331), .B(n2392), .C(n1452), .Y(n2956) );
  OAI21X1 U1977 ( .A(n2331), .B(n2394), .C(n1454), .Y(n2955) );
  OAI21X1 U1978 ( .A(n2331), .B(n2396), .C(n1456), .Y(n2954) );
  OAI21X1 U1979 ( .A(n2331), .B(n2398), .C(n1458), .Y(n2953) );
  OAI21X1 U1980 ( .A(n2331), .B(n2400), .C(n1460), .Y(n2952) );
  OAI21X1 U1981 ( .A(n2331), .B(n2402), .C(n1462), .Y(n2951) );
  OAI21X1 U1982 ( .A(n2331), .B(n2404), .C(n1464), .Y(n2950) );
  OAI21X1 U1983 ( .A(n2332), .B(n2405), .C(n1466), .Y(n2949) );
  OAI21X1 U1984 ( .A(n2332), .B(n2407), .C(n1468), .Y(n2948) );
  OAI21X1 U1985 ( .A(n2332), .B(n2409), .C(n1470), .Y(n2947) );
  OAI21X1 U1986 ( .A(n2332), .B(n2411), .C(n1472), .Y(n2946) );
  OAI21X1 U1987 ( .A(n2332), .B(n2413), .C(n1474), .Y(n2945) );
  OAI21X1 U1988 ( .A(n2332), .B(n2415), .C(n1476), .Y(n2944) );
  OAI21X1 U1989 ( .A(n2332), .B(n2417), .C(n1478), .Y(n2943) );
  OAI21X1 U1990 ( .A(n2332), .B(n2419), .C(n1480), .Y(n2942) );
  NAND3X1 U1991 ( .A(n2422), .B(n2425), .C(n2424), .Y(n2434) );
  OAI21X1 U1992 ( .A(n2333), .B(n2389), .C(n142), .Y(n2941) );
  OAI21X1 U1993 ( .A(n2333), .B(n2392), .C(n1482), .Y(n2940) );
  OAI21X1 U1994 ( .A(n2394), .B(n2333), .C(n1484), .Y(n2939) );
  OAI21X1 U1995 ( .A(n2333), .B(n2396), .C(n1486), .Y(n2938) );
  OAI21X1 U1996 ( .A(n2333), .B(n2398), .C(n1488), .Y(n2937) );
  OAI21X1 U1997 ( .A(n2333), .B(n2400), .C(n1490), .Y(n2936) );
  OAI21X1 U1998 ( .A(n2333), .B(n2402), .C(n1492), .Y(n2935) );
  OAI21X1 U1999 ( .A(n2333), .B(n2404), .C(n1494), .Y(n2934) );
  OAI21X1 U2000 ( .A(n2334), .B(n2406), .C(n1496), .Y(n2933) );
  OAI21X1 U2001 ( .A(n2334), .B(n2408), .C(n1498), .Y(n2932) );
  OAI21X1 U2002 ( .A(n2334), .B(n2410), .C(n1500), .Y(n2931) );
  OAI21X1 U2003 ( .A(n2334), .B(n2412), .C(n1502), .Y(n2930) );
  OAI21X1 U2004 ( .A(n2334), .B(n2414), .C(n1504), .Y(n2929) );
  OAI21X1 U2005 ( .A(n2334), .B(n2416), .C(n1506), .Y(n2928) );
  OAI21X1 U2006 ( .A(n2334), .B(n2418), .C(n1508), .Y(n2927) );
  OAI21X1 U2007 ( .A(n2334), .B(n2420), .C(n1510), .Y(n2926) );
  NAND3X1 U2008 ( .A(n2425), .B(n2424), .C(n2423), .Y(n2436) );
  OAI21X1 U2009 ( .A(n2335), .B(n2389), .C(n144), .Y(n2925) );
  OAI21X1 U2010 ( .A(n2335), .B(n2391), .C(n1512), .Y(n2924) );
  OAI21X1 U2011 ( .A(n2335), .B(n2393), .C(n1514), .Y(n2923) );
  OAI21X1 U2012 ( .A(n2335), .B(n2395), .C(n1516), .Y(n2922) );
  OAI21X1 U2013 ( .A(n2335), .B(n2397), .C(n1518), .Y(n2921) );
  OAI21X1 U2014 ( .A(n2335), .B(n2399), .C(n1520), .Y(n2920) );
  OAI21X1 U2015 ( .A(n2335), .B(n2401), .C(n1522), .Y(n2919) );
  OAI21X1 U2016 ( .A(n2335), .B(n2403), .C(n1524), .Y(n2918) );
  OAI21X1 U2017 ( .A(n2336), .B(n2405), .C(n1526), .Y(n2917) );
  OAI21X1 U2018 ( .A(n2336), .B(n2407), .C(n1528), .Y(n2916) );
  OAI21X1 U2019 ( .A(n2336), .B(n2409), .C(n1530), .Y(n2915) );
  OAI21X1 U2020 ( .A(n2336), .B(n2411), .C(n1532), .Y(n2914) );
  OAI21X1 U2021 ( .A(n2336), .B(n2413), .C(n1534), .Y(n2913) );
  OAI21X1 U2022 ( .A(n2336), .B(n2415), .C(n1536), .Y(n2912) );
  OAI21X1 U2023 ( .A(n2336), .B(n2417), .C(n1538), .Y(n2911) );
  OAI21X1 U2024 ( .A(n2336), .B(n2419), .C(n1540), .Y(n2910) );
  NAND3X1 U2025 ( .A(n2422), .B(n2292), .C(n2426), .Y(n2438) );
  OAI21X1 U2026 ( .A(n2337), .B(n2389), .C(n146), .Y(n2909) );
  OAI21X1 U2027 ( .A(n2337), .B(n2392), .C(n1542), .Y(n2908) );
  OAI21X1 U2028 ( .A(n2337), .B(n2394), .C(n1544), .Y(n2907) );
  OAI21X1 U2029 ( .A(n2337), .B(n2396), .C(n1546), .Y(n2906) );
  OAI21X1 U2030 ( .A(n2337), .B(n2398), .C(n1548), .Y(n2905) );
  OAI21X1 U2031 ( .A(n2337), .B(n2400), .C(n1550), .Y(n2904) );
  OAI21X1 U2032 ( .A(n2337), .B(n2402), .C(n1552), .Y(n2903) );
  OAI21X1 U2033 ( .A(n2337), .B(n2404), .C(n1554), .Y(n2902) );
  OAI21X1 U2034 ( .A(n2338), .B(n2406), .C(n1556), .Y(n2901) );
  OAI21X1 U2035 ( .A(n2338), .B(n2408), .C(n1558), .Y(n2900) );
  OAI21X1 U2036 ( .A(n2338), .B(n2410), .C(n1560), .Y(n2899) );
  OAI21X1 U2037 ( .A(n2338), .B(n2412), .C(n1562), .Y(n2898) );
  OAI21X1 U2038 ( .A(n2338), .B(n2414), .C(n1564), .Y(n2897) );
  OAI21X1 U2039 ( .A(n2338), .B(n2416), .C(n1566), .Y(n2896) );
  OAI21X1 U2040 ( .A(n2338), .B(n2418), .C(n1568), .Y(n2895) );
  OAI21X1 U2041 ( .A(n2338), .B(n2420), .C(n1570), .Y(n2894) );
  NAND3X1 U2042 ( .A(n2426), .B(n2292), .C(n2423), .Y(n2440) );
  OAI21X1 U2043 ( .A(n2339), .B(n2389), .C(n148), .Y(n2893) );
  OAI21X1 U2044 ( .A(n2339), .B(n2391), .C(n1572), .Y(n2892) );
  OAI21X1 U2045 ( .A(n2339), .B(n2394), .C(n1574), .Y(n2891) );
  OAI21X1 U2046 ( .A(n2339), .B(n2395), .C(n1576), .Y(n2890) );
  OAI21X1 U2047 ( .A(n2339), .B(n2397), .C(n1578), .Y(n2889) );
  OAI21X1 U2048 ( .A(n2339), .B(n2399), .C(n1580), .Y(n2888) );
  OAI21X1 U2049 ( .A(n2339), .B(n2401), .C(n1582), .Y(n2887) );
  OAI21X1 U2050 ( .A(n2339), .B(n2403), .C(n1584), .Y(n2886) );
  OAI21X1 U2051 ( .A(n2340), .B(n2405), .C(n1586), .Y(n2885) );
  OAI21X1 U2052 ( .A(n2340), .B(n2407), .C(n1588), .Y(n2884) );
  OAI21X1 U2053 ( .A(n2340), .B(n2409), .C(n1590), .Y(n2883) );
  OAI21X1 U2054 ( .A(n2340), .B(n2411), .C(n1592), .Y(n2882) );
  OAI21X1 U2055 ( .A(n2340), .B(n2413), .C(n1594), .Y(n2881) );
  OAI21X1 U2056 ( .A(n2340), .B(n2415), .C(n1596), .Y(n2880) );
  OAI21X1 U2057 ( .A(n2340), .B(n2417), .C(n1598), .Y(n2879) );
  OAI21X1 U2058 ( .A(n2340), .B(n2419), .C(n1600), .Y(n2878) );
  NAND3X1 U2059 ( .A(n2422), .B(n2426), .C(n2424), .Y(n2442) );
  OAI21X1 U2060 ( .A(n2341), .B(n2389), .C(n150), .Y(n2877) );
  OAI21X1 U2061 ( .A(n2341), .B(n2392), .C(n1602), .Y(n2876) );
  OAI21X1 U2062 ( .A(n2341), .B(n2394), .C(n1604), .Y(n2875) );
  OAI21X1 U2063 ( .A(n2341), .B(n2396), .C(n1606), .Y(n2874) );
  OAI21X1 U2064 ( .A(n2341), .B(n2398), .C(n1608), .Y(n2873) );
  OAI21X1 U2065 ( .A(n2341), .B(n2400), .C(n1610), .Y(n2872) );
  OAI21X1 U2066 ( .A(n2341), .B(n2402), .C(n1612), .Y(n2871) );
  OAI21X1 U2067 ( .A(n2341), .B(n2404), .C(n1614), .Y(n2870) );
  OAI21X1 U2068 ( .A(n2342), .B(n2406), .C(n1616), .Y(n2869) );
  OAI21X1 U2069 ( .A(n2342), .B(n2408), .C(n1618), .Y(n2868) );
  OAI21X1 U2070 ( .A(n2342), .B(n2410), .C(n1620), .Y(n2867) );
  OAI21X1 U2071 ( .A(n2342), .B(n2412), .C(n1622), .Y(n2866) );
  OAI21X1 U2072 ( .A(n2342), .B(n2414), .C(n1624), .Y(n2865) );
  OAI21X1 U2073 ( .A(n2342), .B(n2416), .C(n1626), .Y(n2864) );
  OAI21X1 U2074 ( .A(n2342), .B(n2418), .C(n1628), .Y(n2863) );
  OAI21X1 U2075 ( .A(n2342), .B(n2420), .C(n1630), .Y(n2862) );
  NOR3X1 U2076 ( .A(n2422), .B(n2292), .C(n2425), .Y(n2460) );
  OAI21X1 U2077 ( .A(n2343), .B(n2389), .C(n152), .Y(n2861) );
  OAI21X1 U2078 ( .A(n2343), .B(n2391), .C(n1632), .Y(n2860) );
  OAI21X1 U2079 ( .A(n2343), .B(n2394), .C(n1634), .Y(n2859) );
  OAI21X1 U2080 ( .A(n2343), .B(n2395), .C(n1636), .Y(n2858) );
  OAI21X1 U2081 ( .A(n2343), .B(n2397), .C(n1638), .Y(n2857) );
  OAI21X1 U2082 ( .A(n2343), .B(n2399), .C(n1640), .Y(n2856) );
  OAI21X1 U2083 ( .A(n2343), .B(n2401), .C(n1642), .Y(n2855) );
  OAI21X1 U2084 ( .A(n2343), .B(n2403), .C(n1644), .Y(n2854) );
  OAI21X1 U2085 ( .A(n2343), .B(n2405), .C(n1646), .Y(n2853) );
  OAI21X1 U2086 ( .A(n2343), .B(n2407), .C(n1648), .Y(n2852) );
  OAI21X1 U2087 ( .A(n2343), .B(n2409), .C(n1650), .Y(n2851) );
  OAI21X1 U2088 ( .A(n2343), .B(n2411), .C(n1652), .Y(n2850) );
  OAI21X1 U2089 ( .A(n2343), .B(n2413), .C(n1654), .Y(n2849) );
  OAI21X1 U2090 ( .A(n2343), .B(n2415), .C(n1656), .Y(n2848) );
  OAI21X1 U2091 ( .A(n2343), .B(n2417), .C(n1658), .Y(n2847) );
  OAI21X1 U2092 ( .A(n2343), .B(n2419), .C(n1660), .Y(n2846) );
  OAI21X1 U2093 ( .A(n2344), .B(n2389), .C(n154), .Y(n2845) );
  OAI21X1 U2094 ( .A(n2344), .B(n2392), .C(n156), .Y(n2844) );
  OAI21X1 U2095 ( .A(n2344), .B(n2394), .C(n158), .Y(n2843) );
  OAI21X1 U2096 ( .A(n2344), .B(n2396), .C(n160), .Y(n2842) );
  OAI21X1 U2097 ( .A(n2344), .B(n2398), .C(n162), .Y(n2841) );
  OAI21X1 U2098 ( .A(n2344), .B(n2400), .C(n164), .Y(n2840) );
  OAI21X1 U2099 ( .A(n2344), .B(n2402), .C(n166), .Y(n2839) );
  OAI21X1 U2100 ( .A(n2344), .B(n2404), .C(n168), .Y(n2838) );
  OAI21X1 U2101 ( .A(n2345), .B(n2406), .C(n170), .Y(n2837) );
  OAI21X1 U2102 ( .A(n2345), .B(n2408), .C(n172), .Y(n2836) );
  OAI21X1 U2103 ( .A(n2345), .B(n2410), .C(n174), .Y(n2835) );
  OAI21X1 U2104 ( .A(n2345), .B(n2412), .C(n176), .Y(n2834) );
  OAI21X1 U2105 ( .A(n2345), .B(n2414), .C(n178), .Y(n2833) );
  OAI21X1 U2106 ( .A(n2345), .B(n2416), .C(n180), .Y(n2832) );
  OAI21X1 U2107 ( .A(n2345), .B(n2418), .C(n182), .Y(n2831) );
  OAI21X1 U2108 ( .A(n2345), .B(n2420), .C(n184), .Y(n2830) );
  OAI21X1 U2109 ( .A(n2346), .B(n2389), .C(n186), .Y(n2829) );
  OAI21X1 U2110 ( .A(n2346), .B(n2392), .C(n188), .Y(n2828) );
  OAI21X1 U2111 ( .A(n2346), .B(n2394), .C(n190), .Y(n2827) );
  OAI21X1 U2112 ( .A(n2346), .B(n2396), .C(n192), .Y(n2826) );
  OAI21X1 U2113 ( .A(n2346), .B(n2398), .C(n194), .Y(n2825) );
  OAI21X1 U2114 ( .A(n2346), .B(n2400), .C(n196), .Y(n2824) );
  OAI21X1 U2115 ( .A(n2346), .B(n2402), .C(n198), .Y(n2823) );
  OAI21X1 U2116 ( .A(n2346), .B(n2404), .C(n200), .Y(n2822) );
  OAI21X1 U2117 ( .A(n2347), .B(n2406), .C(n202), .Y(n2821) );
  OAI21X1 U2118 ( .A(n2347), .B(n2408), .C(n204), .Y(n2820) );
  OAI21X1 U2119 ( .A(n2347), .B(n2410), .C(n206), .Y(n2819) );
  OAI21X1 U2120 ( .A(n2347), .B(n2412), .C(n208), .Y(n2818) );
  OAI21X1 U2121 ( .A(n2347), .B(n2414), .C(n210), .Y(n2817) );
  OAI21X1 U2122 ( .A(n2347), .B(n2416), .C(n212), .Y(n2816) );
  OAI21X1 U2123 ( .A(n2347), .B(n2418), .C(n215), .Y(n2815) );
  OAI21X1 U2124 ( .A(n2347), .B(n2420), .C(n217), .Y(n2814) );
  OAI21X1 U2125 ( .A(n2348), .B(n2389), .C(n219), .Y(n2813) );
  OAI21X1 U2126 ( .A(n2348), .B(n2392), .C(n221), .Y(n2812) );
  OAI21X1 U2127 ( .A(n2348), .B(n2393), .C(n223), .Y(n2811) );
  OAI21X1 U2128 ( .A(n2348), .B(n2396), .C(n225), .Y(n2810) );
  OAI21X1 U2129 ( .A(n2348), .B(n2398), .C(n227), .Y(n2809) );
  OAI21X1 U2130 ( .A(n2348), .B(n2400), .C(n229), .Y(n2808) );
  OAI21X1 U2131 ( .A(n2348), .B(n2402), .C(n231), .Y(n2807) );
  OAI21X1 U2132 ( .A(n2348), .B(n2404), .C(n233), .Y(n2806) );
  OAI21X1 U2133 ( .A(n2349), .B(n2406), .C(n235), .Y(n2805) );
  OAI21X1 U2134 ( .A(n2349), .B(n2408), .C(n237), .Y(n2804) );
  OAI21X1 U2135 ( .A(n2349), .B(n2410), .C(n239), .Y(n2803) );
  OAI21X1 U2136 ( .A(n2349), .B(n2412), .C(n241), .Y(n2802) );
  OAI21X1 U2137 ( .A(n2349), .B(n2414), .C(n243), .Y(n2801) );
  OAI21X1 U2138 ( .A(n2349), .B(n2416), .C(n245), .Y(n2800) );
  OAI21X1 U2139 ( .A(n2349), .B(n2418), .C(n247), .Y(n2799) );
  OAI21X1 U2140 ( .A(n2349), .B(n2420), .C(n249), .Y(n2798) );
  OAI21X1 U2141 ( .A(n2350), .B(n2389), .C(n251), .Y(n2797) );
  OAI21X1 U2142 ( .A(n2350), .B(n2392), .C(n253), .Y(n2796) );
  OAI21X1 U2143 ( .A(n2350), .B(n2393), .C(n255), .Y(n2795) );
  OAI21X1 U2144 ( .A(n2350), .B(n2396), .C(n257), .Y(n2794) );
  OAI21X1 U2145 ( .A(n2350), .B(n2398), .C(n259), .Y(n2793) );
  OAI21X1 U2146 ( .A(n2350), .B(n2400), .C(n261), .Y(n2792) );
  OAI21X1 U2147 ( .A(n2350), .B(n2402), .C(n263), .Y(n2791) );
  OAI21X1 U2148 ( .A(n2350), .B(n2404), .C(n265), .Y(n2790) );
  OAI21X1 U2149 ( .A(n2351), .B(n2406), .C(n267), .Y(n2789) );
  OAI21X1 U2150 ( .A(n2351), .B(n2408), .C(n269), .Y(n2788) );
  OAI21X1 U2151 ( .A(n2351), .B(n2410), .C(n271), .Y(n2787) );
  OAI21X1 U2152 ( .A(n2351), .B(n2412), .C(n273), .Y(n2786) );
  OAI21X1 U2153 ( .A(n2351), .B(n2414), .C(n275), .Y(n2785) );
  OAI21X1 U2154 ( .A(n2351), .B(n2416), .C(n277), .Y(n2784) );
  OAI21X1 U2155 ( .A(n2351), .B(n2418), .C(n279), .Y(n2783) );
  OAI21X1 U2156 ( .A(n2351), .B(n2420), .C(n281), .Y(n2782) );
  OAI21X1 U2157 ( .A(n2352), .B(n2390), .C(n283), .Y(n2781) );
  OAI21X1 U2158 ( .A(n2352), .B(n2392), .C(n285), .Y(n2780) );
  OAI21X1 U2159 ( .A(n2352), .B(n2394), .C(n287), .Y(n2779) );
  OAI21X1 U2160 ( .A(n2352), .B(n2396), .C(n289), .Y(n2778) );
  OAI21X1 U2161 ( .A(n2352), .B(n2398), .C(n291), .Y(n2777) );
  OAI21X1 U2162 ( .A(n2352), .B(n2400), .C(n293), .Y(n2776) );
  OAI21X1 U2163 ( .A(n2352), .B(n2402), .C(n295), .Y(n2775) );
  OAI21X1 U2164 ( .A(n2352), .B(n2404), .C(n297), .Y(n2774) );
  OAI21X1 U2165 ( .A(n2353), .B(n2406), .C(n299), .Y(n2773) );
  OAI21X1 U2166 ( .A(n2353), .B(n2408), .C(n301), .Y(n2772) );
  OAI21X1 U2167 ( .A(n2353), .B(n2410), .C(n303), .Y(n2771) );
  OAI21X1 U2168 ( .A(n2353), .B(n2412), .C(n305), .Y(n2770) );
  OAI21X1 U2169 ( .A(n2353), .B(n2414), .C(n307), .Y(n2769) );
  OAI21X1 U2170 ( .A(n2353), .B(n2416), .C(n309), .Y(n2768) );
  OAI21X1 U2171 ( .A(n2353), .B(n2418), .C(n311), .Y(n2767) );
  OAI21X1 U2172 ( .A(n2353), .B(n2420), .C(n313), .Y(n2766) );
  OAI21X1 U2173 ( .A(n2354), .B(n2390), .C(n315), .Y(n2765) );
  OAI21X1 U2174 ( .A(n2354), .B(n2392), .C(n317), .Y(n2764) );
  OAI21X1 U2175 ( .A(n2354), .B(n2393), .C(n319), .Y(n2763) );
  OAI21X1 U2176 ( .A(n2354), .B(n2396), .C(n321), .Y(n2762) );
  OAI21X1 U2177 ( .A(n2354), .B(n2398), .C(n323), .Y(n2761) );
  OAI21X1 U2178 ( .A(n2354), .B(n2400), .C(n325), .Y(n2760) );
  OAI21X1 U2179 ( .A(n2354), .B(n2402), .C(n327), .Y(n2759) );
  OAI21X1 U2180 ( .A(n2354), .B(n2404), .C(n329), .Y(n2758) );
  OAI21X1 U2181 ( .A(n2355), .B(n2406), .C(n331), .Y(n2757) );
  OAI21X1 U2182 ( .A(n2355), .B(n2408), .C(n333), .Y(n2756) );
  OAI21X1 U2183 ( .A(n2355), .B(n2410), .C(n335), .Y(n2755) );
  OAI21X1 U2184 ( .A(n2355), .B(n2412), .C(n337), .Y(n2754) );
  OAI21X1 U2185 ( .A(n2355), .B(n2414), .C(n339), .Y(n2753) );
  OAI21X1 U2186 ( .A(n2355), .B(n2416), .C(n341), .Y(n2752) );
  OAI21X1 U2187 ( .A(n2355), .B(n2418), .C(n343), .Y(n2751) );
  OAI21X1 U2188 ( .A(n2355), .B(n2420), .C(n345), .Y(n2750) );
  OAI21X1 U2189 ( .A(n2356), .B(n2390), .C(n347), .Y(n2749) );
  OAI21X1 U2190 ( .A(n2356), .B(n2392), .C(n349), .Y(n2748) );
  OAI21X1 U2191 ( .A(n2356), .B(n2394), .C(n351), .Y(n2747) );
  OAI21X1 U2192 ( .A(n2356), .B(n2396), .C(n353), .Y(n2746) );
  OAI21X1 U2193 ( .A(n2356), .B(n2398), .C(n355), .Y(n2745) );
  OAI21X1 U2194 ( .A(n2356), .B(n2400), .C(n357), .Y(n2744) );
  OAI21X1 U2195 ( .A(n2356), .B(n2402), .C(n359), .Y(n2743) );
  OAI21X1 U2196 ( .A(n2356), .B(n2404), .C(n361), .Y(n2742) );
  OAI21X1 U2197 ( .A(n2357), .B(n2406), .C(n363), .Y(n2741) );
  OAI21X1 U2198 ( .A(n2357), .B(n2408), .C(n365), .Y(n2740) );
  OAI21X1 U2199 ( .A(n2357), .B(n2410), .C(n367), .Y(n2739) );
  OAI21X1 U2200 ( .A(n2357), .B(n2412), .C(n369), .Y(n2738) );
  OAI21X1 U2201 ( .A(n2357), .B(n2414), .C(n371), .Y(n2737) );
  OAI21X1 U2202 ( .A(n2357), .B(n2416), .C(n373), .Y(n2736) );
  OAI21X1 U2203 ( .A(n2357), .B(n2418), .C(n375), .Y(n2735) );
  OAI21X1 U2204 ( .A(n2357), .B(n2420), .C(n377), .Y(n2734) );
  OAI21X1 U2205 ( .A(n2358), .B(n2390), .C(n379), .Y(n2733) );
  OAI21X1 U2206 ( .A(n2358), .B(n2391), .C(n381), .Y(n2732) );
  OAI21X1 U2207 ( .A(n2358), .B(n2394), .C(n383), .Y(n2731) );
  OAI21X1 U2208 ( .A(n2358), .B(n2395), .C(n385), .Y(n2730) );
  OAI21X1 U2209 ( .A(n2358), .B(n2397), .C(n387), .Y(n2729) );
  OAI21X1 U2210 ( .A(n2358), .B(n2399), .C(n389), .Y(n2728) );
  OAI21X1 U2211 ( .A(n2358), .B(n2402), .C(n391), .Y(n2727) );
  OAI21X1 U2212 ( .A(n2358), .B(n2403), .C(n393), .Y(n2726) );
  OAI21X1 U2213 ( .A(n2358), .B(n2406), .C(n395), .Y(n2725) );
  OAI21X1 U2214 ( .A(n2358), .B(n2408), .C(n397), .Y(n2724) );
  OAI21X1 U2215 ( .A(n2358), .B(n2410), .C(n399), .Y(n2723) );
  OAI21X1 U2216 ( .A(n2358), .B(n2412), .C(n401), .Y(n2722) );
  OAI21X1 U2217 ( .A(n2358), .B(n2414), .C(n403), .Y(n2721) );
  OAI21X1 U2218 ( .A(n2358), .B(n2416), .C(n405), .Y(n2720) );
  OAI21X1 U2219 ( .A(n2358), .B(n2418), .C(n407), .Y(n2719) );
  OAI21X1 U2220 ( .A(n2358), .B(n2420), .C(n409), .Y(n2718) );
  NAND3X1 U2221 ( .A(n2427), .B(n2974), .C(n2430), .Y(n2450) );
  OAI21X1 U2222 ( .A(n2359), .B(n2390), .C(n411), .Y(n2717) );
  OAI21X1 U2223 ( .A(n2359), .B(n2392), .C(n413), .Y(n2716) );
  OAI21X1 U2224 ( .A(n2359), .B(n2393), .C(n415), .Y(n2715) );
  OAI21X1 U2225 ( .A(n2359), .B(n2396), .C(n417), .Y(n2714) );
  OAI21X1 U2226 ( .A(n2359), .B(n2398), .C(n419), .Y(n2713) );
  OAI21X1 U2227 ( .A(n2359), .B(n2400), .C(n421), .Y(n2712) );
  OAI21X1 U2228 ( .A(n2359), .B(n2402), .C(n423), .Y(n2711) );
  OAI21X1 U2229 ( .A(n2359), .B(n2404), .C(n425), .Y(n2710) );
  OAI21X1 U2230 ( .A(n2360), .B(n2406), .C(n427), .Y(n2709) );
  OAI21X1 U2231 ( .A(n2360), .B(n2408), .C(n429), .Y(n2708) );
  OAI21X1 U2232 ( .A(n2360), .B(n2410), .C(n431), .Y(n2707) );
  OAI21X1 U2233 ( .A(n2360), .B(n2412), .C(n433), .Y(n2706) );
  OAI21X1 U2234 ( .A(n2360), .B(n2414), .C(n435), .Y(n2705) );
  OAI21X1 U2235 ( .A(n2360), .B(n2416), .C(n437), .Y(n2704) );
  OAI21X1 U2236 ( .A(n2360), .B(n2418), .C(n439), .Y(n2703) );
  OAI21X1 U2237 ( .A(n2360), .B(n2420), .C(n441), .Y(n2702) );
  OAI21X1 U2238 ( .A(n2361), .B(n2390), .C(n443), .Y(n2701) );
  OAI21X1 U2239 ( .A(n2361), .B(n2392), .C(n445), .Y(n2700) );
  OAI21X1 U2240 ( .A(n2361), .B(n2393), .C(n447), .Y(n2699) );
  OAI21X1 U2241 ( .A(n2361), .B(n2396), .C(n449), .Y(n2698) );
  OAI21X1 U2242 ( .A(n2361), .B(n2398), .C(n451), .Y(n2697) );
  OAI21X1 U2243 ( .A(n2361), .B(n2400), .C(n453), .Y(n2696) );
  OAI21X1 U2244 ( .A(n2361), .B(n2402), .C(n455), .Y(n2695) );
  OAI21X1 U2245 ( .A(n2361), .B(n2404), .C(n457), .Y(n2694) );
  OAI21X1 U2246 ( .A(n2362), .B(n2406), .C(n459), .Y(n2693) );
  OAI21X1 U2247 ( .A(n2362), .B(n2408), .C(n461), .Y(n2692) );
  OAI21X1 U2248 ( .A(n2362), .B(n2410), .C(n463), .Y(n2691) );
  OAI21X1 U2249 ( .A(n2362), .B(n2412), .C(n465), .Y(n2690) );
  OAI21X1 U2250 ( .A(n2362), .B(n2414), .C(n467), .Y(n2689) );
  OAI21X1 U2251 ( .A(n2362), .B(n2416), .C(n469), .Y(n2688) );
  OAI21X1 U2252 ( .A(n2362), .B(n2418), .C(n471), .Y(n2687) );
  OAI21X1 U2253 ( .A(n2362), .B(n2420), .C(n473), .Y(n2686) );
  OAI21X1 U2254 ( .A(n2363), .B(n2390), .C(n475), .Y(n2685) );
  OAI21X1 U2255 ( .A(n2363), .B(n2392), .C(n477), .Y(n2684) );
  OAI21X1 U2256 ( .A(n2363), .B(n2393), .C(n479), .Y(n2683) );
  OAI21X1 U2257 ( .A(n2363), .B(n2396), .C(n481), .Y(n2682) );
  OAI21X1 U2258 ( .A(n2363), .B(n2398), .C(n483), .Y(n2681) );
  OAI21X1 U2259 ( .A(n2363), .B(n2400), .C(n485), .Y(n2680) );
  OAI21X1 U2260 ( .A(n2363), .B(n2402), .C(n487), .Y(n2679) );
  OAI21X1 U2261 ( .A(n2363), .B(n2404), .C(n489), .Y(n2678) );
  OAI21X1 U2262 ( .A(n2364), .B(n2406), .C(n491), .Y(n2677) );
  OAI21X1 U2263 ( .A(n2364), .B(n2408), .C(n493), .Y(n2676) );
  OAI21X1 U2264 ( .A(n2364), .B(n2410), .C(n495), .Y(n2675) );
  OAI21X1 U2265 ( .A(n2364), .B(n2412), .C(n497), .Y(n2674) );
  OAI21X1 U2266 ( .A(n2364), .B(n2414), .C(n499), .Y(n2673) );
  OAI21X1 U2267 ( .A(n2364), .B(n2416), .C(n501), .Y(n2672) );
  OAI21X1 U2268 ( .A(n2364), .B(n2418), .C(n503), .Y(n2671) );
  OAI21X1 U2269 ( .A(n2364), .B(n2420), .C(n505), .Y(n2670) );
  OAI21X1 U2270 ( .A(n2365), .B(n2390), .C(n507), .Y(n2669) );
  OAI21X1 U2271 ( .A(n2365), .B(n2392), .C(n509), .Y(n2668) );
  OAI21X1 U2272 ( .A(n2365), .B(n2394), .C(n511), .Y(n2667) );
  OAI21X1 U2273 ( .A(n2365), .B(n2396), .C(n513), .Y(n2666) );
  OAI21X1 U2274 ( .A(n2365), .B(n2398), .C(n515), .Y(n2665) );
  OAI21X1 U2275 ( .A(n2365), .B(n2400), .C(n517), .Y(n2664) );
  OAI21X1 U2276 ( .A(n2365), .B(n2402), .C(n519), .Y(n2663) );
  OAI21X1 U2277 ( .A(n2365), .B(n2404), .C(n521), .Y(n2662) );
  OAI21X1 U2278 ( .A(n2366), .B(n2406), .C(n523), .Y(n2661) );
  OAI21X1 U2279 ( .A(n2366), .B(n2408), .C(n525), .Y(n2660) );
  OAI21X1 U2280 ( .A(n2366), .B(n2410), .C(n527), .Y(n2659) );
  OAI21X1 U2281 ( .A(n2366), .B(n2412), .C(n529), .Y(n2658) );
  OAI21X1 U2282 ( .A(n2366), .B(n2414), .C(n531), .Y(n2657) );
  OAI21X1 U2283 ( .A(n2366), .B(n2416), .C(n533), .Y(n2656) );
  OAI21X1 U2284 ( .A(n2366), .B(n2418), .C(n535), .Y(n2655) );
  OAI21X1 U2285 ( .A(n2366), .B(n2420), .C(n537), .Y(n2654) );
  OAI21X1 U2286 ( .A(n2367), .B(n2390), .C(n539), .Y(n2653) );
  OAI21X1 U2287 ( .A(n2367), .B(n2391), .C(n541), .Y(n2652) );
  OAI21X1 U2288 ( .A(n2367), .B(n2393), .C(n543), .Y(n2651) );
  OAI21X1 U2289 ( .A(n2367), .B(n2395), .C(n545), .Y(n2650) );
  OAI21X1 U2290 ( .A(n2367), .B(n2397), .C(n547), .Y(n2649) );
  OAI21X1 U2291 ( .A(n2367), .B(n2399), .C(n549), .Y(n2648) );
  OAI21X1 U2292 ( .A(n2367), .B(n2401), .C(n551), .Y(n2647) );
  OAI21X1 U2293 ( .A(n2367), .B(n2403), .C(n553), .Y(n2646) );
  OAI21X1 U2294 ( .A(n2368), .B(n2405), .C(n555), .Y(n2645) );
  OAI21X1 U2295 ( .A(n2368), .B(n2407), .C(n557), .Y(n2644) );
  OAI21X1 U2296 ( .A(n2368), .B(n2409), .C(n559), .Y(n2643) );
  OAI21X1 U2297 ( .A(n2368), .B(n2411), .C(n561), .Y(n2642) );
  OAI21X1 U2298 ( .A(n2368), .B(n2413), .C(n563), .Y(n2641) );
  OAI21X1 U2299 ( .A(n2368), .B(n2415), .C(n565), .Y(n2640) );
  OAI21X1 U2300 ( .A(n2368), .B(n2417), .C(n567), .Y(n2639) );
  OAI21X1 U2301 ( .A(n2368), .B(n2419), .C(n569), .Y(n2638) );
  OAI21X1 U2302 ( .A(n2369), .B(n2390), .C(n571), .Y(n2637) );
  OAI21X1 U2303 ( .A(n2369), .B(n2391), .C(n573), .Y(n2636) );
  OAI21X1 U2304 ( .A(n2369), .B(n2393), .C(n575), .Y(n2635) );
  OAI21X1 U2305 ( .A(n2369), .B(n2395), .C(n577), .Y(n2634) );
  OAI21X1 U2306 ( .A(n2369), .B(n2397), .C(n579), .Y(n2633) );
  OAI21X1 U2307 ( .A(n2369), .B(n2399), .C(n581), .Y(n2632) );
  OAI21X1 U2308 ( .A(n2369), .B(n2401), .C(n583), .Y(n2631) );
  OAI21X1 U2309 ( .A(n2369), .B(n2403), .C(n585), .Y(n2630) );
  OAI21X1 U2310 ( .A(n2370), .B(n2405), .C(n587), .Y(n2629) );
  OAI21X1 U2311 ( .A(n2370), .B(n2407), .C(n589), .Y(n2628) );
  OAI21X1 U2312 ( .A(n2370), .B(n2409), .C(n591), .Y(n2627) );
  OAI21X1 U2313 ( .A(n2370), .B(n2411), .C(n593), .Y(n2626) );
  OAI21X1 U2314 ( .A(n2370), .B(n2413), .C(n595), .Y(n2625) );
  OAI21X1 U2315 ( .A(n2370), .B(n2415), .C(n597), .Y(n2624) );
  OAI21X1 U2316 ( .A(n2370), .B(n2417), .C(n599), .Y(n2623) );
  OAI21X1 U2317 ( .A(n2370), .B(n2419), .C(n601), .Y(n2622) );
  OAI21X1 U2318 ( .A(n2371), .B(n2390), .C(n603), .Y(n2621) );
  OAI21X1 U2319 ( .A(n2371), .B(n2391), .C(n605), .Y(n2620) );
  OAI21X1 U2320 ( .A(n2371), .B(n2393), .C(n607), .Y(n2619) );
  OAI21X1 U2321 ( .A(n2371), .B(n2395), .C(n609), .Y(n2618) );
  OAI21X1 U2322 ( .A(n2371), .B(n2397), .C(n611), .Y(n2617) );
  OAI21X1 U2323 ( .A(n2371), .B(n2399), .C(n613), .Y(n2616) );
  OAI21X1 U2324 ( .A(n2371), .B(n2401), .C(n615), .Y(n2615) );
  OAI21X1 U2325 ( .A(n2371), .B(n2403), .C(n617), .Y(n2614) );
  OAI21X1 U2326 ( .A(n2372), .B(n2405), .C(n619), .Y(n2613) );
  OAI21X1 U2327 ( .A(n2372), .B(n2407), .C(n621), .Y(n2612) );
  OAI21X1 U2328 ( .A(n2372), .B(n2409), .C(n623), .Y(n2611) );
  OAI21X1 U2329 ( .A(n2372), .B(n2411), .C(n625), .Y(n2610) );
  OAI21X1 U2330 ( .A(n2372), .B(n2413), .C(n627), .Y(n2609) );
  OAI21X1 U2331 ( .A(n2372), .B(n2415), .C(n629), .Y(n2608) );
  OAI21X1 U2332 ( .A(n2372), .B(n2417), .C(n631), .Y(n2607) );
  OAI21X1 U2333 ( .A(n2372), .B(n2419), .C(n633), .Y(n2606) );
  OAI21X1 U2334 ( .A(n2373), .B(n2390), .C(n635), .Y(n2605) );
  OAI21X1 U2335 ( .A(n2373), .B(n2391), .C(n637), .Y(n2604) );
  OAI21X1 U2336 ( .A(n2373), .B(n2394), .C(n639), .Y(n2603) );
  OAI21X1 U2337 ( .A(n2373), .B(n2395), .C(n641), .Y(n2602) );
  OAI21X1 U2338 ( .A(n2373), .B(n2397), .C(n643), .Y(n2601) );
  OAI21X1 U2339 ( .A(n2373), .B(n2399), .C(n645), .Y(n2600) );
  OAI21X1 U2340 ( .A(n2373), .B(n2401), .C(n647), .Y(n2599) );
  OAI21X1 U2341 ( .A(n2373), .B(n2403), .C(n649), .Y(n2598) );
  OAI21X1 U2342 ( .A(n2373), .B(n2405), .C(n1163), .Y(n2597) );
  OAI21X1 U2343 ( .A(n2373), .B(n2407), .C(n1165), .Y(n2596) );
  OAI21X1 U2344 ( .A(n2373), .B(n2409), .C(n1167), .Y(n2595) );
  OAI21X1 U2345 ( .A(n2373), .B(n2411), .C(n1169), .Y(n2594) );
  OAI21X1 U2346 ( .A(n2373), .B(n2413), .C(n1171), .Y(n2593) );
  OAI21X1 U2347 ( .A(n2373), .B(n2415), .C(n1173), .Y(n2592) );
  OAI21X1 U2348 ( .A(n2373), .B(n2417), .C(n1175), .Y(n2591) );
  OAI21X1 U2349 ( .A(n2373), .B(n2419), .C(n1177), .Y(n2590) );
  NAND3X1 U2350 ( .A(n2428), .B(n2974), .C(n2430), .Y(n2453) );
  OAI21X1 U2351 ( .A(n2374), .B(n2389), .C(n1662), .Y(n2589) );
  OAI21X1 U2352 ( .A(n2374), .B(n2391), .C(n1179), .Y(n2588) );
  OAI21X1 U2353 ( .A(n2374), .B(n2393), .C(n1181), .Y(n2587) );
  OAI21X1 U2354 ( .A(n2374), .B(n2395), .C(n1183), .Y(n2586) );
  OAI21X1 U2355 ( .A(n2374), .B(n2397), .C(n1185), .Y(n2585) );
  OAI21X1 U2356 ( .A(n2374), .B(n2399), .C(n1187), .Y(n2584) );
  OAI21X1 U2357 ( .A(n2374), .B(n2401), .C(n1189), .Y(n2583) );
  OAI21X1 U2358 ( .A(n2374), .B(n2403), .C(n1191), .Y(n2582) );
  OAI21X1 U2359 ( .A(n2375), .B(n2405), .C(n1193), .Y(n2581) );
  OAI21X1 U2360 ( .A(n2375), .B(n2407), .C(n1195), .Y(n2580) );
  OAI21X1 U2361 ( .A(n2375), .B(n2409), .C(n1197), .Y(n2579) );
  OAI21X1 U2362 ( .A(n2375), .B(n2411), .C(n1199), .Y(n2578) );
  OAI21X1 U2363 ( .A(n2375), .B(n2413), .C(n1201), .Y(n2577) );
  OAI21X1 U2364 ( .A(n2375), .B(n2415), .C(n1203), .Y(n2576) );
  OAI21X1 U2365 ( .A(n2375), .B(n2417), .C(n1205), .Y(n2575) );
  OAI21X1 U2366 ( .A(n2375), .B(n2419), .C(n1207), .Y(n2574) );
  OAI21X1 U2367 ( .A(n2376), .B(n2390), .C(n1664), .Y(n2573) );
  OAI21X1 U2368 ( .A(n2376), .B(n2391), .C(n1209), .Y(n2572) );
  OAI21X1 U2369 ( .A(n2376), .B(n2393), .C(n1211), .Y(n2571) );
  OAI21X1 U2370 ( .A(n2376), .B(n2395), .C(n1213), .Y(n2570) );
  OAI21X1 U2371 ( .A(n2376), .B(n2397), .C(n1215), .Y(n2569) );
  OAI21X1 U2372 ( .A(n2376), .B(n2399), .C(n1217), .Y(n2568) );
  OAI21X1 U2373 ( .A(n2376), .B(n2401), .C(n1219), .Y(n2567) );
  OAI21X1 U2374 ( .A(n2376), .B(n2403), .C(n1221), .Y(n2566) );
  OAI21X1 U2375 ( .A(n2377), .B(n2405), .C(n1223), .Y(n2565) );
  OAI21X1 U2376 ( .A(n2377), .B(n2407), .C(n1225), .Y(n2564) );
  OAI21X1 U2377 ( .A(n2377), .B(n2409), .C(n1227), .Y(n2563) );
  OAI21X1 U2378 ( .A(n2377), .B(n2411), .C(n1229), .Y(n2562) );
  OAI21X1 U2379 ( .A(n2377), .B(n2413), .C(n1231), .Y(n2561) );
  OAI21X1 U2380 ( .A(n2377), .B(n2415), .C(n1233), .Y(n2560) );
  OAI21X1 U2381 ( .A(n2377), .B(n2417), .C(n1235), .Y(n2559) );
  OAI21X1 U2382 ( .A(n2377), .B(n2419), .C(n1237), .Y(n2558) );
  OAI21X1 U2383 ( .A(n2378), .B(n2389), .C(n1666), .Y(n2557) );
  OAI21X1 U2384 ( .A(n2378), .B(n2391), .C(n1239), .Y(n2556) );
  OAI21X1 U2385 ( .A(n2378), .B(n2394), .C(n1241), .Y(n2555) );
  OAI21X1 U2386 ( .A(n2378), .B(n2395), .C(n1243), .Y(n2554) );
  OAI21X1 U2387 ( .A(n2378), .B(n2397), .C(n1245), .Y(n2553) );
  OAI21X1 U2388 ( .A(n2378), .B(n2399), .C(n1247), .Y(n2552) );
  OAI21X1 U2389 ( .A(n2378), .B(n2401), .C(n1249), .Y(n2551) );
  OAI21X1 U2390 ( .A(n2378), .B(n2403), .C(n1251), .Y(n2550) );
  OAI21X1 U2391 ( .A(n2379), .B(n2405), .C(n1253), .Y(n2549) );
  OAI21X1 U2392 ( .A(n2379), .B(n2407), .C(n1255), .Y(n2548) );
  OAI21X1 U2393 ( .A(n2379), .B(n2409), .C(n1257), .Y(n2547) );
  OAI21X1 U2394 ( .A(n2379), .B(n2411), .C(n1259), .Y(n2546) );
  OAI21X1 U2395 ( .A(n2379), .B(n2413), .C(n1261), .Y(n2545) );
  OAI21X1 U2396 ( .A(n2379), .B(n2415), .C(n1263), .Y(n2544) );
  OAI21X1 U2397 ( .A(n2379), .B(n2417), .C(n1265), .Y(n2543) );
  OAI21X1 U2398 ( .A(n2379), .B(n2419), .C(n1267), .Y(n2542) );
  OAI21X1 U2399 ( .A(n2380), .B(n2390), .C(n1668), .Y(n2541) );
  OAI21X1 U2400 ( .A(n2380), .B(n2391), .C(n1269), .Y(n2540) );
  OAI21X1 U2401 ( .A(n2380), .B(n2393), .C(n1271), .Y(n2539) );
  OAI21X1 U2402 ( .A(n2380), .B(n2395), .C(n1273), .Y(n2538) );
  OAI21X1 U2403 ( .A(n2380), .B(n2397), .C(n1275), .Y(n2537) );
  OAI21X1 U2404 ( .A(n2380), .B(n2399), .C(n1277), .Y(n2536) );
  OAI21X1 U2405 ( .A(n2380), .B(n2401), .C(n1279), .Y(n2535) );
  OAI21X1 U2406 ( .A(n2380), .B(n2403), .C(n1281), .Y(n2534) );
  OAI21X1 U2407 ( .A(n2381), .B(n2405), .C(n1283), .Y(n2533) );
  OAI21X1 U2408 ( .A(n2381), .B(n2407), .C(n1285), .Y(n2532) );
  OAI21X1 U2409 ( .A(n2381), .B(n2409), .C(n1287), .Y(n2531) );
  OAI21X1 U2410 ( .A(n2381), .B(n2411), .C(n1289), .Y(n2530) );
  OAI21X1 U2411 ( .A(n2381), .B(n2413), .C(n1291), .Y(n2529) );
  OAI21X1 U2412 ( .A(n2381), .B(n2415), .C(n1293), .Y(n2528) );
  OAI21X1 U2413 ( .A(n2381), .B(n2417), .C(n1295), .Y(n2527) );
  OAI21X1 U2414 ( .A(n2381), .B(n2419), .C(n1297), .Y(n2526) );
  OAI21X1 U2415 ( .A(n2382), .B(n2389), .C(n1670), .Y(n2525) );
  OAI21X1 U2416 ( .A(n2382), .B(n2391), .C(n1299), .Y(n2524) );
  OAI21X1 U2417 ( .A(n2382), .B(n2393), .C(n1301), .Y(n2523) );
  OAI21X1 U2418 ( .A(n2382), .B(n2395), .C(n1303), .Y(n2522) );
  OAI21X1 U2419 ( .A(n2382), .B(n2397), .C(n1305), .Y(n2521) );
  OAI21X1 U2420 ( .A(n2382), .B(n2399), .C(n1307), .Y(n2520) );
  OAI21X1 U2421 ( .A(n2382), .B(n2401), .C(n1309), .Y(n2519) );
  OAI21X1 U2422 ( .A(n2382), .B(n2403), .C(n1311), .Y(n2518) );
  OAI21X1 U2423 ( .A(n2383), .B(n2405), .C(n1313), .Y(n2517) );
  OAI21X1 U2424 ( .A(n2383), .B(n2407), .C(n1315), .Y(n2516) );
  OAI21X1 U2425 ( .A(n2383), .B(n2409), .C(n1317), .Y(n2515) );
  OAI21X1 U2426 ( .A(n2383), .B(n2411), .C(n1319), .Y(n2514) );
  OAI21X1 U2427 ( .A(n2383), .B(n2413), .C(n1321), .Y(n2513) );
  OAI21X1 U2428 ( .A(n2383), .B(n2415), .C(n1323), .Y(n2512) );
  OAI21X1 U2429 ( .A(n2383), .B(n2417), .C(n1325), .Y(n2511) );
  OAI21X1 U2430 ( .A(n2383), .B(n2419), .C(n1327), .Y(n2510) );
  OAI21X1 U2431 ( .A(n2384), .B(n2390), .C(n1672), .Y(n2509) );
  OAI21X1 U2432 ( .A(n2384), .B(n2391), .C(n1329), .Y(n2508) );
  OAI21X1 U2433 ( .A(n2384), .B(n2393), .C(n1331), .Y(n2507) );
  OAI21X1 U2434 ( .A(n2384), .B(n2395), .C(n1333), .Y(n2506) );
  OAI21X1 U2435 ( .A(n2384), .B(n2397), .C(n1335), .Y(n2505) );
  OAI21X1 U2436 ( .A(n2384), .B(n2399), .C(n1337), .Y(n2504) );
  OAI21X1 U2437 ( .A(n2384), .B(n2401), .C(n1339), .Y(n2503) );
  OAI21X1 U2438 ( .A(n2384), .B(n2403), .C(n1341), .Y(n2502) );
  OAI21X1 U2439 ( .A(n2385), .B(n2405), .C(n1343), .Y(n2501) );
  OAI21X1 U2440 ( .A(n2385), .B(n2407), .C(n1345), .Y(n2500) );
  OAI21X1 U2441 ( .A(n2385), .B(n2409), .C(n1347), .Y(n2499) );
  OAI21X1 U2442 ( .A(n2385), .B(n2411), .C(n1349), .Y(n2498) );
  OAI21X1 U2443 ( .A(n2385), .B(n2413), .C(n1351), .Y(n2497) );
  OAI21X1 U2444 ( .A(n2385), .B(n2415), .C(n1353), .Y(n2496) );
  OAI21X1 U2445 ( .A(n2385), .B(n2417), .C(n1355), .Y(n2495) );
  OAI21X1 U2446 ( .A(n2385), .B(n2419), .C(n1357), .Y(n2494) );
  OAI21X1 U2447 ( .A(n2386), .B(n2390), .C(n1674), .Y(n2493) );
  OAI21X1 U2448 ( .A(n2386), .B(n2391), .C(n1359), .Y(n2492) );
  OAI21X1 U2449 ( .A(n2386), .B(n2393), .C(n1361), .Y(n2491) );
  OAI21X1 U2450 ( .A(n2386), .B(n2395), .C(n1363), .Y(n2490) );
  OAI21X1 U2451 ( .A(n2386), .B(n2397), .C(n1365), .Y(n2489) );
  OAI21X1 U2452 ( .A(n2386), .B(n2399), .C(n1367), .Y(n2488) );
  OAI21X1 U2453 ( .A(n2386), .B(n2401), .C(n1369), .Y(n2487) );
  OAI21X1 U2454 ( .A(n2386), .B(n2403), .C(n1371), .Y(n2486) );
  OAI21X1 U2455 ( .A(n2387), .B(n2405), .C(n1373), .Y(n2485) );
  OAI21X1 U2456 ( .A(n2387), .B(n2407), .C(n1375), .Y(n2484) );
  OAI21X1 U2457 ( .A(n2387), .B(n2409), .C(n1377), .Y(n2483) );
  OAI21X1 U2458 ( .A(n2387), .B(n2411), .C(n1379), .Y(n2482) );
  OAI21X1 U2459 ( .A(n2387), .B(n2413), .C(n1381), .Y(n2481) );
  OAI21X1 U2460 ( .A(n2387), .B(n2415), .C(n1383), .Y(n2480) );
  OAI21X1 U2461 ( .A(n2387), .B(n2417), .C(n1385), .Y(n2479) );
  OAI21X1 U2462 ( .A(n2387), .B(n2419), .C(n1387), .Y(n2478) );
  OAI21X1 U2463 ( .A(n2388), .B(n2389), .C(n1676), .Y(n2477) );
  OAI21X1 U2464 ( .A(n2388), .B(n2391), .C(n1389), .Y(n2476) );
  OAI21X1 U2465 ( .A(n2388), .B(n2394), .C(n1391), .Y(n2475) );
  OAI21X1 U2466 ( .A(n2388), .B(n2395), .C(n1393), .Y(n2474) );
  OAI21X1 U2467 ( .A(n2388), .B(n2397), .C(n1395), .Y(n2473) );
  OAI21X1 U2468 ( .A(n2388), .B(n2399), .C(n1397), .Y(n2472) );
  OAI21X1 U2469 ( .A(n2388), .B(n2401), .C(n1399), .Y(n2471) );
  OAI21X1 U2470 ( .A(n2388), .B(n2403), .C(n1401), .Y(n2470) );
  OAI21X1 U2471 ( .A(n2388), .B(n2405), .C(n1403), .Y(n2469) );
  OAI21X1 U2472 ( .A(n2388), .B(n2407), .C(n1405), .Y(n2468) );
  OAI21X1 U2473 ( .A(n2388), .B(n2409), .C(n1407), .Y(n2467) );
  OAI21X1 U2474 ( .A(n2388), .B(n2411), .C(n1409), .Y(n2466) );
  OAI21X1 U2475 ( .A(n2388), .B(n2413), .C(n1411), .Y(n2465) );
  OAI21X1 U2476 ( .A(n2388), .B(n2415), .C(n1413), .Y(n2464) );
  OAI21X1 U2477 ( .A(n2388), .B(n2417), .C(n1415), .Y(n2463) );
  OAI21X1 U2478 ( .A(n2388), .B(n2419), .C(n1417), .Y(n2462) );
endmodule


module memc_Size16_5 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, net89253, net89251, net89385, net89383, net89545,
         net90019, net90763, net90761, net90943, \C2334/net90829 ,
         \C2334/net90835 , \C2334/net90347 , \C2334/net90349 ,
         \C2334/net90351 , \C2334/net90353 , \C2334/net90355 ,
         \C2334/net90357 , \C2334/net90359 , \C2334/net90363 ,
         \C2334/net90365 , \C2334/net90367 , \C2334/net90369 ,
         \C2334/net90371 , \C2334/net90373 , \C2334/net90375 ,
         \C2334/net90377 , \C2334/net90381 , \C2334/net90383 ,
         \C2334/net90385 , \C2334/net90387 , \C2334/net90389 ,
         \C2334/net90391 , \C2334/net90393 , \C2334/net90397 ,
         \C2334/net90399 , \C2334/net90401 , \C2334/net90405 ,
         \C2334/net90085 , \C2334/net89817 , \C2334/net89819 ,
         \C2334/net89821 , \C2334/net89823 , \C2334/net89825 ,
         \C2334/net89827 , \C2334/net89829 , \C2334/net89831 ,
         \C2334/net89833 , \C2334/net89835 , \C2334/net89837 ,
         \C2334/net89839 , \C2334/net89841 , \C2334/net89619 ,
         \C2334/net89621 , \C2334/net89623 , \C2334/net89625 ,
         \C2334/net89627 , \C2334/net89629 , \C2334/net89441 ,
         \C2334/net89443 , \C2334/net89445 , \C2334/net89303 ,
         \C2334/net89305 , net125642, net130272, net130271, N22, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n305, n307, n309, n311, n313, n315, n317, n319, n321,
         n323, n325, n327, n329, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;
  assign \data_out<10>  = net125642;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2052), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2053), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2054), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2055), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2056), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2057), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2058), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2059), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2060), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2061), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2062), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2063), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2064), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2065), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2066), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2067), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2068), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2069), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2070), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2071), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2072), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2073), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2074), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2075), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2076), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2077), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2078), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2079), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2080), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2081), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2082), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2083), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2084), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2085), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2086), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2087), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2088), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2089), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2090), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2091), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2092), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2093), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2094), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2095), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2096), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2097), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2098), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2099), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2100), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2101), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2102), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2103), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2104), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2105), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2106), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2107), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2108), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2109), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2110), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2111), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2112), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2113), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2114), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2115), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2116), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2117), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2118), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2119), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2120), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2121), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2122), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2123), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2124), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2125), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2126), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2127), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2128), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2129), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2130), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2131), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2132), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2133), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2134), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2135), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2136), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2137), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2138), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2139), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2140), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2141), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2142), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2143), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2144), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2145), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2146), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2147), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2148), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2149), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2150), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2151), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2152), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2153), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2154), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2155), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2156), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2157), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2158), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2159), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2160), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2161), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2162), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2163), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2164), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2165), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2166), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2167), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2168), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2169), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2170), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2171), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2172), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2173), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2174), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2175), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2176), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2177), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2178), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2179), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2180), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2181), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2182), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2183), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2184), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2185), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2186), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2187), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2188), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2189), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2190), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2191), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2192), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2193), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2194), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2195), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2196), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2197), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2198), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2199), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2200), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2201), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2202), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2203), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2204), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2205), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2206), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2207), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2208), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2209), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2210), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2211), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2212), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2213), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2214), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2215), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2216), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2217), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2218), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2219), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2220), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2221), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2222), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2223), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2224), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2225), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2226), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2227), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2228), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2229), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2230), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2231), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2232), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2233), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2234), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2235), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2236), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2237), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2238), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2239), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2240), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2241), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2242), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2243), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2244), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2245), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2246), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2247), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2248), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2249), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2250), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2251), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2252), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2253), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2254), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2255), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2256), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2257), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2258), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2259), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2260), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2261), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2262), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2263), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2264), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2265), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2266), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2267), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2268), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2269), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2270), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2271), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2272), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2273), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2274), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2275), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2276), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2277), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2278), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2279), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2280), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2281), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2282), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2283), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2284), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2285), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2286), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2287), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2288), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2289), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2290), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2291), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2292), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2293), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2294), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2295), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2296), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2297), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2298), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2299), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2300), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2301), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2302), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2303), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2304), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2305), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2306), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2307), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2308), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2309), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2310), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2311), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2312), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2313), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2314), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2315), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2316), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2317), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2318), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2319), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2320), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2321), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2322), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2323), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2324), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2325), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2326), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2327), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2328), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2329), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2330), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2331), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2332), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2333), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2334), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2335), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2336), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2337), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2338), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2339), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2340), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2341), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2342), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2343), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2344), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2345), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2346), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2347), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2348), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2349), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2350), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2351), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2352), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2353), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2354), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2355), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2356), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2357), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2358), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2359), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2360), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2361), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2362), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2363), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2364), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2365), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2366), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2367), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2368), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2369), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2370), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2371), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2372), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2373), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2374), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2375), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2376), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2377), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2378), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2379), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2380), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2381), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2382), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2383), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2384), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2385), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2386), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2387), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2388), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2389), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2390), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2391), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2392), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2393), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2394), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2395), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2396), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2397), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2398), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2399), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2400), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2401), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2402), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2403), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2404), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2405), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2406), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2407), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2408), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2409), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2410), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2411), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2412), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2413), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2414), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2415), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2416), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2417), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2418), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2419), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2420), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2421), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2422), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2423), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2424), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2425), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2426), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2427), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2428), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2429), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2430), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2431), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2432), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2433), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2434), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2435), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2436), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2437), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2438), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2439), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2440), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2441), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2442), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2443), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2444), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2445), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2446), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2447), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2448), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2449), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2450), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2451), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2452), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2453), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2454), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2455), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2456), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2457), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2458), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2459), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2460), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2461), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2462), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2463), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2464), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2465), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2466), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2467), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2468), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2469), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2470), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2471), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2472), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2473), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2474), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2475), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2476), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2477), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2478), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2479), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2480), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2481), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2482), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2483), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2484), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2485), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2486), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2487), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2488), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2489), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2490), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2491), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2492), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2493), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2494), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2495), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2496), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2497), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2498), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2499), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2500), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2501), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2502), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2503), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2504), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2505), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2506), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2507), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2508), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2509), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2510), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2511), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2512), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2513), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2514), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2515), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2516), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2517), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2518), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2519), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2520), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2521), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2522), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2523), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2524), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2525), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2526), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2527), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2528), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2529), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2530), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2531), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2532), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2533), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2534), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2535), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2536), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2537), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2538), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2539), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2540), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2541), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2542), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2543), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2544), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2545), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2546), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2547), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2548), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2549), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2550), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2551), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2552), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2553), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2554), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2555), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2556), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2557), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2558), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2559), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2560), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2561), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2562), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2563), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2564) );
  INVX1 U2 ( .A(write), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n422), .Y(n3) );
  INVX1 U5 ( .A(n421), .Y(n4) );
  INVX1 U6 ( .A(n420), .Y(n5) );
  AND2X2 U7 ( .A(n1646), .B(\data_in<15> ), .Y(n6) );
  INVX4 U8 ( .A(n424), .Y(n7) );
  INVX4 U9 ( .A(n424), .Y(n1678) );
  INVX2 U10 ( .A(n369), .Y(n8) );
  INVX2 U11 ( .A(n369), .Y(n9) );
  INVX2 U12 ( .A(n369), .Y(n370) );
  INVX2 U13 ( .A(n367), .Y(n10) );
  INVX2 U14 ( .A(n367), .Y(n11) );
  INVX2 U15 ( .A(n367), .Y(n368) );
  INVX2 U16 ( .A(n365), .Y(n12) );
  INVX2 U17 ( .A(n365), .Y(n13) );
  INVX2 U18 ( .A(n365), .Y(n366) );
  INVX2 U19 ( .A(n363), .Y(n14) );
  INVX2 U20 ( .A(n363), .Y(n15) );
  INVX2 U21 ( .A(n363), .Y(n364) );
  INVX2 U22 ( .A(n361), .Y(n16) );
  INVX2 U23 ( .A(n361), .Y(n17) );
  INVX2 U24 ( .A(n361), .Y(n362) );
  INVX2 U25 ( .A(n359), .Y(n18) );
  INVX2 U26 ( .A(n359), .Y(n19) );
  INVX2 U27 ( .A(n359), .Y(n360) );
  INVX2 U28 ( .A(n357), .Y(n20) );
  INVX2 U29 ( .A(n357), .Y(n21) );
  INVX2 U30 ( .A(n357), .Y(n358) );
  INVX2 U31 ( .A(n353), .Y(n22) );
  INVX2 U32 ( .A(n353), .Y(n23) );
  INVX2 U33 ( .A(n353), .Y(n354) );
  INVX2 U34 ( .A(n351), .Y(n24) );
  INVX2 U35 ( .A(n351), .Y(n25) );
  INVX2 U36 ( .A(n351), .Y(n352) );
  INVX2 U37 ( .A(n349), .Y(n26) );
  INVX2 U38 ( .A(n349), .Y(n27) );
  INVX2 U39 ( .A(n349), .Y(n350) );
  INVX2 U40 ( .A(n347), .Y(n28) );
  INVX2 U41 ( .A(n347), .Y(n29) );
  INVX2 U42 ( .A(n347), .Y(n348) );
  INVX2 U43 ( .A(n345), .Y(n30) );
  INVX2 U44 ( .A(n345), .Y(n31) );
  INVX2 U45 ( .A(n345), .Y(n346) );
  INVX2 U46 ( .A(n343), .Y(n32) );
  INVX2 U47 ( .A(n343), .Y(n33) );
  INVX2 U48 ( .A(n343), .Y(n344) );
  INVX2 U49 ( .A(n341), .Y(n34) );
  INVX2 U50 ( .A(n341), .Y(n35) );
  INVX2 U51 ( .A(n341), .Y(n342) );
  INVX2 U52 ( .A(n337), .Y(n36) );
  INVX2 U53 ( .A(n337), .Y(n37) );
  INVX2 U54 ( .A(n337), .Y(n338) );
  INVX2 U55 ( .A(n335), .Y(n38) );
  INVX2 U56 ( .A(n335), .Y(n39) );
  INVX2 U57 ( .A(n335), .Y(n336) );
  INVX2 U58 ( .A(n333), .Y(n40) );
  INVX2 U59 ( .A(n333), .Y(n41) );
  INVX2 U60 ( .A(n333), .Y(n334) );
  INVX2 U61 ( .A(n355), .Y(n42) );
  INVX2 U62 ( .A(n355), .Y(n43) );
  INVX2 U63 ( .A(n355), .Y(n356) );
  INVX1 U64 ( .A(n423), .Y(n44) );
  INVX1 U65 ( .A(n422), .Y(n45) );
  INVX1 U66 ( .A(n421), .Y(n46) );
  INVX1 U67 ( .A(n420), .Y(n47) );
  INVX2 U68 ( .A(n371), .Y(n48) );
  INVX2 U69 ( .A(n371), .Y(n49) );
  INVX2 U70 ( .A(n371), .Y(n372) );
  INVX8 U71 ( .A(n1647), .Y(n1646) );
  INVX1 U72 ( .A(net89545), .Y(\C2334/net89621 ) );
  INVX1 U73 ( .A(net89545), .Y(\C2334/net89623 ) );
  INVX1 U74 ( .A(net89545), .Y(\C2334/net89625 ) );
  INVX1 U75 ( .A(net89545), .Y(\C2334/net89627 ) );
  INVX1 U76 ( .A(net89253), .Y(\C2334/net89305 ) );
  INVX1 U77 ( .A(net89385), .Y(\C2334/net89445 ) );
  INVX1 U78 ( .A(net89385), .Y(\C2334/net89441 ) );
  INVX1 U79 ( .A(net89385), .Y(\C2334/net89443 ) );
  INVX1 U80 ( .A(net89253), .Y(\C2334/net89303 ) );
  INVX2 U81 ( .A(\C2334/net89841 ), .Y(\C2334/net89829 ) );
  INVX1 U82 ( .A(\C2334/net90085 ), .Y(\C2334/net89839 ) );
  INVX2 U83 ( .A(\C2334/net89841 ), .Y(\C2334/net89823 ) );
  INVX2 U84 ( .A(\C2334/net89839 ), .Y(\C2334/net89821 ) );
  INVX2 U85 ( .A(\C2334/net89841 ), .Y(\C2334/net89819 ) );
  INVX2 U86 ( .A(\C2334/net89839 ), .Y(\C2334/net89817 ) );
  INVX2 U87 ( .A(net90019), .Y(\C2334/net90085 ) );
  INVX1 U88 ( .A(net89545), .Y(\C2334/net89619 ) );
  INVX2 U89 ( .A(\C2334/net89841 ), .Y(\C2334/net89827 ) );
  INVX2 U90 ( .A(\C2334/net89839 ), .Y(\C2334/net89825 ) );
  INVX1 U91 ( .A(n1575), .Y(N26) );
  INVX1 U92 ( .A(n80), .Y(N22) );
  INVX1 U93 ( .A(n1580), .Y(N20) );
  INVX1 U94 ( .A(n1582), .Y(N18) );
  INVX1 U95 ( .A(n1569), .Y(N32) );
  INVX1 U96 ( .A(n1570), .Y(N31) );
  INVX1 U97 ( .A(n1571), .Y(N30) );
  INVX1 U98 ( .A(n1572), .Y(N29) );
  INVX1 U99 ( .A(n1573), .Y(N28) );
  INVX1 U100 ( .A(n1574), .Y(N27) );
  INVX1 U101 ( .A(n1576), .Y(N25) );
  INVX1 U102 ( .A(n1577), .Y(N24) );
  INVX1 U103 ( .A(n1578), .Y(N23) );
  INVX1 U104 ( .A(n1579), .Y(N21) );
  INVX1 U105 ( .A(n1581), .Y(N19) );
  INVX1 U106 ( .A(n1583), .Y(N17) );
  BUFX2 U107 ( .A(n552), .Y(n1585) );
  BUFX2 U108 ( .A(n554), .Y(n1587) );
  BUFX2 U109 ( .A(n556), .Y(n1589) );
  BUFX2 U110 ( .A(n558), .Y(n1591) );
  BUFX2 U111 ( .A(n560), .Y(n1593) );
  BUFX2 U112 ( .A(n562), .Y(n1595) );
  BUFX2 U113 ( .A(n564), .Y(n1597) );
  BUFX2 U114 ( .A(n566), .Y(n1600) );
  BUFX2 U115 ( .A(n568), .Y(n1602) );
  BUFX2 U116 ( .A(n570), .Y(n1604) );
  BUFX2 U117 ( .A(n572), .Y(n1606) );
  BUFX2 U118 ( .A(n574), .Y(n1608) );
  BUFX2 U119 ( .A(n576), .Y(n1610) );
  BUFX2 U120 ( .A(n578), .Y(n1612) );
  BUFX2 U121 ( .A(n580), .Y(n1615) );
  BUFX2 U122 ( .A(n582), .Y(n1617) );
  BUFX2 U123 ( .A(n584), .Y(n1619) );
  BUFX2 U124 ( .A(n586), .Y(n1621) );
  BUFX2 U125 ( .A(n588), .Y(n1623) );
  BUFX2 U126 ( .A(n590), .Y(n1625) );
  BUFX2 U127 ( .A(n592), .Y(n1627) );
  BUFX2 U128 ( .A(n594), .Y(n1630) );
  BUFX2 U129 ( .A(n596), .Y(n1632) );
  BUFX2 U130 ( .A(n598), .Y(n1634) );
  BUFX2 U131 ( .A(n600), .Y(n1636) );
  BUFX2 U132 ( .A(n602), .Y(n1638) );
  BUFX2 U133 ( .A(n604), .Y(n1640) );
  BUFX2 U134 ( .A(n606), .Y(n1642) );
  INVX1 U135 ( .A(n84), .Y(net125642) );
  OR2X2 U136 ( .A(write), .B(n83), .Y(n84) );
  INVX1 U137 ( .A(n82), .Y(n83) );
  AND2X1 U138 ( .A(N22), .B(net90943), .Y(n82) );
  MUX2X1 U139 ( .B(n77), .A(n62), .S(\C2334/net89303 ), .Y(n80) );
  MUX2X1 U140 ( .B(n78), .A(n79), .S(\C2334/net89443 ), .Y(n77) );
  MUX2X1 U141 ( .B(n74), .A(n71), .S(\C2334/net89625 ), .Y(n78) );
  MUX2X1 U142 ( .B(n75), .A(n76), .S(\C2334/net89823 ), .Y(n74) );
  MUX2X1 U143 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(\C2334/net90359 ), .Y(
        n75) );
  INVX8 U144 ( .A(\C2334/net90401 ), .Y(\C2334/net90359 ) );
  MUX2X1 U145 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(\C2334/net90359 ), .Y(
        n76) );
  MUX2X1 U146 ( .B(n72), .A(n73), .S(\C2334/net89823 ), .Y(n71) );
  MUX2X1 U147 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(\C2334/net90359 ), .Y(
        n72) );
  MUX2X1 U148 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(\C2334/net90359 ), .Y(
        n73) );
  MUX2X1 U149 ( .B(n68), .A(n65), .S(\C2334/net89625 ), .Y(n79) );
  MUX2X1 U150 ( .B(n69), .A(n70), .S(\C2334/net89823 ), .Y(n68) );
  MUX2X1 U151 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n81), .Y(n69) );
  INVX8 U152 ( .A(\C2334/net90399 ), .Y(n81) );
  MUX2X1 U153 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n81), .Y(n70) );
  MUX2X1 U154 ( .B(n66), .A(n67), .S(\C2334/net89823 ), .Y(n65) );
  MUX2X1 U155 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n81), .Y(n66) );
  MUX2X1 U156 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n81), .Y(n67) );
  MUX2X1 U157 ( .B(n63), .A(n64), .S(\C2334/net89443 ), .Y(n62) );
  MUX2X1 U158 ( .B(n59), .A(n56), .S(\C2334/net89625 ), .Y(n63) );
  MUX2X1 U159 ( .B(n60), .A(n61), .S(\C2334/net89823 ), .Y(n59) );
  MUX2X1 U160 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n81), .Y(n60) );
  MUX2X1 U161 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n81), .Y(n61) );
  MUX2X1 U162 ( .B(n57), .A(n58), .S(\C2334/net89823 ), .Y(n56) );
  MUX2X1 U163 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n81), .Y(n57) );
  MUX2X1 U164 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n81), .Y(n58) );
  MUX2X1 U165 ( .B(n53), .A(n50), .S(\C2334/net89625 ), .Y(n64) );
  MUX2X1 U166 ( .B(n54), .A(n55), .S(\C2334/net89823 ), .Y(n53) );
  MUX2X1 U167 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n81), .Y(n54) );
  MUX2X1 U168 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n81), .Y(n55) );
  MUX2X1 U169 ( .B(n51), .A(n52), .S(\C2334/net89823 ), .Y(n50) );
  MUX2X1 U170 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n81), .Y(n51) );
  MUX2X1 U171 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n81), .Y(n52) );
  INVX1 U172 ( .A(rst), .Y(net90943) );
  INVX2 U173 ( .A(\C2334/net89841 ), .Y(\C2334/net89831 ) );
  INVX1 U174 ( .A(net89545), .Y(\C2334/net89629 ) );
  INVX2 U175 ( .A(N12), .Y(net89545) );
  INVX2 U176 ( .A(net90761), .Y(\C2334/net90835 ) );
  INVX1 U177 ( .A(net89253), .Y(net89251) );
  INVX1 U178 ( .A(N14), .Y(net89253) );
  INVX1 U179 ( .A(net89385), .Y(net89383) );
  INVX1 U180 ( .A(N13), .Y(net89385) );
  INVX1 U181 ( .A(n549), .Y(n1629) );
  INVX1 U182 ( .A(n550), .Y(n1644) );
  BUFX2 U183 ( .A(n572), .Y(n1607) );
  BUFX2 U184 ( .A(n574), .Y(n1609) );
  BUFX2 U185 ( .A(n576), .Y(n1611) );
  BUFX2 U186 ( .A(n578), .Y(n1613) );
  BUFX2 U187 ( .A(n580), .Y(n1616) );
  BUFX2 U188 ( .A(n582), .Y(n1618) );
  BUFX2 U189 ( .A(n584), .Y(n1620) );
  BUFX2 U190 ( .A(n586), .Y(n1622) );
  BUFX2 U191 ( .A(n588), .Y(n1624) );
  BUFX2 U192 ( .A(n590), .Y(n1626) );
  BUFX2 U193 ( .A(n592), .Y(n1628) );
  BUFX2 U194 ( .A(n552), .Y(n1586) );
  BUFX2 U195 ( .A(n570), .Y(n1605) );
  BUFX2 U196 ( .A(n594), .Y(n1631) );
  BUFX2 U197 ( .A(n596), .Y(n1633) );
  BUFX2 U198 ( .A(n598), .Y(n1635) );
  BUFX2 U199 ( .A(n600), .Y(n1637) );
  BUFX2 U200 ( .A(n602), .Y(n1639) );
  BUFX2 U201 ( .A(n604), .Y(n1641) );
  BUFX2 U202 ( .A(n606), .Y(n1643) );
  BUFX2 U203 ( .A(n554), .Y(n1588) );
  BUFX2 U204 ( .A(n556), .Y(n1590) );
  BUFX2 U205 ( .A(n558), .Y(n1592) );
  BUFX2 U206 ( .A(n560), .Y(n1594) );
  BUFX2 U207 ( .A(n562), .Y(n1596) );
  BUFX2 U208 ( .A(n564), .Y(n1598) );
  BUFX2 U209 ( .A(n566), .Y(n1601) );
  BUFX2 U210 ( .A(n568), .Y(n1603) );
  INVX1 U211 ( .A(n548), .Y(n1614) );
  INVX1 U212 ( .A(n547), .Y(n1599) );
  INVX1 U213 ( .A(n423), .Y(n1676) );
  INVX1 U214 ( .A(n420), .Y(n1670) );
  INVX1 U215 ( .A(n421), .Y(n1672) );
  INVX1 U216 ( .A(n422), .Y(n1674) );
  INVX4 U217 ( .A(n1647), .Y(n1645) );
  INVX4 U218 ( .A(n1584), .Y(n1647) );
  INVX4 U219 ( .A(n389), .Y(n390) );
  INVX4 U220 ( .A(n407), .Y(n408) );
  INVX4 U221 ( .A(n405), .Y(n406) );
  INVX4 U222 ( .A(n401), .Y(n402) );
  INVX4 U223 ( .A(n399), .Y(n400) );
  INVX4 U224 ( .A(n397), .Y(n398) );
  INVX4 U225 ( .A(n395), .Y(n396) );
  INVX4 U226 ( .A(n393), .Y(n394) );
  INVX4 U227 ( .A(n391), .Y(n392) );
  INVX4 U228 ( .A(n403), .Y(n404) );
  INVX4 U229 ( .A(n301), .Y(n302) );
  AND2X2 U230 ( .A(net130271), .B(n515), .Y(\data_out<4> ) );
  INVX1 U231 ( .A(write), .Y(net130271) );
  INVX1 U232 ( .A(net130271), .Y(net130272) );
  AND2X2 U233 ( .A(\mem<20><8> ), .B(n332), .Y(n86) );
  INVX1 U234 ( .A(n86), .Y(n87) );
  AND2X2 U235 ( .A(\mem<20><9> ), .B(n332), .Y(n88) );
  INVX1 U236 ( .A(n88), .Y(n89) );
  AND2X2 U237 ( .A(\mem<20><10> ), .B(n332), .Y(n90) );
  INVX1 U238 ( .A(n90), .Y(n91) );
  AND2X2 U239 ( .A(\mem<20><11> ), .B(n332), .Y(n92) );
  INVX1 U240 ( .A(n92), .Y(n93) );
  AND2X2 U241 ( .A(\mem<20><12> ), .B(n332), .Y(n94) );
  INVX1 U242 ( .A(n94), .Y(n95) );
  AND2X2 U243 ( .A(\mem<20><13> ), .B(n332), .Y(n96) );
  INVX1 U244 ( .A(n96), .Y(n97) );
  AND2X2 U245 ( .A(\mem<20><14> ), .B(n332), .Y(n98) );
  INVX1 U246 ( .A(n98), .Y(n99) );
  AND2X2 U247 ( .A(\mem<19><8> ), .B(n334), .Y(n100) );
  INVX1 U248 ( .A(n100), .Y(n101) );
  AND2X2 U249 ( .A(\mem<19><9> ), .B(n40), .Y(n102) );
  INVX1 U250 ( .A(n102), .Y(n103) );
  AND2X2 U251 ( .A(n334), .B(\mem<19><10> ), .Y(n104) );
  INVX1 U252 ( .A(n104), .Y(n105) );
  AND2X2 U253 ( .A(\mem<19><11> ), .B(n334), .Y(n106) );
  INVX1 U254 ( .A(n106), .Y(n107) );
  AND2X2 U255 ( .A(\mem<19><12> ), .B(n40), .Y(n108) );
  INVX1 U256 ( .A(n108), .Y(n109) );
  AND2X2 U257 ( .A(\mem<19><13> ), .B(n334), .Y(n110) );
  INVX1 U258 ( .A(n110), .Y(n111) );
  AND2X2 U259 ( .A(\mem<19><14> ), .B(n334), .Y(n112) );
  INVX1 U260 ( .A(n112), .Y(n113) );
  AND2X2 U261 ( .A(\mem<18><8> ), .B(n336), .Y(n114) );
  INVX1 U262 ( .A(n114), .Y(n115) );
  AND2X2 U263 ( .A(\mem<18><9> ), .B(n38), .Y(n116) );
  INVX1 U264 ( .A(n116), .Y(n117) );
  AND2X2 U265 ( .A(n336), .B(\mem<18><10> ), .Y(n118) );
  INVX1 U266 ( .A(n118), .Y(n119) );
  AND2X2 U267 ( .A(\mem<18><11> ), .B(n336), .Y(n120) );
  INVX1 U268 ( .A(n120), .Y(n121) );
  AND2X2 U269 ( .A(\mem<18><12> ), .B(n38), .Y(n122) );
  INVX1 U270 ( .A(n122), .Y(n123) );
  AND2X2 U271 ( .A(\mem<18><13> ), .B(n336), .Y(n124) );
  INVX1 U272 ( .A(n124), .Y(n125) );
  AND2X2 U273 ( .A(\mem<18><14> ), .B(n336), .Y(n126) );
  INVX1 U274 ( .A(n126), .Y(n127) );
  AND2X2 U275 ( .A(\mem<17><8> ), .B(n338), .Y(n128) );
  INVX1 U276 ( .A(n128), .Y(n129) );
  AND2X2 U277 ( .A(\mem<17><9> ), .B(n36), .Y(n130) );
  INVX1 U278 ( .A(n130), .Y(n131) );
  AND2X2 U279 ( .A(n338), .B(\mem<17><10> ), .Y(n132) );
  INVX1 U280 ( .A(n132), .Y(n133) );
  AND2X2 U281 ( .A(\mem<17><11> ), .B(n338), .Y(n134) );
  INVX1 U282 ( .A(n134), .Y(n135) );
  AND2X2 U283 ( .A(\mem<17><12> ), .B(n36), .Y(n136) );
  INVX1 U284 ( .A(n136), .Y(n137) );
  AND2X2 U285 ( .A(\mem<17><13> ), .B(n338), .Y(n138) );
  INVX1 U286 ( .A(n138), .Y(n139) );
  AND2X2 U287 ( .A(\mem<17><14> ), .B(n338), .Y(n140) );
  INVX1 U288 ( .A(n140), .Y(n141) );
  AND2X2 U289 ( .A(\mem<16><8> ), .B(n340), .Y(n142) );
  INVX1 U290 ( .A(n142), .Y(n143) );
  AND2X2 U291 ( .A(\mem<16><9> ), .B(n340), .Y(n144) );
  INVX1 U292 ( .A(n144), .Y(n145) );
  AND2X2 U293 ( .A(\mem<16><10> ), .B(n340), .Y(n146) );
  INVX1 U294 ( .A(n146), .Y(n147) );
  AND2X2 U295 ( .A(\mem<16><11> ), .B(n340), .Y(n148) );
  INVX1 U296 ( .A(n148), .Y(n149) );
  AND2X2 U297 ( .A(\mem<16><12> ), .B(n340), .Y(n150) );
  INVX1 U298 ( .A(n150), .Y(n151) );
  AND2X2 U299 ( .A(\mem<16><13> ), .B(n340), .Y(n152) );
  INVX1 U300 ( .A(n152), .Y(n153) );
  AND2X2 U301 ( .A(\mem<16><15> ), .B(n340), .Y(n154) );
  INVX1 U302 ( .A(n154), .Y(n155) );
  AND2X2 U303 ( .A(\mem<15><8> ), .B(n342), .Y(n156) );
  INVX1 U304 ( .A(n156), .Y(n157) );
  AND2X2 U305 ( .A(\mem<15><9> ), .B(n34), .Y(n158) );
  INVX1 U306 ( .A(n158), .Y(n159) );
  AND2X2 U307 ( .A(n342), .B(\mem<15><10> ), .Y(n160) );
  INVX1 U308 ( .A(n160), .Y(n161) );
  AND2X2 U309 ( .A(\mem<15><11> ), .B(n342), .Y(n162) );
  INVX1 U310 ( .A(n162), .Y(n163) );
  AND2X2 U311 ( .A(\mem<15><12> ), .B(n34), .Y(n164) );
  INVX1 U312 ( .A(n164), .Y(n165) );
  AND2X2 U313 ( .A(\mem<15><13> ), .B(n342), .Y(n166) );
  INVX1 U314 ( .A(n166), .Y(n167) );
  AND2X2 U315 ( .A(\mem<15><14> ), .B(n342), .Y(n168) );
  INVX1 U316 ( .A(n168), .Y(n169) );
  AND2X2 U317 ( .A(\mem<14><8> ), .B(n344), .Y(n170) );
  INVX1 U318 ( .A(n170), .Y(n171) );
  AND2X2 U319 ( .A(\mem<14><9> ), .B(n32), .Y(n172) );
  INVX1 U320 ( .A(n172), .Y(n173) );
  AND2X2 U321 ( .A(n344), .B(\mem<14><10> ), .Y(n174) );
  INVX1 U322 ( .A(n174), .Y(n175) );
  AND2X2 U323 ( .A(\mem<14><11> ), .B(n344), .Y(n176) );
  INVX1 U324 ( .A(n176), .Y(n177) );
  AND2X2 U325 ( .A(\mem<14><12> ), .B(n32), .Y(n178) );
  INVX1 U326 ( .A(n178), .Y(n179) );
  AND2X2 U327 ( .A(\mem<14><13> ), .B(n344), .Y(n180) );
  INVX1 U328 ( .A(n180), .Y(n181) );
  AND2X2 U329 ( .A(\mem<14><14> ), .B(n344), .Y(n182) );
  INVX1 U330 ( .A(n182), .Y(n183) );
  AND2X2 U331 ( .A(\mem<13><8> ), .B(n346), .Y(n184) );
  INVX1 U332 ( .A(n184), .Y(n185) );
  AND2X2 U333 ( .A(\mem<13><9> ), .B(n30), .Y(n186) );
  INVX1 U334 ( .A(n186), .Y(n187) );
  AND2X2 U335 ( .A(n346), .B(\mem<13><10> ), .Y(n188) );
  INVX1 U336 ( .A(n188), .Y(n189) );
  AND2X2 U337 ( .A(\mem<13><11> ), .B(n346), .Y(n190) );
  INVX1 U338 ( .A(n190), .Y(n191) );
  AND2X2 U339 ( .A(\mem<13><12> ), .B(n30), .Y(n192) );
  INVX1 U340 ( .A(n192), .Y(n193) );
  AND2X2 U341 ( .A(\mem<13><13> ), .B(n346), .Y(n194) );
  INVX1 U342 ( .A(n194), .Y(n195) );
  AND2X2 U343 ( .A(\mem<13><14> ), .B(n346), .Y(n196) );
  INVX1 U344 ( .A(n196), .Y(n197) );
  AND2X2 U345 ( .A(\mem<12><8> ), .B(n348), .Y(n198) );
  INVX1 U346 ( .A(n198), .Y(n199) );
  AND2X2 U347 ( .A(\mem<12><9> ), .B(n28), .Y(n200) );
  INVX1 U348 ( .A(n200), .Y(n201) );
  AND2X2 U349 ( .A(n348), .B(\mem<12><10> ), .Y(n202) );
  INVX1 U350 ( .A(n202), .Y(n203) );
  AND2X2 U351 ( .A(\mem<12><11> ), .B(n348), .Y(n204) );
  INVX1 U352 ( .A(n204), .Y(n205) );
  AND2X2 U353 ( .A(\mem<12><12> ), .B(n28), .Y(n206) );
  INVX1 U354 ( .A(n206), .Y(n207) );
  AND2X2 U355 ( .A(\mem<12><13> ), .B(n348), .Y(n208) );
  INVX1 U356 ( .A(n208), .Y(n209) );
  AND2X2 U357 ( .A(\mem<12><14> ), .B(n348), .Y(n210) );
  INVX1 U358 ( .A(n210), .Y(n211) );
  AND2X2 U359 ( .A(\mem<11><8> ), .B(n350), .Y(n212) );
  INVX1 U360 ( .A(n212), .Y(n213) );
  AND2X2 U361 ( .A(\mem<11><9> ), .B(n26), .Y(n215) );
  INVX1 U362 ( .A(n215), .Y(n216) );
  AND2X2 U363 ( .A(n350), .B(\mem<11><10> ), .Y(n217) );
  INVX1 U364 ( .A(n217), .Y(n218) );
  AND2X2 U365 ( .A(\mem<11><11> ), .B(n350), .Y(n219) );
  INVX1 U366 ( .A(n219), .Y(n220) );
  AND2X2 U367 ( .A(\mem<11><12> ), .B(n26), .Y(n221) );
  INVX1 U368 ( .A(n221), .Y(n222) );
  AND2X2 U369 ( .A(\mem<11><13> ), .B(n350), .Y(n223) );
  INVX1 U370 ( .A(n223), .Y(n224) );
  AND2X2 U371 ( .A(\mem<11><14> ), .B(n350), .Y(n225) );
  INVX1 U372 ( .A(n225), .Y(n226) );
  AND2X2 U373 ( .A(\mem<10><8> ), .B(n352), .Y(n227) );
  INVX1 U374 ( .A(n227), .Y(n228) );
  AND2X2 U375 ( .A(\mem<10><9> ), .B(n24), .Y(n229) );
  INVX1 U376 ( .A(n229), .Y(n230) );
  AND2X2 U377 ( .A(n352), .B(\mem<10><10> ), .Y(n231) );
  INVX1 U378 ( .A(n231), .Y(n232) );
  AND2X2 U379 ( .A(\mem<10><11> ), .B(n352), .Y(n233) );
  INVX1 U380 ( .A(n233), .Y(n234) );
  AND2X2 U381 ( .A(\mem<10><12> ), .B(n24), .Y(n235) );
  INVX1 U382 ( .A(n235), .Y(n236) );
  AND2X2 U383 ( .A(\mem<10><13> ), .B(n352), .Y(n237) );
  INVX1 U384 ( .A(n237), .Y(n238) );
  AND2X2 U385 ( .A(\mem<10><14> ), .B(n352), .Y(n239) );
  INVX1 U386 ( .A(n239), .Y(n240) );
  AND2X2 U387 ( .A(\mem<9><8> ), .B(n354), .Y(n241) );
  INVX1 U388 ( .A(n241), .Y(n242) );
  AND2X2 U389 ( .A(\mem<9><9> ), .B(n22), .Y(n243) );
  INVX1 U390 ( .A(n243), .Y(n244) );
  AND2X2 U391 ( .A(n354), .B(\mem<9><10> ), .Y(n245) );
  INVX1 U392 ( .A(n245), .Y(n246) );
  AND2X2 U393 ( .A(\mem<9><11> ), .B(n354), .Y(n247) );
  INVX1 U394 ( .A(n247), .Y(n248) );
  AND2X2 U395 ( .A(\mem<9><12> ), .B(n22), .Y(n249) );
  INVX1 U396 ( .A(n249), .Y(n250) );
  AND2X2 U397 ( .A(\mem<9><13> ), .B(n354), .Y(n251) );
  INVX1 U398 ( .A(n251), .Y(n252) );
  AND2X2 U399 ( .A(\mem<9><14> ), .B(n354), .Y(n253) );
  INVX1 U400 ( .A(n253), .Y(n254) );
  AND2X2 U401 ( .A(\mem<8><8> ), .B(n356), .Y(n255) );
  INVX1 U402 ( .A(n255), .Y(n256) );
  AND2X2 U403 ( .A(\mem<8><9> ), .B(n43), .Y(n257) );
  INVX1 U404 ( .A(n257), .Y(n258) );
  AND2X2 U405 ( .A(\mem<7><8> ), .B(n358), .Y(n259) );
  INVX1 U406 ( .A(n259), .Y(n260) );
  AND2X2 U407 ( .A(n21), .B(\mem<7><9> ), .Y(n261) );
  INVX1 U408 ( .A(n261), .Y(n262) );
  AND2X2 U409 ( .A(\mem<6><8> ), .B(n360), .Y(n263) );
  INVX1 U410 ( .A(n263), .Y(n264) );
  AND2X2 U411 ( .A(n19), .B(\mem<6><9> ), .Y(n265) );
  INVX1 U412 ( .A(n265), .Y(n266) );
  AND2X2 U413 ( .A(\mem<5><8> ), .B(n362), .Y(n267) );
  INVX1 U414 ( .A(n267), .Y(n268) );
  AND2X2 U415 ( .A(n17), .B(\mem<5><9> ), .Y(n269) );
  INVX1 U416 ( .A(n269), .Y(n270) );
  AND2X2 U417 ( .A(\mem<4><8> ), .B(n364), .Y(n271) );
  INVX1 U418 ( .A(n271), .Y(n272) );
  AND2X2 U419 ( .A(n15), .B(\mem<4><9> ), .Y(n273) );
  INVX1 U420 ( .A(n273), .Y(n274) );
  AND2X2 U421 ( .A(\mem<3><8> ), .B(n366), .Y(n275) );
  INVX1 U422 ( .A(n275), .Y(n276) );
  AND2X2 U423 ( .A(n13), .B(\mem<3><9> ), .Y(n277) );
  INVX1 U424 ( .A(n277), .Y(n278) );
  AND2X2 U425 ( .A(\mem<2><8> ), .B(n368), .Y(n279) );
  INVX1 U426 ( .A(n279), .Y(n280) );
  AND2X2 U427 ( .A(n11), .B(\mem<2><9> ), .Y(n281) );
  INVX1 U428 ( .A(n281), .Y(n282) );
  AND2X2 U429 ( .A(\mem<1><8> ), .B(n370), .Y(n283) );
  INVX1 U430 ( .A(n283), .Y(n284) );
  AND2X2 U431 ( .A(n9), .B(\mem<1><9> ), .Y(n285) );
  INVX1 U432 ( .A(n285), .Y(n286) );
  AND2X2 U433 ( .A(\mem<0><8> ), .B(n372), .Y(n287) );
  INVX1 U434 ( .A(n287), .Y(n288) );
  AND2X2 U435 ( .A(\mem<0><9> ), .B(n372), .Y(n289) );
  INVX1 U436 ( .A(n289), .Y(n290) );
  AND2X2 U437 ( .A(\mem<0><10> ), .B(n372), .Y(n291) );
  INVX1 U438 ( .A(n291), .Y(n292) );
  AND2X2 U439 ( .A(\mem<0><11> ), .B(n372), .Y(n293) );
  INVX1 U440 ( .A(n293), .Y(n294) );
  AND2X2 U441 ( .A(\mem<0><12> ), .B(n372), .Y(n295) );
  INVX1 U442 ( .A(n295), .Y(n296) );
  AND2X2 U443 ( .A(\mem<0><13> ), .B(n372), .Y(n297) );
  INVX1 U444 ( .A(n297), .Y(n298) );
  AND2X2 U445 ( .A(\mem<0><15> ), .B(n49), .Y(n299) );
  INVX1 U446 ( .A(n299), .Y(n300) );
  AND2X2 U447 ( .A(n1645), .B(n569), .Y(n301) );
  INVX4 U448 ( .A(n331), .Y(n332) );
  INVX4 U449 ( .A(n339), .Y(n340) );
  OR2X2 U450 ( .A(write), .B(n508), .Y(n303) );
  INVX1 U451 ( .A(n303), .Y(\data_out<0> ) );
  OR2X2 U452 ( .A(write), .B(n510), .Y(n305) );
  INVX1 U453 ( .A(n305), .Y(\data_out<1> ) );
  OR2X2 U454 ( .A(write), .B(n512), .Y(n307) );
  INVX1 U455 ( .A(n307), .Y(\data_out<2> ) );
  OR2X2 U456 ( .A(write), .B(n514), .Y(n309) );
  INVX1 U457 ( .A(n309), .Y(\data_out<3> ) );
  OR2X2 U458 ( .A(write), .B(n517), .Y(n311) );
  INVX1 U459 ( .A(n311), .Y(\data_out<5> ) );
  OR2X2 U460 ( .A(write), .B(n519), .Y(n313) );
  INVX1 U461 ( .A(n313), .Y(\data_out<6> ) );
  OR2X2 U462 ( .A(write), .B(n533), .Y(n315) );
  INVX1 U463 ( .A(n315), .Y(\data_out<7> ) );
  OR2X2 U464 ( .A(n2), .B(n535), .Y(n317) );
  INVX1 U465 ( .A(n317), .Y(\data_out<8> ) );
  OR2X2 U466 ( .A(write), .B(n521), .Y(n319) );
  INVX1 U467 ( .A(n319), .Y(\data_out<9> ) );
  OR2X2 U468 ( .A(write), .B(n523), .Y(n321) );
  INVX1 U469 ( .A(n321), .Y(\data_out<11> ) );
  OR2X2 U470 ( .A(write), .B(n525), .Y(n323) );
  INVX1 U471 ( .A(n323), .Y(\data_out<12> ) );
  OR2X2 U472 ( .A(write), .B(n527), .Y(n325) );
  INVX1 U473 ( .A(n325), .Y(\data_out<13> ) );
  OR2X2 U474 ( .A(write), .B(n529), .Y(n327) );
  INVX1 U475 ( .A(n327), .Y(\data_out<14> ) );
  OR2X2 U476 ( .A(write), .B(n531), .Y(n329) );
  INVX1 U477 ( .A(n329), .Y(\data_out<15> ) );
  AND2X2 U478 ( .A(n1646), .B(n571), .Y(n331) );
  AND2X2 U479 ( .A(n1645), .B(n573), .Y(n333) );
  AND2X2 U480 ( .A(n1645), .B(n575), .Y(n335) );
  AND2X2 U481 ( .A(n1645), .B(n577), .Y(n337) );
  AND2X2 U482 ( .A(n1645), .B(n548), .Y(n339) );
  AND2X2 U483 ( .A(n1645), .B(n579), .Y(n341) );
  AND2X2 U484 ( .A(n1645), .B(n581), .Y(n343) );
  AND2X2 U485 ( .A(n1645), .B(n583), .Y(n345) );
  AND2X2 U486 ( .A(n1645), .B(n585), .Y(n347) );
  AND2X2 U487 ( .A(n1645), .B(n587), .Y(n349) );
  AND2X2 U488 ( .A(n1645), .B(n589), .Y(n351) );
  AND2X2 U489 ( .A(n1645), .B(n591), .Y(n353) );
  AND2X2 U490 ( .A(n1645), .B(n549), .Y(n355) );
  AND2X2 U491 ( .A(n1645), .B(n593), .Y(n357) );
  AND2X2 U492 ( .A(n1645), .B(n595), .Y(n359) );
  AND2X2 U493 ( .A(n1645), .B(n597), .Y(n361) );
  AND2X2 U494 ( .A(n1645), .B(n599), .Y(n363) );
  AND2X2 U495 ( .A(n1645), .B(n601), .Y(n365) );
  AND2X2 U496 ( .A(n1645), .B(n603), .Y(n367) );
  AND2X2 U497 ( .A(n1645), .B(n605), .Y(n369) );
  AND2X2 U498 ( .A(n1646), .B(n550), .Y(n371) );
  AND2X2 U499 ( .A(\mem<8><10> ), .B(n356), .Y(n373) );
  INVX1 U500 ( .A(n373), .Y(n374) );
  AND2X2 U501 ( .A(\mem<7><10> ), .B(n358), .Y(n375) );
  INVX1 U502 ( .A(n375), .Y(n376) );
  AND2X2 U503 ( .A(\mem<6><10> ), .B(n360), .Y(n377) );
  INVX1 U504 ( .A(n377), .Y(n378) );
  AND2X2 U505 ( .A(\mem<5><10> ), .B(n362), .Y(n379) );
  INVX1 U506 ( .A(n379), .Y(n380) );
  AND2X2 U507 ( .A(\mem<4><10> ), .B(n364), .Y(n381) );
  INVX1 U508 ( .A(n381), .Y(n382) );
  AND2X2 U509 ( .A(\mem<3><10> ), .B(n366), .Y(n383) );
  INVX1 U510 ( .A(n383), .Y(n384) );
  AND2X2 U511 ( .A(\mem<2><10> ), .B(n368), .Y(n385) );
  INVX1 U512 ( .A(n385), .Y(n386) );
  AND2X2 U513 ( .A(\mem<1><10> ), .B(n370), .Y(n387) );
  INVX1 U514 ( .A(n387), .Y(n388) );
  AND2X2 U515 ( .A(n1645), .B(n551), .Y(n389) );
  AND2X2 U516 ( .A(n1645), .B(n553), .Y(n391) );
  AND2X2 U517 ( .A(n1645), .B(n555), .Y(n393) );
  AND2X2 U518 ( .A(n1645), .B(n557), .Y(n395) );
  AND2X2 U519 ( .A(n1645), .B(n559), .Y(n397) );
  AND2X2 U520 ( .A(n1645), .B(n561), .Y(n399) );
  AND2X2 U521 ( .A(n1645), .B(n563), .Y(n401) );
  AND2X2 U522 ( .A(n1645), .B(n547), .Y(n403) );
  AND2X2 U523 ( .A(n1645), .B(n565), .Y(n405) );
  AND2X2 U524 ( .A(n1646), .B(n567), .Y(n407) );
  AND2X2 U525 ( .A(n1646), .B(\data_in<0> ), .Y(n409) );
  AND2X2 U526 ( .A(n1646), .B(\data_in<1> ), .Y(n410) );
  AND2X2 U527 ( .A(n1646), .B(\data_in<2> ), .Y(n411) );
  AND2X2 U528 ( .A(n1646), .B(\data_in<3> ), .Y(n412) );
  AND2X2 U529 ( .A(n1646), .B(\data_in<4> ), .Y(n413) );
  AND2X2 U530 ( .A(n1646), .B(\data_in<5> ), .Y(n414) );
  AND2X2 U531 ( .A(n1646), .B(\data_in<6> ), .Y(n415) );
  AND2X2 U532 ( .A(n1646), .B(\data_in<7> ), .Y(n416) );
  AND2X2 U533 ( .A(n1646), .B(\data_in<8> ), .Y(n417) );
  AND2X2 U534 ( .A(n1646), .B(\data_in<9> ), .Y(n418) );
  AND2X2 U535 ( .A(n1646), .B(\data_in<10> ), .Y(n419) );
  AND2X2 U536 ( .A(n1646), .B(\data_in<11> ), .Y(n420) );
  AND2X2 U537 ( .A(n1646), .B(\data_in<12> ), .Y(n421) );
  AND2X2 U538 ( .A(n1646), .B(\data_in<13> ), .Y(n422) );
  AND2X2 U539 ( .A(n1646), .B(\data_in<14> ), .Y(n423) );
  AND2X2 U540 ( .A(n1646), .B(\data_in<15> ), .Y(n424) );
  AND2X2 U541 ( .A(\mem<8><11> ), .B(n43), .Y(n425) );
  INVX1 U542 ( .A(n425), .Y(n426) );
  AND2X2 U543 ( .A(n42), .B(\mem<8><12> ), .Y(n427) );
  INVX1 U544 ( .A(n427), .Y(n428) );
  AND2X2 U545 ( .A(n43), .B(\mem<8><13> ), .Y(n429) );
  INVX1 U546 ( .A(n429), .Y(n430) );
  AND2X2 U547 ( .A(\mem<8><14> ), .B(n356), .Y(n431) );
  INVX1 U548 ( .A(n431), .Y(n432) );
  AND2X2 U549 ( .A(n42), .B(\mem<8><15> ), .Y(n433) );
  INVX1 U550 ( .A(n433), .Y(n434) );
  AND2X2 U551 ( .A(\mem<7><11> ), .B(n20), .Y(n435) );
  INVX1 U552 ( .A(n435), .Y(n436) );
  AND2X2 U553 ( .A(\mem<7><12> ), .B(n358), .Y(n437) );
  INVX1 U554 ( .A(n437), .Y(n438) );
  AND2X2 U555 ( .A(\mem<7><13> ), .B(n20), .Y(n439) );
  INVX1 U556 ( .A(n439), .Y(n440) );
  AND2X2 U557 ( .A(\mem<7><14> ), .B(n358), .Y(n441) );
  INVX1 U558 ( .A(n441), .Y(n442) );
  AND2X2 U559 ( .A(\mem<7><15> ), .B(n358), .Y(n443) );
  INVX1 U560 ( .A(n443), .Y(n444) );
  AND2X2 U561 ( .A(\mem<6><11> ), .B(n18), .Y(n445) );
  INVX1 U562 ( .A(n445), .Y(n446) );
  AND2X2 U563 ( .A(\mem<6><12> ), .B(n360), .Y(n447) );
  INVX1 U564 ( .A(n447), .Y(n448) );
  AND2X2 U565 ( .A(\mem<6><13> ), .B(n18), .Y(n449) );
  INVX1 U566 ( .A(n449), .Y(n450) );
  AND2X2 U567 ( .A(\mem<6><14> ), .B(n360), .Y(n451) );
  INVX1 U568 ( .A(n451), .Y(n452) );
  AND2X2 U569 ( .A(\mem<6><15> ), .B(n360), .Y(n453) );
  INVX1 U570 ( .A(n453), .Y(n454) );
  AND2X2 U571 ( .A(\mem<5><11> ), .B(n16), .Y(n455) );
  INVX1 U572 ( .A(n455), .Y(n456) );
  AND2X2 U573 ( .A(\mem<5><12> ), .B(n362), .Y(n457) );
  INVX1 U574 ( .A(n457), .Y(n458) );
  AND2X2 U575 ( .A(\mem<5><13> ), .B(n16), .Y(n459) );
  INVX1 U576 ( .A(n459), .Y(n460) );
  AND2X2 U577 ( .A(\mem<5><14> ), .B(n362), .Y(n461) );
  INVX1 U578 ( .A(n461), .Y(n462) );
  AND2X2 U579 ( .A(\mem<5><15> ), .B(n362), .Y(n463) );
  INVX1 U580 ( .A(n463), .Y(n464) );
  AND2X2 U581 ( .A(\mem<4><11> ), .B(n14), .Y(n465) );
  INVX1 U582 ( .A(n465), .Y(n466) );
  AND2X2 U583 ( .A(\mem<4><12> ), .B(n364), .Y(n467) );
  INVX1 U584 ( .A(n467), .Y(n468) );
  AND2X2 U585 ( .A(\mem<4><13> ), .B(n14), .Y(n469) );
  INVX1 U586 ( .A(n469), .Y(n470) );
  AND2X2 U587 ( .A(\mem<4><14> ), .B(n364), .Y(n471) );
  INVX1 U588 ( .A(n471), .Y(n472) );
  AND2X2 U589 ( .A(\mem<4><15> ), .B(n364), .Y(n473) );
  INVX1 U590 ( .A(n473), .Y(n474) );
  AND2X2 U591 ( .A(\mem<3><11> ), .B(n12), .Y(n475) );
  INVX1 U592 ( .A(n475), .Y(n476) );
  AND2X2 U593 ( .A(\mem<3><12> ), .B(n366), .Y(n477) );
  INVX1 U594 ( .A(n477), .Y(n478) );
  AND2X2 U595 ( .A(\mem<3><13> ), .B(n12), .Y(n479) );
  INVX1 U596 ( .A(n479), .Y(n480) );
  AND2X2 U597 ( .A(\mem<3><14> ), .B(n366), .Y(n481) );
  INVX1 U598 ( .A(n481), .Y(n482) );
  AND2X2 U599 ( .A(\mem<3><15> ), .B(n366), .Y(n483) );
  INVX1 U600 ( .A(n483), .Y(n484) );
  AND2X2 U601 ( .A(\mem<2><11> ), .B(n10), .Y(n485) );
  INVX1 U602 ( .A(n485), .Y(n486) );
  AND2X2 U603 ( .A(\mem<2><12> ), .B(n368), .Y(n487) );
  INVX1 U604 ( .A(n487), .Y(n488) );
  AND2X2 U605 ( .A(\mem<2><13> ), .B(n10), .Y(n489) );
  INVX1 U606 ( .A(n489), .Y(n490) );
  AND2X2 U607 ( .A(\mem<2><14> ), .B(n368), .Y(n491) );
  INVX1 U608 ( .A(n491), .Y(n492) );
  AND2X2 U609 ( .A(\mem<2><15> ), .B(n368), .Y(n493) );
  INVX1 U610 ( .A(n493), .Y(n494) );
  AND2X2 U611 ( .A(\mem<1><11> ), .B(n8), .Y(n495) );
  INVX1 U612 ( .A(n495), .Y(n496) );
  AND2X2 U613 ( .A(\mem<1><12> ), .B(n370), .Y(n497) );
  INVX1 U614 ( .A(n497), .Y(n498) );
  AND2X2 U615 ( .A(\mem<1><13> ), .B(n8), .Y(n499) );
  INVX1 U616 ( .A(n499), .Y(n500) );
  AND2X2 U617 ( .A(\mem<1><14> ), .B(n370), .Y(n501) );
  INVX1 U618 ( .A(n501), .Y(n502) );
  AND2X2 U619 ( .A(\mem<1><15> ), .B(n370), .Y(n503) );
  INVX1 U620 ( .A(n503), .Y(n504) );
  INVX1 U621 ( .A(net90763), .Y(net90761) );
  AND2X1 U622 ( .A(\C2334/net89629 ), .B(\C2334/net89831 ), .Y(n505) );
  AND2X1 U623 ( .A(n2564), .B(net89251), .Y(n506) );
  AND2X1 U624 ( .A(N32), .B(net90943), .Y(n507) );
  INVX1 U625 ( .A(n507), .Y(n508) );
  AND2X1 U626 ( .A(N31), .B(net90943), .Y(n509) );
  INVX1 U627 ( .A(n509), .Y(n510) );
  AND2X1 U628 ( .A(N30), .B(net90943), .Y(n511) );
  INVX1 U629 ( .A(n511), .Y(n512) );
  AND2X1 U630 ( .A(N29), .B(net90943), .Y(n513) );
  INVX1 U631 ( .A(n513), .Y(n514) );
  AND2X1 U632 ( .A(N28), .B(net90943), .Y(n515) );
  AND2X1 U633 ( .A(N27), .B(net90943), .Y(n516) );
  INVX1 U634 ( .A(n516), .Y(n517) );
  AND2X1 U635 ( .A(N26), .B(net90943), .Y(n518) );
  INVX1 U636 ( .A(n518), .Y(n519) );
  AND2X1 U637 ( .A(N23), .B(net90943), .Y(n520) );
  INVX1 U638 ( .A(n520), .Y(n521) );
  AND2X1 U639 ( .A(N21), .B(net90943), .Y(n522) );
  INVX1 U640 ( .A(n522), .Y(n523) );
  AND2X1 U641 ( .A(N20), .B(net90943), .Y(n524) );
  INVX1 U642 ( .A(n524), .Y(n525) );
  AND2X1 U643 ( .A(N19), .B(net90943), .Y(n526) );
  INVX1 U644 ( .A(n526), .Y(n527) );
  AND2X1 U645 ( .A(N18), .B(net90943), .Y(n528) );
  INVX1 U646 ( .A(n528), .Y(n529) );
  AND2X1 U647 ( .A(N17), .B(net90943), .Y(n530) );
  INVX1 U648 ( .A(n530), .Y(n531) );
  AND2X1 U649 ( .A(N25), .B(net90943), .Y(n532) );
  INVX1 U650 ( .A(n532), .Y(n533) );
  AND2X1 U651 ( .A(N24), .B(net90943), .Y(n534) );
  INVX1 U652 ( .A(n534), .Y(n535) );
  BUFX2 U653 ( .A(n1712), .Y(n536) );
  INVX1 U654 ( .A(n536), .Y(n1996) );
  BUFX2 U655 ( .A(n1729), .Y(n537) );
  INVX1 U656 ( .A(n537), .Y(n2005) );
  BUFX2 U657 ( .A(n1746), .Y(n538) );
  INVX1 U658 ( .A(n538), .Y(n2014) );
  BUFX2 U659 ( .A(n1763), .Y(n539) );
  INVX1 U660 ( .A(n539), .Y(n2023) );
  BUFX2 U661 ( .A(n1780), .Y(n540) );
  INVX1 U662 ( .A(n540), .Y(n2032) );
  BUFX2 U663 ( .A(n1906), .Y(n541) );
  INVX1 U664 ( .A(n541), .Y(n1970) );
  BUFX2 U665 ( .A(n1979), .Y(n542) );
  INVX1 U666 ( .A(n542), .Y(n2041) );
  AND2X1 U667 ( .A(net90761), .B(n505), .Y(n543) );
  AND2X1 U668 ( .A(net89383), .B(n506), .Y(n544) );
  AND2X1 U669 ( .A(net90763), .B(n505), .Y(n545) );
  AND2X1 U670 ( .A(net89385), .B(n506), .Y(n546) );
  AND2X1 U671 ( .A(n544), .B(n2042), .Y(n547) );
  AND2X1 U672 ( .A(n2042), .B(n546), .Y(n548) );
  AND2X1 U673 ( .A(n2042), .B(n1970), .Y(n549) );
  AND2X1 U674 ( .A(n2042), .B(n2041), .Y(n550) );
  AND2X1 U675 ( .A(n543), .B(n544), .Y(n551) );
  INVX1 U676 ( .A(n551), .Y(n552) );
  AND2X1 U677 ( .A(n544), .B(n545), .Y(n553) );
  INVX1 U678 ( .A(n553), .Y(n554) );
  AND2X1 U679 ( .A(n544), .B(n1996), .Y(n555) );
  INVX1 U680 ( .A(n555), .Y(n556) );
  AND2X1 U681 ( .A(n544), .B(n2005), .Y(n557) );
  INVX1 U682 ( .A(n557), .Y(n558) );
  AND2X1 U683 ( .A(n544), .B(n2014), .Y(n559) );
  INVX1 U684 ( .A(n559), .Y(n560) );
  AND2X1 U685 ( .A(n544), .B(n2023), .Y(n561) );
  INVX1 U686 ( .A(n561), .Y(n562) );
  AND2X1 U687 ( .A(n544), .B(n2032), .Y(n563) );
  INVX1 U688 ( .A(n563), .Y(n564) );
  AND2X1 U689 ( .A(n543), .B(n546), .Y(n565) );
  INVX1 U690 ( .A(n565), .Y(n566) );
  AND2X1 U691 ( .A(n545), .B(n546), .Y(n567) );
  INVX1 U692 ( .A(n567), .Y(n568) );
  AND2X1 U693 ( .A(n1996), .B(n546), .Y(n569) );
  INVX1 U694 ( .A(n569), .Y(n570) );
  AND2X1 U695 ( .A(n2005), .B(n546), .Y(n571) );
  INVX1 U696 ( .A(n571), .Y(n572) );
  AND2X1 U697 ( .A(n2014), .B(n546), .Y(n573) );
  INVX1 U698 ( .A(n573), .Y(n574) );
  AND2X1 U699 ( .A(n2023), .B(n546), .Y(n575) );
  INVX1 U700 ( .A(n575), .Y(n576) );
  AND2X1 U701 ( .A(n2032), .B(n546), .Y(n577) );
  INVX1 U702 ( .A(n577), .Y(n578) );
  AND2X1 U703 ( .A(n543), .B(n1970), .Y(n579) );
  INVX1 U704 ( .A(n579), .Y(n580) );
  AND2X1 U705 ( .A(n545), .B(n1970), .Y(n581) );
  INVX1 U706 ( .A(n581), .Y(n582) );
  AND2X1 U707 ( .A(n1996), .B(n1970), .Y(n583) );
  INVX1 U708 ( .A(n583), .Y(n584) );
  AND2X1 U709 ( .A(n2005), .B(n1970), .Y(n585) );
  INVX1 U710 ( .A(n585), .Y(n586) );
  AND2X1 U711 ( .A(n2014), .B(n1970), .Y(n587) );
  INVX1 U712 ( .A(n587), .Y(n588) );
  AND2X1 U713 ( .A(n2023), .B(n1970), .Y(n589) );
  INVX1 U714 ( .A(n589), .Y(n590) );
  AND2X1 U715 ( .A(n2032), .B(n1970), .Y(n591) );
  INVX1 U716 ( .A(n591), .Y(n592) );
  AND2X1 U717 ( .A(n543), .B(n2041), .Y(n593) );
  INVX1 U718 ( .A(n593), .Y(n594) );
  AND2X1 U719 ( .A(n545), .B(n2041), .Y(n595) );
  INVX1 U720 ( .A(n595), .Y(n596) );
  AND2X1 U721 ( .A(n1996), .B(n2041), .Y(n597) );
  INVX1 U722 ( .A(n597), .Y(n598) );
  AND2X1 U723 ( .A(n2005), .B(n2041), .Y(n599) );
  INVX1 U724 ( .A(n599), .Y(n600) );
  AND2X1 U725 ( .A(n2014), .B(n2041), .Y(n601) );
  INVX1 U726 ( .A(n601), .Y(n602) );
  AND2X1 U727 ( .A(n2023), .B(n2041), .Y(n603) );
  INVX1 U728 ( .A(n603), .Y(n604) );
  AND2X1 U729 ( .A(n2032), .B(n2041), .Y(n605) );
  INVX1 U730 ( .A(n605), .Y(n606) );
  INVX1 U731 ( .A(N11), .Y(net90019) );
  MUX2X1 U732 ( .B(n608), .A(n609), .S(\C2334/net89837 ), .Y(n607) );
  MUX2X1 U733 ( .B(n611), .A(n612), .S(\C2334/net89837 ), .Y(n610) );
  MUX2X1 U734 ( .B(n614), .A(n615), .S(\C2334/net89837 ), .Y(n613) );
  MUX2X1 U735 ( .B(n617), .A(n618), .S(\C2334/net89837 ), .Y(n616) );
  MUX2X1 U736 ( .B(n620), .A(n621), .S(\C2334/net89441 ), .Y(n619) );
  MUX2X1 U737 ( .B(n623), .A(n624), .S(\C2334/net89837 ), .Y(n622) );
  MUX2X1 U738 ( .B(n626), .A(n627), .S(\C2334/net89837 ), .Y(n625) );
  MUX2X1 U739 ( .B(n629), .A(n630), .S(\C2334/net89837 ), .Y(n628) );
  MUX2X1 U740 ( .B(n632), .A(n633), .S(\C2334/net89837 ), .Y(n631) );
  MUX2X1 U741 ( .B(n635), .A(n636), .S(\C2334/net89441 ), .Y(n634) );
  MUX2X1 U742 ( .B(n638), .A(n639), .S(\C2334/net89835 ), .Y(n637) );
  MUX2X1 U743 ( .B(n641), .A(n642), .S(\C2334/net89835 ), .Y(n640) );
  MUX2X1 U744 ( .B(n644), .A(n645), .S(\C2334/net89835 ), .Y(n643) );
  MUX2X1 U745 ( .B(n647), .A(n648), .S(\C2334/net89835 ), .Y(n646) );
  MUX2X1 U746 ( .B(n650), .A(n1163), .S(\C2334/net89441 ), .Y(n649) );
  MUX2X1 U747 ( .B(n1165), .A(n1166), .S(\C2334/net89835 ), .Y(n1164) );
  MUX2X1 U748 ( .B(n1168), .A(n1169), .S(\C2334/net89835 ), .Y(n1167) );
  MUX2X1 U749 ( .B(n1171), .A(n1172), .S(\C2334/net89835 ), .Y(n1170) );
  MUX2X1 U750 ( .B(n1174), .A(n1175), .S(\C2334/net89835 ), .Y(n1173) );
  MUX2X1 U751 ( .B(n1177), .A(n1178), .S(\C2334/net89441 ), .Y(n1176) );
  MUX2X1 U752 ( .B(n1180), .A(n1181), .S(\C2334/net89835 ), .Y(n1179) );
  MUX2X1 U753 ( .B(n1183), .A(n1184), .S(\C2334/net89835 ), .Y(n1182) );
  MUX2X1 U754 ( .B(n1186), .A(n1187), .S(\C2334/net89835 ), .Y(n1185) );
  MUX2X1 U755 ( .B(n1189), .A(n1190), .S(\C2334/net89835 ), .Y(n1188) );
  MUX2X1 U756 ( .B(n1192), .A(n1193), .S(\C2334/net89441 ), .Y(n1191) );
  MUX2X1 U757 ( .B(n1195), .A(n1196), .S(\C2334/net89833 ), .Y(n1194) );
  MUX2X1 U758 ( .B(n1198), .A(n1199), .S(\C2334/net89833 ), .Y(n1197) );
  MUX2X1 U759 ( .B(n1201), .A(n1202), .S(\C2334/net89833 ), .Y(n1200) );
  MUX2X1 U760 ( .B(n1204), .A(n1205), .S(\C2334/net89833 ), .Y(n1203) );
  MUX2X1 U761 ( .B(n1207), .A(n1208), .S(\C2334/net89441 ), .Y(n1206) );
  MUX2X1 U762 ( .B(n1210), .A(n1211), .S(\C2334/net89833 ), .Y(n1209) );
  MUX2X1 U763 ( .B(n1213), .A(n1214), .S(\C2334/net89833 ), .Y(n1212) );
  MUX2X1 U764 ( .B(n1216), .A(n1217), .S(\C2334/net89833 ), .Y(n1215) );
  MUX2X1 U765 ( .B(n1219), .A(n1220), .S(\C2334/net89833 ), .Y(n1218) );
  MUX2X1 U766 ( .B(n1222), .A(n1223), .S(\C2334/net89441 ), .Y(n1221) );
  MUX2X1 U767 ( .B(n1225), .A(n1226), .S(\C2334/net89833 ), .Y(n1224) );
  MUX2X1 U768 ( .B(n1228), .A(n1229), .S(\C2334/net89833 ), .Y(n1227) );
  MUX2X1 U769 ( .B(n1231), .A(n1232), .S(\C2334/net89833 ), .Y(n1230) );
  MUX2X1 U770 ( .B(n1234), .A(n1235), .S(\C2334/net89833 ), .Y(n1233) );
  MUX2X1 U771 ( .B(n1237), .A(n1238), .S(\C2334/net89441 ), .Y(n1236) );
  MUX2X1 U772 ( .B(n1240), .A(n1241), .S(\C2334/net89831 ), .Y(n1239) );
  MUX2X1 U773 ( .B(n1243), .A(n1244), .S(\C2334/net89831 ), .Y(n1242) );
  MUX2X1 U774 ( .B(n1246), .A(n1247), .S(\C2334/net89831 ), .Y(n1245) );
  MUX2X1 U775 ( .B(n1249), .A(n1250), .S(\C2334/net89831 ), .Y(n1248) );
  MUX2X1 U776 ( .B(n1252), .A(n1253), .S(\C2334/net89441 ), .Y(n1251) );
  MUX2X1 U777 ( .B(n1255), .A(n1256), .S(\C2334/net89831 ), .Y(n1254) );
  MUX2X1 U778 ( .B(n1258), .A(n1259), .S(\C2334/net89831 ), .Y(n1257) );
  MUX2X1 U779 ( .B(n1261), .A(n1262), .S(\C2334/net89831 ), .Y(n1260) );
  MUX2X1 U780 ( .B(n1264), .A(n1265), .S(\C2334/net89831 ), .Y(n1263) );
  MUX2X1 U781 ( .B(n1267), .A(n1268), .S(\C2334/net89441 ), .Y(n1266) );
  MUX2X1 U782 ( .B(n1270), .A(n1271), .S(\C2334/net89831 ), .Y(n1269) );
  MUX2X1 U783 ( .B(n1273), .A(n1274), .S(\C2334/net89831 ), .Y(n1272) );
  MUX2X1 U784 ( .B(n1276), .A(n1277), .S(\C2334/net89831 ), .Y(n1275) );
  MUX2X1 U785 ( .B(n1279), .A(n1280), .S(\C2334/net89831 ), .Y(n1278) );
  MUX2X1 U786 ( .B(n1282), .A(n1283), .S(\C2334/net89441 ), .Y(n1281) );
  MUX2X1 U787 ( .B(n1285), .A(n1286), .S(\C2334/net89829 ), .Y(n1284) );
  MUX2X1 U788 ( .B(n1288), .A(n1289), .S(\C2334/net89829 ), .Y(n1287) );
  MUX2X1 U789 ( .B(n1291), .A(n1292), .S(\C2334/net89829 ), .Y(n1290) );
  MUX2X1 U790 ( .B(n1294), .A(n1295), .S(\C2334/net89829 ), .Y(n1293) );
  MUX2X1 U791 ( .B(n1297), .A(n1298), .S(\C2334/net89441 ), .Y(n1296) );
  MUX2X1 U792 ( .B(n1300), .A(n1301), .S(\C2334/net89829 ), .Y(n1299) );
  MUX2X1 U793 ( .B(n1303), .A(n1304), .S(\C2334/net89829 ), .Y(n1302) );
  MUX2X1 U794 ( .B(n1306), .A(n1307), .S(\C2334/net89829 ), .Y(n1305) );
  MUX2X1 U795 ( .B(n1309), .A(n1310), .S(\C2334/net89829 ), .Y(n1308) );
  MUX2X1 U796 ( .B(n1312), .A(n1313), .S(\C2334/net89443 ), .Y(n1311) );
  MUX2X1 U797 ( .B(n1315), .A(n1316), .S(\C2334/net89829 ), .Y(n1314) );
  MUX2X1 U798 ( .B(n1318), .A(n1319), .S(\C2334/net89829 ), .Y(n1317) );
  MUX2X1 U799 ( .B(n1321), .A(n1322), .S(\C2334/net89829 ), .Y(n1320) );
  MUX2X1 U800 ( .B(n1324), .A(n1325), .S(\C2334/net89829 ), .Y(n1323) );
  MUX2X1 U801 ( .B(n1327), .A(n1328), .S(\C2334/net89443 ), .Y(n1326) );
  MUX2X1 U802 ( .B(n1330), .A(n1331), .S(\C2334/net89827 ), .Y(n1329) );
  MUX2X1 U803 ( .B(n1333), .A(n1334), .S(\C2334/net89827 ), .Y(n1332) );
  MUX2X1 U804 ( .B(n1336), .A(n1337), .S(\C2334/net89827 ), .Y(n1335) );
  MUX2X1 U805 ( .B(n1339), .A(n1340), .S(\C2334/net89827 ), .Y(n1338) );
  MUX2X1 U806 ( .B(n1342), .A(n1343), .S(\C2334/net89443 ), .Y(n1341) );
  MUX2X1 U807 ( .B(n1345), .A(n1346), .S(\C2334/net89827 ), .Y(n1344) );
  MUX2X1 U808 ( .B(n1348), .A(n1349), .S(\C2334/net89827 ), .Y(n1347) );
  MUX2X1 U809 ( .B(n1351), .A(n1352), .S(\C2334/net89827 ), .Y(n1350) );
  MUX2X1 U810 ( .B(n1354), .A(n1355), .S(\C2334/net89827 ), .Y(n1353) );
  MUX2X1 U811 ( .B(n1357), .A(n1358), .S(\C2334/net89443 ), .Y(n1356) );
  MUX2X1 U812 ( .B(n1360), .A(n1361), .S(\C2334/net89827 ), .Y(n1359) );
  MUX2X1 U813 ( .B(n1363), .A(n1364), .S(\C2334/net89827 ), .Y(n1362) );
  MUX2X1 U814 ( .B(n1366), .A(n1367), .S(\C2334/net89827 ), .Y(n1365) );
  MUX2X1 U815 ( .B(n1369), .A(n1370), .S(\C2334/net89827 ), .Y(n1368) );
  MUX2X1 U816 ( .B(n1372), .A(n1373), .S(\C2334/net89443 ), .Y(n1371) );
  MUX2X1 U817 ( .B(n1375), .A(n1376), .S(\C2334/net89825 ), .Y(n1374) );
  MUX2X1 U818 ( .B(n1378), .A(n1379), .S(\C2334/net89825 ), .Y(n1377) );
  MUX2X1 U819 ( .B(n1381), .A(n1382), .S(\C2334/net89825 ), .Y(n1380) );
  MUX2X1 U820 ( .B(n1384), .A(n1385), .S(\C2334/net89825 ), .Y(n1383) );
  MUX2X1 U821 ( .B(n1387), .A(n1388), .S(\C2334/net89443 ), .Y(n1386) );
  MUX2X1 U822 ( .B(n1390), .A(n1391), .S(\C2334/net89825 ), .Y(n1389) );
  MUX2X1 U823 ( .B(n1393), .A(n1394), .S(\C2334/net89825 ), .Y(n1392) );
  MUX2X1 U824 ( .B(n1396), .A(n1397), .S(\C2334/net89825 ), .Y(n1395) );
  MUX2X1 U825 ( .B(n1399), .A(n1400), .S(\C2334/net89825 ), .Y(n1398) );
  MUX2X1 U826 ( .B(n1402), .A(n1403), .S(\C2334/net89443 ), .Y(n1401) );
  MUX2X1 U827 ( .B(n1405), .A(n1406), .S(\C2334/net89825 ), .Y(n1404) );
  MUX2X1 U828 ( .B(n1408), .A(n1409), .S(\C2334/net89825 ), .Y(n1407) );
  MUX2X1 U829 ( .B(n1411), .A(n1412), .S(\C2334/net89825 ), .Y(n1410) );
  MUX2X1 U830 ( .B(n1414), .A(n1415), .S(\C2334/net89825 ), .Y(n1413) );
  MUX2X1 U831 ( .B(n1417), .A(n1418), .S(\C2334/net89443 ), .Y(n1416) );
  MUX2X1 U832 ( .B(n1420), .A(n1421), .S(\C2334/net89823 ), .Y(n1419) );
  MUX2X1 U833 ( .B(n1423), .A(n1424), .S(\C2334/net89823 ), .Y(n1422) );
  MUX2X1 U834 ( .B(n1426), .A(n1427), .S(\C2334/net89823 ), .Y(n1425) );
  MUX2X1 U835 ( .B(n1429), .A(n1430), .S(\C2334/net89823 ), .Y(n1428) );
  MUX2X1 U836 ( .B(n1432), .A(n1433), .S(\C2334/net89443 ), .Y(n1431) );
  MUX2X1 U837 ( .B(n1435), .A(n1436), .S(\C2334/net89821 ), .Y(n1434) );
  MUX2X1 U838 ( .B(n1438), .A(n1439), .S(\C2334/net89821 ), .Y(n1437) );
  MUX2X1 U839 ( .B(n1441), .A(n1442), .S(\C2334/net89821 ), .Y(n1440) );
  MUX2X1 U840 ( .B(n1444), .A(n1445), .S(\C2334/net89821 ), .Y(n1443) );
  MUX2X1 U841 ( .B(n1447), .A(n1448), .S(\C2334/net89443 ), .Y(n1446) );
  MUX2X1 U842 ( .B(n1450), .A(n1451), .S(\C2334/net89821 ), .Y(n1449) );
  MUX2X1 U843 ( .B(n1453), .A(n1454), .S(\C2334/net89821 ), .Y(n1452) );
  MUX2X1 U844 ( .B(n1456), .A(n1457), .S(\C2334/net89821 ), .Y(n1455) );
  MUX2X1 U845 ( .B(n1459), .A(n1460), .S(\C2334/net89821 ), .Y(n1458) );
  MUX2X1 U846 ( .B(n1462), .A(n1463), .S(\C2334/net89445 ), .Y(n1461) );
  MUX2X1 U847 ( .B(n1465), .A(n1466), .S(\C2334/net89821 ), .Y(n1464) );
  MUX2X1 U848 ( .B(n1468), .A(n1469), .S(\C2334/net89821 ), .Y(n1467) );
  MUX2X1 U849 ( .B(n1471), .A(n1472), .S(\C2334/net89821 ), .Y(n1470) );
  MUX2X1 U850 ( .B(n1474), .A(n1475), .S(\C2334/net89821 ), .Y(n1473) );
  MUX2X1 U851 ( .B(n1477), .A(n1478), .S(\C2334/net89445 ), .Y(n1476) );
  MUX2X1 U852 ( .B(n1480), .A(n1481), .S(\C2334/net89819 ), .Y(n1479) );
  MUX2X1 U853 ( .B(n1483), .A(n1484), .S(\C2334/net89819 ), .Y(n1482) );
  MUX2X1 U854 ( .B(n1486), .A(n1487), .S(\C2334/net89819 ), .Y(n1485) );
  MUX2X1 U855 ( .B(n1489), .A(n1490), .S(\C2334/net89819 ), .Y(n1488) );
  MUX2X1 U856 ( .B(n1492), .A(n1493), .S(\C2334/net89445 ), .Y(n1491) );
  MUX2X1 U857 ( .B(n1495), .A(n1496), .S(\C2334/net89819 ), .Y(n1494) );
  MUX2X1 U858 ( .B(n1498), .A(n1499), .S(\C2334/net89819 ), .Y(n1497) );
  MUX2X1 U859 ( .B(n1501), .A(n1502), .S(\C2334/net89819 ), .Y(n1500) );
  MUX2X1 U860 ( .B(n1504), .A(n1505), .S(\C2334/net89819 ), .Y(n1503) );
  MUX2X1 U861 ( .B(n1507), .A(n1508), .S(\C2334/net89445 ), .Y(n1506) );
  MUX2X1 U862 ( .B(n1510), .A(n1511), .S(\C2334/net89819 ), .Y(n1509) );
  MUX2X1 U863 ( .B(n1513), .A(n1514), .S(\C2334/net89819 ), .Y(n1512) );
  MUX2X1 U864 ( .B(n1516), .A(n1517), .S(\C2334/net89819 ), .Y(n1515) );
  MUX2X1 U865 ( .B(n1519), .A(n1520), .S(\C2334/net89819 ), .Y(n1518) );
  MUX2X1 U866 ( .B(n1522), .A(n1523), .S(\C2334/net89445 ), .Y(n1521) );
  MUX2X1 U867 ( .B(n1525), .A(n1526), .S(\C2334/net89817 ), .Y(n1524) );
  MUX2X1 U868 ( .B(n1528), .A(n1529), .S(\C2334/net89817 ), .Y(n1527) );
  MUX2X1 U869 ( .B(n1531), .A(n1532), .S(\C2334/net89817 ), .Y(n1530) );
  MUX2X1 U870 ( .B(n1534), .A(n1535), .S(\C2334/net89817 ), .Y(n1533) );
  MUX2X1 U871 ( .B(n1537), .A(n1538), .S(\C2334/net89445 ), .Y(n1536) );
  MUX2X1 U872 ( .B(n1540), .A(n1541), .S(\C2334/net89817 ), .Y(n1539) );
  MUX2X1 U873 ( .B(n1543), .A(n1544), .S(\C2334/net89817 ), .Y(n1542) );
  MUX2X1 U874 ( .B(n1546), .A(n1547), .S(\C2334/net89817 ), .Y(n1545) );
  MUX2X1 U875 ( .B(n1549), .A(n1550), .S(\C2334/net89817 ), .Y(n1548) );
  MUX2X1 U876 ( .B(n1552), .A(n1553), .S(\C2334/net89445 ), .Y(n1551) );
  MUX2X1 U877 ( .B(n1555), .A(n1556), .S(\C2334/net89817 ), .Y(n1554) );
  MUX2X1 U878 ( .B(n1558), .A(n1559), .S(\C2334/net89817 ), .Y(n1557) );
  MUX2X1 U879 ( .B(n1561), .A(n1562), .S(\C2334/net89817 ), .Y(n1560) );
  MUX2X1 U880 ( .B(n1564), .A(n1565), .S(\C2334/net89817 ), .Y(n1563) );
  MUX2X1 U881 ( .B(n1567), .A(n1568), .S(\C2334/net89445 ), .Y(n1566) );
  MUX2X1 U882 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(\C2334/net90389 ), .Y(
        n609) );
  MUX2X1 U883 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(\C2334/net90389 ), .Y(
        n608) );
  MUX2X1 U884 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(\C2334/net90389 ), .Y(
        n612) );
  MUX2X1 U885 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(\C2334/net90389 ), .Y(
        n611) );
  MUX2X1 U886 ( .B(n610), .A(n607), .S(\C2334/net89619 ), .Y(n621) );
  MUX2X1 U887 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(\C2334/net90387 ), .Y(
        n615) );
  MUX2X1 U888 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(\C2334/net90387 ), .Y(
        n614) );
  MUX2X1 U889 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(\C2334/net90387 ), .Y(
        n618) );
  MUX2X1 U890 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(\C2334/net90387 ), .Y(
        n617) );
  MUX2X1 U891 ( .B(n616), .A(n613), .S(\C2334/net89619 ), .Y(n620) );
  MUX2X1 U892 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(\C2334/net90387 ), .Y(
        n624) );
  MUX2X1 U893 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(\C2334/net90387 ), .Y(
        n623) );
  MUX2X1 U894 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(\C2334/net90387 ), .Y(
        n627) );
  MUX2X1 U895 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(\C2334/net90387 ), .Y(
        n626) );
  MUX2X1 U896 ( .B(n625), .A(n622), .S(\C2334/net89619 ), .Y(n636) );
  MUX2X1 U897 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(\C2334/net90387 ), .Y(
        n630) );
  MUX2X1 U898 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(\C2334/net90387 ), .Y(
        n629) );
  MUX2X1 U899 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(\C2334/net90387 ), .Y(
        n633) );
  MUX2X1 U900 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(\C2334/net90387 ), .Y(
        n632) );
  MUX2X1 U901 ( .B(n631), .A(n628), .S(\C2334/net89619 ), .Y(n635) );
  MUX2X1 U902 ( .B(n634), .A(n619), .S(\C2334/net89303 ), .Y(n1569) );
  MUX2X1 U903 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(\C2334/net90385 ), .Y(
        n639) );
  MUX2X1 U904 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(\C2334/net90385 ), .Y(
        n638) );
  MUX2X1 U905 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(\C2334/net90385 ), .Y(
        n642) );
  MUX2X1 U906 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(\C2334/net90385 ), .Y(
        n641) );
  MUX2X1 U907 ( .B(n640), .A(n637), .S(\C2334/net89619 ), .Y(n1163) );
  MUX2X1 U908 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(\C2334/net90385 ), .Y(
        n645) );
  MUX2X1 U909 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(\C2334/net90385 ), .Y(
        n644) );
  MUX2X1 U910 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(\C2334/net90385 ), .Y(
        n648) );
  MUX2X1 U911 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(\C2334/net90385 ), .Y(
        n647) );
  MUX2X1 U912 ( .B(n646), .A(n643), .S(\C2334/net89619 ), .Y(n650) );
  MUX2X1 U913 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(\C2334/net90385 ), .Y(
        n1166) );
  MUX2X1 U914 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(\C2334/net90385 ), .Y(
        n1165) );
  MUX2X1 U915 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(\C2334/net90385 ), .Y(
        n1169) );
  MUX2X1 U916 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(\C2334/net90385 ), .Y(
        n1168) );
  MUX2X1 U917 ( .B(n1167), .A(n1164), .S(\C2334/net89619 ), .Y(n1178) );
  MUX2X1 U918 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(\C2334/net90383 ), .Y(
        n1172) );
  MUX2X1 U919 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(\C2334/net90383 ), .Y(
        n1171) );
  MUX2X1 U920 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(\C2334/net90383 ), .Y(
        n1175) );
  MUX2X1 U921 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(\C2334/net90383 ), .Y(
        n1174) );
  MUX2X1 U922 ( .B(n1173), .A(n1170), .S(\C2334/net89619 ), .Y(n1177) );
  MUX2X1 U923 ( .B(n1176), .A(n649), .S(\C2334/net89303 ), .Y(n1570) );
  MUX2X1 U924 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(\C2334/net90383 ), .Y(
        n1181) );
  MUX2X1 U925 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(\C2334/net90383 ), .Y(
        n1180) );
  MUX2X1 U926 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(\C2334/net90383 ), .Y(
        n1184) );
  MUX2X1 U927 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(\C2334/net90383 ), .Y(
        n1183) );
  MUX2X1 U928 ( .B(n1182), .A(n1179), .S(\C2334/net89619 ), .Y(n1193) );
  MUX2X1 U929 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(\C2334/net90383 ), .Y(
        n1187) );
  MUX2X1 U930 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(\C2334/net90383 ), .Y(
        n1186) );
  MUX2X1 U931 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(\C2334/net90383 ), .Y(
        n1190) );
  MUX2X1 U932 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(\C2334/net90383 ), .Y(
        n1189) );
  MUX2X1 U933 ( .B(n1188), .A(n1185), .S(\C2334/net89619 ), .Y(n1192) );
  MUX2X1 U934 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(\C2334/net90381 ), .Y(
        n1196) );
  MUX2X1 U935 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(\C2334/net90381 ), .Y(
        n1195) );
  MUX2X1 U936 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(\C2334/net90381 ), .Y(
        n1199) );
  MUX2X1 U937 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(\C2334/net90381 ), .Y(
        n1198) );
  MUX2X1 U938 ( .B(n1197), .A(n1194), .S(\C2334/net89619 ), .Y(n1208) );
  MUX2X1 U939 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(\C2334/net90381 ), .Y(
        n1202) );
  MUX2X1 U940 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(\C2334/net90381 ), .Y(
        n1201) );
  MUX2X1 U941 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(\C2334/net90381 ), .Y(
        n1205) );
  MUX2X1 U942 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(\C2334/net90381 ), .Y(
        n1204) );
  MUX2X1 U943 ( .B(n1203), .A(n1200), .S(\C2334/net89619 ), .Y(n1207) );
  MUX2X1 U944 ( .B(n1206), .A(n1191), .S(\C2334/net89303 ), .Y(n1571) );
  MUX2X1 U945 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(\C2334/net90381 ), .Y(
        n1211) );
  MUX2X1 U946 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(\C2334/net90381 ), .Y(
        n1210) );
  MUX2X1 U947 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(\C2334/net90381 ), .Y(
        n1214) );
  MUX2X1 U948 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(\C2334/net90381 ), .Y(
        n1213) );
  MUX2X1 U949 ( .B(n1212), .A(n1209), .S(\C2334/net89621 ), .Y(n1223) );
  MUX2X1 U950 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(\C2334/net90377 ), .Y(
        n1217) );
  MUX2X1 U951 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(\C2334/net90389 ), .Y(
        n1216) );
  MUX2X1 U952 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(\C2334/net90377 ), .Y(
        n1220) );
  MUX2X1 U953 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(\C2334/net90375 ), .Y(
        n1219) );
  MUX2X1 U954 ( .B(n1218), .A(n1215), .S(\C2334/net89621 ), .Y(n1222) );
  MUX2X1 U955 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(\C2334/net90355 ), .Y(
        n1226) );
  MUX2X1 U956 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(\C2334/net90377 ), .Y(
        n1225) );
  MUX2X1 U957 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(\C2334/net90389 ), .Y(
        n1229) );
  MUX2X1 U958 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(\C2334/net90389 ), .Y(
        n1228) );
  MUX2X1 U959 ( .B(n1227), .A(n1224), .S(\C2334/net89621 ), .Y(n1238) );
  MUX2X1 U960 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(\C2334/net90355 ), .Y(
        n1232) );
  MUX2X1 U961 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(\C2334/net90355 ), .Y(
        n1231) );
  MUX2X1 U962 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(\C2334/net90389 ), .Y(
        n1235) );
  MUX2X1 U963 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(\C2334/net90371 ), .Y(
        n1234) );
  MUX2X1 U964 ( .B(n1233), .A(n1230), .S(\C2334/net89621 ), .Y(n1237) );
  MUX2X1 U965 ( .B(n1236), .A(n1221), .S(\C2334/net89303 ), .Y(n1572) );
  MUX2X1 U966 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(\C2334/net90377 ), .Y(
        n1241) );
  MUX2X1 U967 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(\C2334/net90377 ), .Y(
        n1240) );
  MUX2X1 U968 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(\C2334/net90377 ), .Y(
        n1244) );
  MUX2X1 U969 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(\C2334/net90377 ), .Y(
        n1243) );
  MUX2X1 U970 ( .B(n1242), .A(n1239), .S(\C2334/net89621 ), .Y(n1253) );
  MUX2X1 U971 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(\C2334/net90377 ), .Y(
        n1247) );
  MUX2X1 U972 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(\C2334/net90377 ), .Y(
        n1246) );
  MUX2X1 U973 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(\C2334/net90377 ), .Y(
        n1250) );
  MUX2X1 U974 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(\C2334/net90377 ), .Y(
        n1249) );
  MUX2X1 U975 ( .B(n1248), .A(n1245), .S(\C2334/net89621 ), .Y(n1252) );
  MUX2X1 U976 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(\C2334/net90377 ), .Y(
        n1256) );
  MUX2X1 U977 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(\C2334/net90377 ), .Y(
        n1255) );
  MUX2X1 U978 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(\C2334/net90377 ), .Y(
        n1259) );
  MUX2X1 U979 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(\C2334/net90377 ), .Y(
        n1258) );
  MUX2X1 U980 ( .B(n1257), .A(n1254), .S(\C2334/net89621 ), .Y(n1268) );
  MUX2X1 U981 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(\C2334/net90375 ), .Y(
        n1262) );
  MUX2X1 U982 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(\C2334/net90375 ), .Y(
        n1261) );
  MUX2X1 U983 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(\C2334/net90375 ), .Y(
        n1265) );
  MUX2X1 U984 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(\C2334/net90375 ), .Y(
        n1264) );
  MUX2X1 U985 ( .B(n1263), .A(n1260), .S(\C2334/net89621 ), .Y(n1267) );
  MUX2X1 U986 ( .B(n1266), .A(n1251), .S(\C2334/net89303 ), .Y(n1573) );
  MUX2X1 U987 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(\C2334/net90375 ), .Y(
        n1271) );
  MUX2X1 U988 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(\C2334/net90375 ), .Y(
        n1270) );
  MUX2X1 U989 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(\C2334/net90375 ), .Y(
        n1274) );
  MUX2X1 U990 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(\C2334/net90375 ), .Y(
        n1273) );
  MUX2X1 U991 ( .B(n1272), .A(n1269), .S(\C2334/net89621 ), .Y(n1283) );
  MUX2X1 U992 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(\C2334/net90375 ), .Y(
        n1277) );
  MUX2X1 U993 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(\C2334/net90375 ), .Y(
        n1276) );
  MUX2X1 U994 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(\C2334/net90375 ), .Y(
        n1280) );
  MUX2X1 U995 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(\C2334/net90375 ), .Y(
        n1279) );
  MUX2X1 U996 ( .B(n1278), .A(n1275), .S(\C2334/net89621 ), .Y(n1282) );
  MUX2X1 U997 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(\C2334/net90373 ), .Y(
        n1286) );
  MUX2X1 U998 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(\C2334/net90373 ), .Y(
        n1285) );
  MUX2X1 U999 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(\C2334/net90373 ), .Y(
        n1289) );
  MUX2X1 U1000 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(\C2334/net90373 ), .Y(
        n1288) );
  MUX2X1 U1001 ( .B(n1287), .A(n1284), .S(\C2334/net89621 ), .Y(n1298) );
  MUX2X1 U1002 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(\C2334/net90373 ), .Y(
        n1292) );
  MUX2X1 U1003 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(\C2334/net90373 ), .Y(
        n1291) );
  MUX2X1 U1004 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(\C2334/net90373 ), .Y(
        n1295) );
  MUX2X1 U1005 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(\C2334/net90373 ), .Y(
        n1294) );
  MUX2X1 U1006 ( .B(n1293), .A(n1290), .S(\C2334/net89621 ), .Y(n1297) );
  MUX2X1 U1007 ( .B(n1296), .A(n1281), .S(\C2334/net89303 ), .Y(n1574) );
  MUX2X1 U1008 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(\C2334/net90373 ), .Y(
        n1301) );
  MUX2X1 U1009 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(\C2334/net90373 ), .Y(
        n1300) );
  MUX2X1 U1010 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(\C2334/net90373 ), .Y(
        n1304) );
  MUX2X1 U1011 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(\C2334/net90373 ), .Y(
        n1303) );
  MUX2X1 U1012 ( .B(n1302), .A(n1299), .S(\C2334/net89623 ), .Y(n1313) );
  MUX2X1 U1013 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(\C2334/net90371 ), .Y(
        n1307) );
  MUX2X1 U1014 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(\C2334/net90371 ), .Y(
        n1306) );
  MUX2X1 U1015 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(\C2334/net90371 ), .Y(
        n1310) );
  MUX2X1 U1016 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(\C2334/net90371 ), .Y(
        n1309) );
  MUX2X1 U1017 ( .B(n1308), .A(n1305), .S(\C2334/net89623 ), .Y(n1312) );
  MUX2X1 U1018 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(\C2334/net90371 ), .Y(
        n1316) );
  MUX2X1 U1019 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(\C2334/net90371 ), .Y(
        n1315) );
  MUX2X1 U1020 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(\C2334/net90371 ), .Y(
        n1319) );
  MUX2X1 U1021 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(\C2334/net90371 ), .Y(
        n1318) );
  MUX2X1 U1022 ( .B(n1317), .A(n1314), .S(\C2334/net89623 ), .Y(n1328) );
  MUX2X1 U1023 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(\C2334/net90371 ), .Y(
        n1322) );
  MUX2X1 U1024 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(\C2334/net90371 ), .Y(
        n1321) );
  MUX2X1 U1025 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(\C2334/net90371 ), .Y(
        n1325) );
  MUX2X1 U1026 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(\C2334/net90371 ), .Y(
        n1324) );
  MUX2X1 U1027 ( .B(n1323), .A(n1320), .S(\C2334/net89623 ), .Y(n1327) );
  MUX2X1 U1028 ( .B(n1326), .A(n1311), .S(\C2334/net89303 ), .Y(n1575) );
  MUX2X1 U1029 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(\C2334/net90369 ), .Y(
        n1331) );
  MUX2X1 U1030 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(\C2334/net90369 ), .Y(
        n1330) );
  MUX2X1 U1031 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(\C2334/net90369 ), .Y(
        n1334) );
  MUX2X1 U1032 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(\C2334/net90369 ), .Y(
        n1333) );
  MUX2X1 U1033 ( .B(n1332), .A(n1329), .S(\C2334/net89623 ), .Y(n1343) );
  MUX2X1 U1034 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(\C2334/net90369 ), .Y(
        n1337) );
  MUX2X1 U1035 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(\C2334/net90369 ), .Y(
        n1336) );
  MUX2X1 U1036 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(\C2334/net90369 ), .Y(
        n1340) );
  MUX2X1 U1037 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(\C2334/net90369 ), .Y(
        n1339) );
  MUX2X1 U1038 ( .B(n1338), .A(n1335), .S(\C2334/net89623 ), .Y(n1342) );
  MUX2X1 U1039 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(\C2334/net90369 ), .Y(
        n1346) );
  MUX2X1 U1040 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(\C2334/net90369 ), .Y(
        n1345) );
  MUX2X1 U1041 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(\C2334/net90369 ), .Y(
        n1349) );
  MUX2X1 U1042 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(\C2334/net90369 ), .Y(
        n1348) );
  MUX2X1 U1043 ( .B(n1347), .A(n1344), .S(\C2334/net89623 ), .Y(n1358) );
  MUX2X1 U1044 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(\C2334/net90367 ), .Y(
        n1352) );
  MUX2X1 U1045 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(\C2334/net90367 ), .Y(
        n1351) );
  MUX2X1 U1046 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(\C2334/net90367 ), .Y(
        n1355) );
  MUX2X1 U1047 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(\C2334/net90367 ), .Y(
        n1354) );
  MUX2X1 U1048 ( .B(n1353), .A(n1350), .S(\C2334/net89623 ), .Y(n1357) );
  MUX2X1 U1049 ( .B(n1356), .A(n1341), .S(\C2334/net89303 ), .Y(n1576) );
  MUX2X1 U1050 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(\C2334/net90367 ), .Y(
        n1361) );
  MUX2X1 U1051 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(\C2334/net90367 ), .Y(
        n1360) );
  MUX2X1 U1052 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(\C2334/net90367 ), .Y(
        n1364) );
  MUX2X1 U1053 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(\C2334/net90367 ), .Y(
        n1363) );
  MUX2X1 U1054 ( .B(n1362), .A(n1359), .S(\C2334/net89623 ), .Y(n1373) );
  MUX2X1 U1055 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(\C2334/net90367 ), .Y(
        n1367) );
  MUX2X1 U1056 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(\C2334/net90367 ), .Y(
        n1366) );
  MUX2X1 U1057 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(\C2334/net90367 ), .Y(
        n1370) );
  MUX2X1 U1058 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(\C2334/net90367 ), .Y(
        n1369) );
  MUX2X1 U1059 ( .B(n1368), .A(n1365), .S(\C2334/net89623 ), .Y(n1372) );
  MUX2X1 U1060 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(\C2334/net90365 ), .Y(
        n1376) );
  MUX2X1 U1061 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(\C2334/net90365 ), .Y(
        n1375) );
  MUX2X1 U1062 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(\C2334/net90365 ), .Y(
        n1379) );
  MUX2X1 U1063 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(\C2334/net90365 ), .Y(
        n1378) );
  MUX2X1 U1064 ( .B(n1377), .A(n1374), .S(\C2334/net89623 ), .Y(n1388) );
  MUX2X1 U1065 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(\C2334/net90365 ), .Y(
        n1382) );
  MUX2X1 U1066 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(\C2334/net90365 ), .Y(
        n1381) );
  MUX2X1 U1067 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(\C2334/net90365 ), .Y(
        n1385) );
  MUX2X1 U1068 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(\C2334/net90365 ), .Y(
        n1384) );
  MUX2X1 U1069 ( .B(n1383), .A(n1380), .S(\C2334/net89623 ), .Y(n1387) );
  MUX2X1 U1070 ( .B(n1386), .A(n1371), .S(\C2334/net89303 ), .Y(n1577) );
  MUX2X1 U1071 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(\C2334/net90365 ), .Y(
        n1391) );
  MUX2X1 U1072 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(\C2334/net90365 ), .Y(
        n1390) );
  MUX2X1 U1073 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(\C2334/net90365 ), .Y(
        n1394) );
  MUX2X1 U1074 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(\C2334/net90365 ), .Y(
        n1393) );
  MUX2X1 U1075 ( .B(n1392), .A(n1389), .S(\C2334/net89625 ), .Y(n1403) );
  MUX2X1 U1076 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(\C2334/net90363 ), .Y(
        n1397) );
  MUX2X1 U1077 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(\C2334/net90363 ), .Y(
        n1396) );
  MUX2X1 U1078 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(\C2334/net90363 ), .Y(
        n1400) );
  MUX2X1 U1079 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(\C2334/net90363 ), .Y(
        n1399) );
  MUX2X1 U1080 ( .B(n1398), .A(n1395), .S(\C2334/net89625 ), .Y(n1402) );
  MUX2X1 U1081 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(\C2334/net90363 ), .Y(
        n1406) );
  MUX2X1 U1082 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(\C2334/net90363 ), .Y(
        n1405) );
  MUX2X1 U1083 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(\C2334/net90363 ), .Y(
        n1409) );
  MUX2X1 U1084 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(\C2334/net90363 ), .Y(
        n1408) );
  MUX2X1 U1085 ( .B(n1407), .A(n1404), .S(\C2334/net89625 ), .Y(n1418) );
  MUX2X1 U1086 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(\C2334/net90363 ), .Y(
        n1412) );
  MUX2X1 U1087 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(\C2334/net90363 ), .Y(
        n1411) );
  MUX2X1 U1088 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(\C2334/net90363 ), .Y(
        n1415) );
  MUX2X1 U1089 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(\C2334/net90363 ), .Y(
        n1414) );
  MUX2X1 U1090 ( .B(n1413), .A(n1410), .S(\C2334/net89625 ), .Y(n1417) );
  MUX2X1 U1091 ( .B(n1416), .A(n1401), .S(\C2334/net89303 ), .Y(n1578) );
  MUX2X1 U1092 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(\C2334/net90359 ), 
        .Y(n1421) );
  MUX2X1 U1093 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(\C2334/net90359 ), 
        .Y(n1420) );
  MUX2X1 U1094 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(\C2334/net90359 ), 
        .Y(n1424) );
  MUX2X1 U1095 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(\C2334/net90359 ), 
        .Y(n1423) );
  MUX2X1 U1096 ( .B(n1422), .A(n1419), .S(\C2334/net89625 ), .Y(n1433) );
  MUX2X1 U1097 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(\C2334/net90359 ), 
        .Y(n1427) );
  MUX2X1 U1098 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(\C2334/net90359 ), 
        .Y(n1426) );
  MUX2X1 U1099 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(\C2334/net90359 ), 
        .Y(n1430) );
  MUX2X1 U1100 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(\C2334/net90359 ), 
        .Y(n1429) );
  MUX2X1 U1101 ( .B(n1428), .A(n1425), .S(\C2334/net89625 ), .Y(n1432) );
  MUX2X1 U1102 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(\C2334/net90357 ), 
        .Y(n1436) );
  MUX2X1 U1103 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(\C2334/net90357 ), 
        .Y(n1435) );
  MUX2X1 U1104 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(\C2334/net90357 ), 
        .Y(n1439) );
  MUX2X1 U1105 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(\C2334/net90357 ), .Y(
        n1438) );
  MUX2X1 U1106 ( .B(n1437), .A(n1434), .S(\C2334/net89625 ), .Y(n1448) );
  MUX2X1 U1107 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(\C2334/net90357 ), .Y(
        n1442) );
  MUX2X1 U1108 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(\C2334/net90357 ), .Y(
        n1441) );
  MUX2X1 U1109 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(\C2334/net90357 ), .Y(
        n1445) );
  MUX2X1 U1110 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(\C2334/net90357 ), .Y(
        n1444) );
  MUX2X1 U1111 ( .B(n1443), .A(n1440), .S(\C2334/net89625 ), .Y(n1447) );
  MUX2X1 U1112 ( .B(n1446), .A(n1431), .S(\C2334/net89303 ), .Y(n1579) );
  MUX2X1 U1113 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(\C2334/net90357 ), 
        .Y(n1451) );
  MUX2X1 U1114 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(\C2334/net90357 ), 
        .Y(n1450) );
  MUX2X1 U1115 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(\C2334/net90357 ), 
        .Y(n1454) );
  MUX2X1 U1116 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(\C2334/net90357 ), 
        .Y(n1453) );
  MUX2X1 U1117 ( .B(n1452), .A(n1449), .S(\C2334/net89627 ), .Y(n1463) );
  MUX2X1 U1118 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(\C2334/net90355 ), 
        .Y(n1457) );
  MUX2X1 U1119 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(\C2334/net90355 ), 
        .Y(n1456) );
  MUX2X1 U1120 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(\C2334/net90355 ), 
        .Y(n1460) );
  MUX2X1 U1121 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(\C2334/net90355 ), 
        .Y(n1459) );
  MUX2X1 U1122 ( .B(n1458), .A(n1455), .S(\C2334/net89627 ), .Y(n1462) );
  MUX2X1 U1123 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(\C2334/net90355 ), 
        .Y(n1466) );
  MUX2X1 U1124 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(\C2334/net90355 ), 
        .Y(n1465) );
  MUX2X1 U1125 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(\C2334/net90355 ), 
        .Y(n1469) );
  MUX2X1 U1126 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(\C2334/net90355 ), .Y(
        n1468) );
  MUX2X1 U1127 ( .B(n1467), .A(n1464), .S(\C2334/net89627 ), .Y(n1478) );
  MUX2X1 U1128 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(\C2334/net90355 ), .Y(
        n1472) );
  MUX2X1 U1129 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(\C2334/net90355 ), .Y(
        n1471) );
  MUX2X1 U1130 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(\C2334/net90355 ), .Y(
        n1475) );
  MUX2X1 U1131 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(\C2334/net90355 ), .Y(
        n1474) );
  MUX2X1 U1132 ( .B(n1473), .A(n1470), .S(\C2334/net89627 ), .Y(n1477) );
  MUX2X1 U1133 ( .B(n1476), .A(n1461), .S(\C2334/net89305 ), .Y(n1580) );
  MUX2X1 U1134 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(\C2334/net90353 ), 
        .Y(n1481) );
  MUX2X1 U1135 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(\C2334/net90353 ), 
        .Y(n1480) );
  MUX2X1 U1136 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(\C2334/net90353 ), 
        .Y(n1484) );
  MUX2X1 U1137 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(\C2334/net90353 ), 
        .Y(n1483) );
  MUX2X1 U1138 ( .B(n1482), .A(n1479), .S(\C2334/net89627 ), .Y(n1493) );
  MUX2X1 U1139 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(\C2334/net90353 ), 
        .Y(n1487) );
  MUX2X1 U1140 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(\C2334/net90353 ), 
        .Y(n1486) );
  MUX2X1 U1141 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(\C2334/net90353 ), 
        .Y(n1490) );
  MUX2X1 U1142 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(\C2334/net90353 ), 
        .Y(n1489) );
  MUX2X1 U1143 ( .B(n1488), .A(n1485), .S(\C2334/net89627 ), .Y(n1492) );
  MUX2X1 U1144 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(\C2334/net90353 ), 
        .Y(n1496) );
  MUX2X1 U1145 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(\C2334/net90353 ), 
        .Y(n1495) );
  MUX2X1 U1146 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(\C2334/net90353 ), 
        .Y(n1499) );
  MUX2X1 U1147 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(\C2334/net90353 ), .Y(
        n1498) );
  MUX2X1 U1148 ( .B(n1497), .A(n1494), .S(\C2334/net89627 ), .Y(n1508) );
  MUX2X1 U1149 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(\C2334/net90351 ), .Y(
        n1502) );
  MUX2X1 U1150 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(\C2334/net90351 ), .Y(
        n1501) );
  MUX2X1 U1151 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(\C2334/net90351 ), .Y(
        n1505) );
  MUX2X1 U1152 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(\C2334/net90351 ), .Y(
        n1504) );
  MUX2X1 U1153 ( .B(n1503), .A(n1500), .S(\C2334/net89627 ), .Y(n1507) );
  MUX2X1 U1154 ( .B(n1506), .A(n1491), .S(\C2334/net89305 ), .Y(n1581) );
  MUX2X1 U1155 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(\C2334/net90351 ), 
        .Y(n1511) );
  MUX2X1 U1156 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(\C2334/net90351 ), 
        .Y(n1510) );
  MUX2X1 U1157 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(\C2334/net90351 ), 
        .Y(n1514) );
  MUX2X1 U1158 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(\C2334/net90351 ), 
        .Y(n1513) );
  MUX2X1 U1159 ( .B(n1512), .A(n1509), .S(\C2334/net89627 ), .Y(n1523) );
  MUX2X1 U1160 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(\C2334/net90351 ), 
        .Y(n1517) );
  MUX2X1 U1161 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(\C2334/net90351 ), 
        .Y(n1516) );
  MUX2X1 U1162 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(\C2334/net90351 ), 
        .Y(n1520) );
  MUX2X1 U1163 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(\C2334/net90351 ), 
        .Y(n1519) );
  MUX2X1 U1164 ( .B(n1518), .A(n1515), .S(\C2334/net89627 ), .Y(n1522) );
  MUX2X1 U1165 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(\C2334/net90349 ), 
        .Y(n1526) );
  MUX2X1 U1166 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(\C2334/net90349 ), 
        .Y(n1525) );
  MUX2X1 U1167 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(\C2334/net90349 ), 
        .Y(n1529) );
  MUX2X1 U1168 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(\C2334/net90349 ), .Y(
        n1528) );
  MUX2X1 U1169 ( .B(n1527), .A(n1524), .S(\C2334/net89627 ), .Y(n1538) );
  MUX2X1 U1170 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(\C2334/net90349 ), .Y(
        n1532) );
  MUX2X1 U1171 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(\C2334/net90349 ), .Y(
        n1531) );
  MUX2X1 U1172 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(\C2334/net90349 ), .Y(
        n1535) );
  MUX2X1 U1173 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(\C2334/net90349 ), .Y(
        n1534) );
  MUX2X1 U1174 ( .B(n1533), .A(n1530), .S(\C2334/net89627 ), .Y(n1537) );
  MUX2X1 U1175 ( .B(n1536), .A(n1521), .S(\C2334/net89305 ), .Y(n1582) );
  MUX2X1 U1177 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(\C2334/net90349 ), 
        .Y(n1541) );
  MUX2X1 U1178 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(\C2334/net90349 ), 
        .Y(n1540) );
  MUX2X1 U1179 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(\C2334/net90349 ), 
        .Y(n1544) );
  MUX2X1 U1180 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(\C2334/net90349 ), 
        .Y(n1543) );
  MUX2X1 U1181 ( .B(n1542), .A(n1539), .S(\C2334/net89629 ), .Y(n1553) );
  MUX2X1 U1182 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(\C2334/net90347 ), 
        .Y(n1547) );
  MUX2X1 U1183 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(\C2334/net90347 ), 
        .Y(n1546) );
  MUX2X1 U1184 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(\C2334/net90347 ), 
        .Y(n1550) );
  MUX2X1 U1185 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(\C2334/net90347 ), 
        .Y(n1549) );
  MUX2X1 U1186 ( .B(n1548), .A(n1545), .S(\C2334/net89629 ), .Y(n1552) );
  MUX2X1 U1187 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(\C2334/net90347 ), 
        .Y(n1556) );
  MUX2X1 U1188 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(\C2334/net90347 ), 
        .Y(n1555) );
  MUX2X1 U1189 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(\C2334/net90347 ), 
        .Y(n1559) );
  MUX2X1 U1190 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(\C2334/net90347 ), .Y(
        n1558) );
  MUX2X1 U1191 ( .B(n1557), .A(n1554), .S(\C2334/net89629 ), .Y(n1568) );
  MUX2X1 U1192 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(\C2334/net90347 ), .Y(
        n1562) );
  MUX2X1 U1193 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(\C2334/net90347 ), .Y(
        n1561) );
  MUX2X1 U1194 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(\C2334/net90347 ), .Y(
        n1565) );
  MUX2X1 U1195 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(\C2334/net90347 ), .Y(
        n1564) );
  MUX2X1 U1196 ( .B(n1563), .A(n1560), .S(\C2334/net89629 ), .Y(n1567) );
  MUX2X1 U1197 ( .B(n1566), .A(n1551), .S(\C2334/net89305 ), .Y(n1583) );
  INVX8 U1198 ( .A(\C2334/net90085 ), .Y(\C2334/net89841 ) );
  INVX8 U1199 ( .A(\C2334/net89839 ), .Y(\C2334/net89837 ) );
  INVX8 U1200 ( .A(\C2334/net89839 ), .Y(\C2334/net89835 ) );
  INVX8 U1201 ( .A(\C2334/net89839 ), .Y(\C2334/net89833 ) );
  INVX8 U1202 ( .A(\C2334/net90829 ), .Y(\C2334/net90405 ) );
  INVX8 U1203 ( .A(\C2334/net90829 ), .Y(\C2334/net90401 ) );
  INVX8 U1204 ( .A(\C2334/net90829 ), .Y(\C2334/net90399 ) );
  INVX8 U1205 ( .A(\C2334/net90829 ), .Y(\C2334/net90397 ) );
  INVX8 U1206 ( .A(\C2334/net90829 ), .Y(\C2334/net90393 ) );
  INVX8 U1207 ( .A(\C2334/net90829 ), .Y(\C2334/net90391 ) );
  INVX8 U1208 ( .A(\C2334/net90391 ), .Y(\C2334/net90389 ) );
  INVX8 U1209 ( .A(\C2334/net90391 ), .Y(\C2334/net90387 ) );
  INVX8 U1210 ( .A(\C2334/net90391 ), .Y(\C2334/net90385 ) );
  INVX8 U1211 ( .A(\C2334/net90393 ), .Y(\C2334/net90383 ) );
  INVX8 U1212 ( .A(\C2334/net90393 ), .Y(\C2334/net90381 ) );
  INVX8 U1213 ( .A(\C2334/net90393 ), .Y(\C2334/net90377 ) );
  INVX8 U1214 ( .A(\C2334/net90393 ), .Y(\C2334/net90375 ) );
  INVX8 U1215 ( .A(\C2334/net90391 ), .Y(\C2334/net90373 ) );
  INVX8 U1216 ( .A(\C2334/net90397 ), .Y(\C2334/net90371 ) );
  INVX8 U1217 ( .A(\C2334/net90397 ), .Y(\C2334/net90369 ) );
  INVX8 U1218 ( .A(\C2334/net90397 ), .Y(\C2334/net90367 ) );
  INVX8 U1219 ( .A(\C2334/net90399 ), .Y(\C2334/net90365 ) );
  INVX8 U1220 ( .A(\C2334/net90399 ), .Y(\C2334/net90363 ) );
  INVX8 U1221 ( .A(\C2334/net90401 ), .Y(\C2334/net90357 ) );
  INVX8 U1222 ( .A(\C2334/net90401 ), .Y(\C2334/net90355 ) );
  INVX8 U1223 ( .A(\C2334/net90405 ), .Y(\C2334/net90353 ) );
  INVX8 U1224 ( .A(\C2334/net90405 ), .Y(\C2334/net90351 ) );
  INVX8 U1225 ( .A(\C2334/net90405 ), .Y(\C2334/net90349 ) );
  INVX8 U1226 ( .A(\C2334/net90405 ), .Y(\C2334/net90347 ) );
  INVX8 U1227 ( .A(\C2334/net90835 ), .Y(\C2334/net90829 ) );
  INVX1 U1228 ( .A(N10), .Y(net90763) );
  AND2X2 U1229 ( .A(net130272), .B(net90943), .Y(n1584) );
  INVX8 U1230 ( .A(n409), .Y(n1648) );
  INVX8 U1231 ( .A(n409), .Y(n1649) );
  INVX8 U1232 ( .A(n410), .Y(n1650) );
  INVX8 U1233 ( .A(n410), .Y(n1651) );
  INVX8 U1234 ( .A(n411), .Y(n1652) );
  INVX8 U1235 ( .A(n411), .Y(n1653) );
  INVX8 U1236 ( .A(n412), .Y(n1654) );
  INVX8 U1237 ( .A(n412), .Y(n1655) );
  INVX8 U1238 ( .A(n413), .Y(n1656) );
  INVX8 U1239 ( .A(n413), .Y(n1657) );
  INVX8 U1240 ( .A(n414), .Y(n1658) );
  INVX8 U1241 ( .A(n414), .Y(n1659) );
  INVX8 U1242 ( .A(n415), .Y(n1660) );
  INVX8 U1243 ( .A(n415), .Y(n1661) );
  INVX8 U1244 ( .A(n416), .Y(n1662) );
  INVX8 U1245 ( .A(n416), .Y(n1663) );
  INVX8 U1246 ( .A(n417), .Y(n1664) );
  INVX8 U1247 ( .A(n417), .Y(n1665) );
  INVX8 U1248 ( .A(n418), .Y(n1666) );
  INVX8 U1249 ( .A(n418), .Y(n1667) );
  INVX8 U1250 ( .A(n419), .Y(n1668) );
  INVX8 U1251 ( .A(n419), .Y(n1669) );
  INVX8 U1252 ( .A(n420), .Y(n1671) );
  INVX8 U1253 ( .A(n421), .Y(n1673) );
  INVX8 U1254 ( .A(n422), .Y(n1675) );
  INVX8 U1255 ( .A(n423), .Y(n1677) );
  INVX8 U1256 ( .A(n6), .Y(n1679) );
  NAND2X1 U1257 ( .A(\mem<31><0> ), .B(n390), .Y(n1680) );
  OAI21X1 U1258 ( .A(n1586), .B(n1648), .C(n1680), .Y(n2563) );
  NAND2X1 U1259 ( .A(\mem<31><1> ), .B(n390), .Y(n1681) );
  OAI21X1 U1260 ( .A(n1651), .B(n1585), .C(n1681), .Y(n2562) );
  NAND2X1 U1261 ( .A(\mem<31><2> ), .B(n390), .Y(n1682) );
  OAI21X1 U1262 ( .A(n1653), .B(n1585), .C(n1682), .Y(n2561) );
  NAND2X1 U1263 ( .A(\mem<31><3> ), .B(n390), .Y(n1683) );
  OAI21X1 U1264 ( .A(n1655), .B(n1585), .C(n1683), .Y(n2560) );
  NAND2X1 U1265 ( .A(\mem<31><4> ), .B(n390), .Y(n1684) );
  OAI21X1 U1266 ( .A(n1657), .B(n1585), .C(n1684), .Y(n2559) );
  NAND2X1 U1267 ( .A(\mem<31><5> ), .B(n390), .Y(n1685) );
  OAI21X1 U1268 ( .A(n1659), .B(n1585), .C(n1685), .Y(n2558) );
  NAND2X1 U1269 ( .A(\mem<31><6> ), .B(n390), .Y(n1686) );
  OAI21X1 U1270 ( .A(n1661), .B(n1585), .C(n1686), .Y(n2557) );
  NAND2X1 U1271 ( .A(\mem<31><7> ), .B(n390), .Y(n1687) );
  OAI21X1 U1272 ( .A(n1663), .B(n1585), .C(n1687), .Y(n2556) );
  NAND2X1 U1273 ( .A(\mem<31><8> ), .B(n390), .Y(n1688) );
  OAI21X1 U1274 ( .A(n1665), .B(n1585), .C(n1688), .Y(n2555) );
  NAND2X1 U1275 ( .A(\mem<31><9> ), .B(n390), .Y(n1689) );
  OAI21X1 U1276 ( .A(n1667), .B(n1586), .C(n1689), .Y(n2554) );
  NAND2X1 U1277 ( .A(\mem<31><10> ), .B(n390), .Y(n1690) );
  OAI21X1 U1278 ( .A(n1669), .B(n1586), .C(n1690), .Y(n2553) );
  NAND2X1 U1279 ( .A(\mem<31><11> ), .B(n390), .Y(n1691) );
  OAI21X1 U1280 ( .A(n1671), .B(n1586), .C(n1691), .Y(n2552) );
  NAND2X1 U1281 ( .A(\mem<31><12> ), .B(n390), .Y(n1692) );
  OAI21X1 U1282 ( .A(n1673), .B(n1586), .C(n1692), .Y(n2551) );
  NAND2X1 U1283 ( .A(\mem<31><13> ), .B(n390), .Y(n1693) );
  OAI21X1 U1284 ( .A(n1675), .B(n1586), .C(n1693), .Y(n2550) );
  NAND2X1 U1285 ( .A(\mem<31><14> ), .B(n390), .Y(n1694) );
  OAI21X1 U1286 ( .A(n1677), .B(n1586), .C(n1694), .Y(n2549) );
  NAND2X1 U1287 ( .A(\mem<31><15> ), .B(n390), .Y(n1695) );
  OAI21X1 U1288 ( .A(n1679), .B(n1586), .C(n1695), .Y(n2548) );
  NAND2X1 U1289 ( .A(\mem<30><0> ), .B(n392), .Y(n1696) );
  OAI21X1 U1290 ( .A(n1587), .B(n1648), .C(n1696), .Y(n2547) );
  NAND2X1 U1291 ( .A(\mem<30><1> ), .B(n392), .Y(n1697) );
  OAI21X1 U1292 ( .A(n1587), .B(n1651), .C(n1697), .Y(n2546) );
  NAND2X1 U1293 ( .A(\mem<30><2> ), .B(n392), .Y(n1698) );
  OAI21X1 U1294 ( .A(n1587), .B(n1653), .C(n1698), .Y(n2545) );
  NAND2X1 U1295 ( .A(\mem<30><3> ), .B(n392), .Y(n1699) );
  OAI21X1 U1296 ( .A(n1587), .B(n1655), .C(n1699), .Y(n2544) );
  NAND2X1 U1297 ( .A(\mem<30><4> ), .B(n392), .Y(n1700) );
  OAI21X1 U1298 ( .A(n1587), .B(n1657), .C(n1700), .Y(n2543) );
  NAND2X1 U1299 ( .A(\mem<30><5> ), .B(n392), .Y(n1701) );
  OAI21X1 U1300 ( .A(n1587), .B(n1659), .C(n1701), .Y(n2542) );
  NAND2X1 U1301 ( .A(\mem<30><6> ), .B(n392), .Y(n1702) );
  OAI21X1 U1302 ( .A(n1587), .B(n1661), .C(n1702), .Y(n2541) );
  NAND2X1 U1303 ( .A(\mem<30><7> ), .B(n392), .Y(n1703) );
  OAI21X1 U1304 ( .A(n1587), .B(n1663), .C(n1703), .Y(n2540) );
  NAND2X1 U1305 ( .A(\mem<30><8> ), .B(n392), .Y(n1704) );
  OAI21X1 U1306 ( .A(n1588), .B(n1664), .C(n1704), .Y(n2539) );
  NAND2X1 U1307 ( .A(\mem<30><9> ), .B(n392), .Y(n1705) );
  OAI21X1 U1308 ( .A(n1588), .B(n1666), .C(n1705), .Y(n2538) );
  NAND2X1 U1309 ( .A(\mem<30><10> ), .B(n392), .Y(n1706) );
  OAI21X1 U1310 ( .A(n1588), .B(n1668), .C(n1706), .Y(n2537) );
  NAND2X1 U1311 ( .A(\mem<30><11> ), .B(n392), .Y(n1707) );
  OAI21X1 U1312 ( .A(n1588), .B(n1671), .C(n1707), .Y(n2536) );
  NAND2X1 U1313 ( .A(\mem<30><12> ), .B(n392), .Y(n1708) );
  OAI21X1 U1314 ( .A(n1588), .B(n1673), .C(n1708), .Y(n2535) );
  NAND2X1 U1315 ( .A(\mem<30><13> ), .B(n392), .Y(n1709) );
  OAI21X1 U1316 ( .A(n1588), .B(n1675), .C(n1709), .Y(n2534) );
  NAND2X1 U1317 ( .A(\mem<30><14> ), .B(n392), .Y(n1710) );
  OAI21X1 U1318 ( .A(n1588), .B(n1677), .C(n1710), .Y(n2533) );
  NAND2X1 U1319 ( .A(\mem<30><15> ), .B(n392), .Y(n1711) );
  OAI21X1 U1320 ( .A(n1588), .B(n1678), .C(n1711), .Y(n2532) );
  NAND3X1 U1321 ( .A(net90761), .B(\C2334/net89629 ), .C(net90019), .Y(n1712)
         );
  NAND2X1 U1322 ( .A(\mem<29><0> ), .B(n394), .Y(n1713) );
  OAI21X1 U1323 ( .A(n1589), .B(n1648), .C(n1713), .Y(n2531) );
  NAND2X1 U1324 ( .A(\mem<29><1> ), .B(n394), .Y(n1714) );
  OAI21X1 U1325 ( .A(n1589), .B(n1650), .C(n1714), .Y(n2530) );
  NAND2X1 U1326 ( .A(\mem<29><2> ), .B(n394), .Y(n1715) );
  OAI21X1 U1327 ( .A(n1589), .B(n1652), .C(n1715), .Y(n2529) );
  NAND2X1 U1328 ( .A(\mem<29><3> ), .B(n394), .Y(n1716) );
  OAI21X1 U1329 ( .A(n1589), .B(n1654), .C(n1716), .Y(n2528) );
  NAND2X1 U1330 ( .A(\mem<29><4> ), .B(n394), .Y(n1717) );
  OAI21X1 U1331 ( .A(n1589), .B(n1656), .C(n1717), .Y(n2527) );
  NAND2X1 U1332 ( .A(\mem<29><5> ), .B(n394), .Y(n1718) );
  OAI21X1 U1333 ( .A(n1589), .B(n1658), .C(n1718), .Y(n2526) );
  NAND2X1 U1334 ( .A(\mem<29><6> ), .B(n394), .Y(n1719) );
  OAI21X1 U1335 ( .A(n1589), .B(n1660), .C(n1719), .Y(n2525) );
  NAND2X1 U1336 ( .A(\mem<29><7> ), .B(n394), .Y(n1720) );
  OAI21X1 U1337 ( .A(n1589), .B(n1662), .C(n1720), .Y(n2524) );
  NAND2X1 U1338 ( .A(\mem<29><8> ), .B(n394), .Y(n1721) );
  OAI21X1 U1339 ( .A(n1590), .B(n1665), .C(n1721), .Y(n2523) );
  NAND2X1 U1340 ( .A(\mem<29><9> ), .B(n394), .Y(n1722) );
  OAI21X1 U1341 ( .A(n1590), .B(n1667), .C(n1722), .Y(n2522) );
  NAND2X1 U1342 ( .A(\mem<29><10> ), .B(n394), .Y(n1723) );
  OAI21X1 U1343 ( .A(n1590), .B(n1669), .C(n1723), .Y(n2521) );
  NAND2X1 U1344 ( .A(\mem<29><11> ), .B(n394), .Y(n1724) );
  OAI21X1 U1345 ( .A(n1590), .B(n1671), .C(n1724), .Y(n2520) );
  NAND2X1 U1346 ( .A(\mem<29><12> ), .B(n394), .Y(n1725) );
  OAI21X1 U1347 ( .A(n1590), .B(n1673), .C(n1725), .Y(n2519) );
  NAND2X1 U1348 ( .A(\mem<29><13> ), .B(n394), .Y(n1726) );
  OAI21X1 U1349 ( .A(n1590), .B(n1675), .C(n1726), .Y(n2518) );
  NAND2X1 U1350 ( .A(\mem<29><14> ), .B(n394), .Y(n1727) );
  OAI21X1 U1351 ( .A(n1590), .B(n1677), .C(n1727), .Y(n2517) );
  NAND2X1 U1352 ( .A(\mem<29><15> ), .B(n394), .Y(n1728) );
  OAI21X1 U1353 ( .A(n1590), .B(n1679), .C(n1728), .Y(n2516) );
  NAND3X1 U1354 ( .A(\C2334/net89629 ), .B(net90019), .C(net90763), .Y(n1729)
         );
  NAND2X1 U1355 ( .A(\mem<28><0> ), .B(n396), .Y(n1730) );
  OAI21X1 U1356 ( .A(n1591), .B(n1648), .C(n1730), .Y(n2515) );
  NAND2X1 U1357 ( .A(\mem<28><1> ), .B(n396), .Y(n1731) );
  OAI21X1 U1358 ( .A(n1591), .B(n1651), .C(n1731), .Y(n2514) );
  NAND2X1 U1359 ( .A(\mem<28><2> ), .B(n396), .Y(n1732) );
  OAI21X1 U1360 ( .A(n1591), .B(n1653), .C(n1732), .Y(n2513) );
  NAND2X1 U1361 ( .A(\mem<28><3> ), .B(n396), .Y(n1733) );
  OAI21X1 U1362 ( .A(n1591), .B(n1655), .C(n1733), .Y(n2512) );
  NAND2X1 U1363 ( .A(\mem<28><4> ), .B(n396), .Y(n1734) );
  OAI21X1 U1364 ( .A(n1591), .B(n1657), .C(n1734), .Y(n2511) );
  NAND2X1 U1365 ( .A(\mem<28><5> ), .B(n396), .Y(n1735) );
  OAI21X1 U1366 ( .A(n1591), .B(n1659), .C(n1735), .Y(n2510) );
  NAND2X1 U1367 ( .A(\mem<28><6> ), .B(n396), .Y(n1736) );
  OAI21X1 U1368 ( .A(n1591), .B(n1661), .C(n1736), .Y(n2509) );
  NAND2X1 U1369 ( .A(\mem<28><7> ), .B(n396), .Y(n1737) );
  OAI21X1 U1370 ( .A(n1591), .B(n1663), .C(n1737), .Y(n2508) );
  NAND2X1 U1371 ( .A(\mem<28><8> ), .B(n396), .Y(n1738) );
  OAI21X1 U1372 ( .A(n1592), .B(n1664), .C(n1738), .Y(n2507) );
  NAND2X1 U1373 ( .A(\mem<28><9> ), .B(n396), .Y(n1739) );
  OAI21X1 U1374 ( .A(n1592), .B(n1666), .C(n1739), .Y(n2506) );
  NAND2X1 U1375 ( .A(\mem<28><10> ), .B(n396), .Y(n1740) );
  OAI21X1 U1376 ( .A(n1592), .B(n1668), .C(n1740), .Y(n2505) );
  NAND2X1 U1377 ( .A(\mem<28><11> ), .B(n396), .Y(n1741) );
  OAI21X1 U1378 ( .A(n1592), .B(n1671), .C(n1741), .Y(n2504) );
  NAND2X1 U1379 ( .A(\mem<28><12> ), .B(n396), .Y(n1742) );
  OAI21X1 U1380 ( .A(n1592), .B(n1673), .C(n1742), .Y(n2503) );
  NAND2X1 U1381 ( .A(\mem<28><13> ), .B(n396), .Y(n1743) );
  OAI21X1 U1382 ( .A(n1592), .B(n1675), .C(n1743), .Y(n2502) );
  NAND2X1 U1383 ( .A(\mem<28><14> ), .B(n396), .Y(n1744) );
  OAI21X1 U1384 ( .A(n1592), .B(n1677), .C(n1744), .Y(n2501) );
  NAND2X1 U1385 ( .A(\mem<28><15> ), .B(n396), .Y(n1745) );
  OAI21X1 U1386 ( .A(n1592), .B(n7), .C(n1745), .Y(n2500) );
  NAND3X1 U1387 ( .A(net90761), .B(\C2334/net89831 ), .C(net89545), .Y(n1746)
         );
  NAND2X1 U1388 ( .A(\mem<27><0> ), .B(n398), .Y(n1747) );
  OAI21X1 U1389 ( .A(n1593), .B(n1648), .C(n1747), .Y(n2499) );
  NAND2X1 U1390 ( .A(\mem<27><1> ), .B(n398), .Y(n1748) );
  OAI21X1 U1391 ( .A(n1593), .B(n1650), .C(n1748), .Y(n2498) );
  NAND2X1 U1392 ( .A(\mem<27><2> ), .B(n398), .Y(n1749) );
  OAI21X1 U1393 ( .A(n1593), .B(n1652), .C(n1749), .Y(n2497) );
  NAND2X1 U1394 ( .A(\mem<27><3> ), .B(n398), .Y(n1750) );
  OAI21X1 U1395 ( .A(n1593), .B(n1654), .C(n1750), .Y(n2496) );
  NAND2X1 U1396 ( .A(\mem<27><4> ), .B(n398), .Y(n1751) );
  OAI21X1 U1397 ( .A(n1593), .B(n1656), .C(n1751), .Y(n2495) );
  NAND2X1 U1398 ( .A(\mem<27><5> ), .B(n398), .Y(n1752) );
  OAI21X1 U1399 ( .A(n1593), .B(n1658), .C(n1752), .Y(n2494) );
  NAND2X1 U1400 ( .A(\mem<27><6> ), .B(n398), .Y(n1753) );
  OAI21X1 U1401 ( .A(n1593), .B(n1660), .C(n1753), .Y(n2493) );
  NAND2X1 U1402 ( .A(\mem<27><7> ), .B(n398), .Y(n1754) );
  OAI21X1 U1403 ( .A(n1593), .B(n1662), .C(n1754), .Y(n2492) );
  NAND2X1 U1404 ( .A(\mem<27><8> ), .B(n398), .Y(n1755) );
  OAI21X1 U1405 ( .A(n1594), .B(n1665), .C(n1755), .Y(n2491) );
  NAND2X1 U1406 ( .A(\mem<27><9> ), .B(n398), .Y(n1756) );
  OAI21X1 U1407 ( .A(n1594), .B(n1667), .C(n1756), .Y(n2490) );
  NAND2X1 U1408 ( .A(\mem<27><10> ), .B(n398), .Y(n1757) );
  OAI21X1 U1409 ( .A(n1594), .B(n1669), .C(n1757), .Y(n2489) );
  NAND2X1 U1410 ( .A(\mem<27><11> ), .B(n398), .Y(n1758) );
  OAI21X1 U1411 ( .A(n1594), .B(n1671), .C(n1758), .Y(n2488) );
  NAND2X1 U1412 ( .A(\mem<27><12> ), .B(n398), .Y(n1759) );
  OAI21X1 U1413 ( .A(n1594), .B(n1673), .C(n1759), .Y(n2487) );
  NAND2X1 U1414 ( .A(\mem<27><13> ), .B(n398), .Y(n1760) );
  OAI21X1 U1415 ( .A(n1594), .B(n1675), .C(n1760), .Y(n2486) );
  NAND2X1 U1416 ( .A(\mem<27><14> ), .B(n398), .Y(n1761) );
  OAI21X1 U1417 ( .A(n1594), .B(n1677), .C(n1761), .Y(n2485) );
  NAND2X1 U1418 ( .A(\mem<27><15> ), .B(n398), .Y(n1762) );
  OAI21X1 U1419 ( .A(n1594), .B(n1679), .C(n1762), .Y(n2484) );
  NAND3X1 U1420 ( .A(net89545), .B(\C2334/net89831 ), .C(net90763), .Y(n1763)
         );
  NAND2X1 U1421 ( .A(\mem<26><0> ), .B(n400), .Y(n1764) );
  OAI21X1 U1422 ( .A(n1595), .B(n1648), .C(n1764), .Y(n2483) );
  NAND2X1 U1423 ( .A(\mem<26><1> ), .B(n400), .Y(n1765) );
  OAI21X1 U1424 ( .A(n1595), .B(n1651), .C(n1765), .Y(n2482) );
  NAND2X1 U1425 ( .A(\mem<26><2> ), .B(n400), .Y(n1766) );
  OAI21X1 U1426 ( .A(n1595), .B(n1653), .C(n1766), .Y(n2481) );
  NAND2X1 U1427 ( .A(\mem<26><3> ), .B(n400), .Y(n1767) );
  OAI21X1 U1428 ( .A(n1595), .B(n1655), .C(n1767), .Y(n2480) );
  NAND2X1 U1429 ( .A(\mem<26><4> ), .B(n400), .Y(n1768) );
  OAI21X1 U1430 ( .A(n1595), .B(n1657), .C(n1768), .Y(n2479) );
  NAND2X1 U1431 ( .A(\mem<26><5> ), .B(n400), .Y(n1769) );
  OAI21X1 U1432 ( .A(n1595), .B(n1659), .C(n1769), .Y(n2478) );
  NAND2X1 U1433 ( .A(\mem<26><6> ), .B(n400), .Y(n1770) );
  OAI21X1 U1434 ( .A(n1595), .B(n1661), .C(n1770), .Y(n2477) );
  NAND2X1 U1435 ( .A(\mem<26><7> ), .B(n400), .Y(n1771) );
  OAI21X1 U1436 ( .A(n1595), .B(n1663), .C(n1771), .Y(n2476) );
  NAND2X1 U1437 ( .A(\mem<26><8> ), .B(n400), .Y(n1772) );
  OAI21X1 U1438 ( .A(n1596), .B(n1664), .C(n1772), .Y(n2475) );
  NAND2X1 U1439 ( .A(\mem<26><9> ), .B(n400), .Y(n1773) );
  OAI21X1 U1440 ( .A(n1596), .B(n1666), .C(n1773), .Y(n2474) );
  NAND2X1 U1441 ( .A(\mem<26><10> ), .B(n400), .Y(n1774) );
  OAI21X1 U1442 ( .A(n1596), .B(n1668), .C(n1774), .Y(n2473) );
  NAND2X1 U1443 ( .A(\mem<26><11> ), .B(n400), .Y(n1775) );
  OAI21X1 U1444 ( .A(n1596), .B(n1671), .C(n1775), .Y(n2472) );
  NAND2X1 U1445 ( .A(\mem<26><12> ), .B(n400), .Y(n1776) );
  OAI21X1 U1446 ( .A(n1596), .B(n1673), .C(n1776), .Y(n2471) );
  NAND2X1 U1447 ( .A(\mem<26><13> ), .B(n400), .Y(n1777) );
  OAI21X1 U1448 ( .A(n1596), .B(n1675), .C(n1777), .Y(n2470) );
  NAND2X1 U1449 ( .A(\mem<26><14> ), .B(n400), .Y(n1778) );
  OAI21X1 U1450 ( .A(n1596), .B(n1677), .C(n1778), .Y(n2469) );
  NAND2X1 U1451 ( .A(\mem<26><15> ), .B(n400), .Y(n1779) );
  OAI21X1 U1452 ( .A(n1596), .B(n1678), .C(n1779), .Y(n2468) );
  NAND3X1 U1453 ( .A(net90761), .B(net89545), .C(net90019), .Y(n1780) );
  NAND2X1 U1454 ( .A(\mem<25><0> ), .B(n402), .Y(n1781) );
  OAI21X1 U1455 ( .A(n1597), .B(n1648), .C(n1781), .Y(n2467) );
  NAND2X1 U1456 ( .A(\mem<25><1> ), .B(n402), .Y(n1782) );
  OAI21X1 U1457 ( .A(n1597), .B(n1650), .C(n1782), .Y(n2466) );
  NAND2X1 U1458 ( .A(\mem<25><2> ), .B(n402), .Y(n1783) );
  OAI21X1 U1459 ( .A(n1597), .B(n1652), .C(n1783), .Y(n2465) );
  NAND2X1 U1460 ( .A(\mem<25><3> ), .B(n402), .Y(n1784) );
  OAI21X1 U1461 ( .A(n1597), .B(n1654), .C(n1784), .Y(n2464) );
  NAND2X1 U1462 ( .A(\mem<25><4> ), .B(n402), .Y(n1785) );
  OAI21X1 U1463 ( .A(n1597), .B(n1656), .C(n1785), .Y(n2463) );
  NAND2X1 U1464 ( .A(\mem<25><5> ), .B(n402), .Y(n1786) );
  OAI21X1 U1465 ( .A(n1597), .B(n1658), .C(n1786), .Y(n2462) );
  NAND2X1 U1466 ( .A(\mem<25><6> ), .B(n402), .Y(n1787) );
  OAI21X1 U1467 ( .A(n1597), .B(n1660), .C(n1787), .Y(n2461) );
  NAND2X1 U1468 ( .A(\mem<25><7> ), .B(n402), .Y(n1788) );
  OAI21X1 U1469 ( .A(n1597), .B(n1662), .C(n1788), .Y(n2460) );
  NAND2X1 U1470 ( .A(\mem<25><8> ), .B(n402), .Y(n1789) );
  OAI21X1 U1471 ( .A(n1598), .B(n1665), .C(n1789), .Y(n2459) );
  NAND2X1 U1472 ( .A(\mem<25><9> ), .B(n402), .Y(n1790) );
  OAI21X1 U1473 ( .A(n1598), .B(n1667), .C(n1790), .Y(n2458) );
  NAND2X1 U1474 ( .A(\mem<25><10> ), .B(n402), .Y(n1791) );
  OAI21X1 U1475 ( .A(n1598), .B(n1669), .C(n1791), .Y(n2457) );
  NAND2X1 U1476 ( .A(\mem<25><11> ), .B(n402), .Y(n1792) );
  OAI21X1 U1477 ( .A(n1598), .B(n1671), .C(n1792), .Y(n2456) );
  NAND2X1 U1478 ( .A(\mem<25><12> ), .B(n402), .Y(n1793) );
  OAI21X1 U1479 ( .A(n1598), .B(n1673), .C(n1793), .Y(n2455) );
  NAND2X1 U1480 ( .A(\mem<25><13> ), .B(n402), .Y(n1794) );
  OAI21X1 U1481 ( .A(n1598), .B(n1675), .C(n1794), .Y(n2454) );
  NAND2X1 U1482 ( .A(\mem<25><14> ), .B(n402), .Y(n1795) );
  OAI21X1 U1483 ( .A(n1598), .B(n1677), .C(n1795), .Y(n2453) );
  NAND2X1 U1484 ( .A(\mem<25><15> ), .B(n402), .Y(n1796) );
  OAI21X1 U1485 ( .A(n1598), .B(n1679), .C(n1796), .Y(n2452) );
  NOR3X1 U1486 ( .A(net90761), .B(\C2334/net89831 ), .C(\C2334/net89629 ), .Y(
        n2042) );
  NAND2X1 U1487 ( .A(\mem<24><0> ), .B(n404), .Y(n1797) );
  OAI21X1 U1488 ( .A(n1599), .B(n1648), .C(n1797), .Y(n2451) );
  NAND2X1 U1489 ( .A(\mem<24><1> ), .B(n404), .Y(n1798) );
  OAI21X1 U1490 ( .A(n1599), .B(n1650), .C(n1798), .Y(n2450) );
  NAND2X1 U1491 ( .A(\mem<24><2> ), .B(n404), .Y(n1799) );
  OAI21X1 U1492 ( .A(n1599), .B(n1652), .C(n1799), .Y(n2449) );
  NAND2X1 U1493 ( .A(\mem<24><3> ), .B(n404), .Y(n1800) );
  OAI21X1 U1494 ( .A(n1599), .B(n1654), .C(n1800), .Y(n2448) );
  NAND2X1 U1495 ( .A(\mem<24><4> ), .B(n404), .Y(n1801) );
  OAI21X1 U1496 ( .A(n1599), .B(n1656), .C(n1801), .Y(n2447) );
  NAND2X1 U1497 ( .A(\mem<24><5> ), .B(n404), .Y(n1802) );
  OAI21X1 U1498 ( .A(n1599), .B(n1658), .C(n1802), .Y(n2446) );
  NAND2X1 U1499 ( .A(\mem<24><6> ), .B(n404), .Y(n1803) );
  OAI21X1 U1500 ( .A(n1599), .B(n1660), .C(n1803), .Y(n2445) );
  NAND2X1 U1501 ( .A(\mem<24><7> ), .B(n404), .Y(n1804) );
  OAI21X1 U1502 ( .A(n1599), .B(n1662), .C(n1804), .Y(n2444) );
  NAND2X1 U1503 ( .A(\mem<24><8> ), .B(n404), .Y(n1805) );
  OAI21X1 U1504 ( .A(n1599), .B(n1664), .C(n1805), .Y(n2443) );
  NAND2X1 U1505 ( .A(\mem<24><9> ), .B(n404), .Y(n1806) );
  OAI21X1 U1506 ( .A(n1599), .B(n1666), .C(n1806), .Y(n2442) );
  NAND2X1 U1507 ( .A(\mem<24><10> ), .B(n404), .Y(n1807) );
  OAI21X1 U1508 ( .A(n1599), .B(n1668), .C(n1807), .Y(n2441) );
  NAND2X1 U1509 ( .A(\mem<24><11> ), .B(n404), .Y(n1808) );
  OAI21X1 U1510 ( .A(n1599), .B(n1670), .C(n1808), .Y(n2440) );
  NAND2X1 U1511 ( .A(\mem<24><12> ), .B(n404), .Y(n1809) );
  OAI21X1 U1512 ( .A(n1599), .B(n1672), .C(n1809), .Y(n2439) );
  NAND2X1 U1513 ( .A(\mem<24><13> ), .B(n404), .Y(n1810) );
  OAI21X1 U1514 ( .A(n1599), .B(n1674), .C(n1810), .Y(n2438) );
  NAND2X1 U1515 ( .A(\mem<24><14> ), .B(n404), .Y(n1811) );
  OAI21X1 U1516 ( .A(n1599), .B(n1676), .C(n1811), .Y(n2437) );
  NAND2X1 U1517 ( .A(\mem<24><15> ), .B(n404), .Y(n1812) );
  OAI21X1 U1518 ( .A(n1599), .B(n1678), .C(n1812), .Y(n2436) );
  NAND2X1 U1519 ( .A(\mem<23><0> ), .B(n406), .Y(n1813) );
  OAI21X1 U1520 ( .A(n1600), .B(n1648), .C(n1813), .Y(n2435) );
  NAND2X1 U1521 ( .A(\mem<23><1> ), .B(n406), .Y(n1814) );
  OAI21X1 U1522 ( .A(n1600), .B(n1651), .C(n1814), .Y(n2434) );
  NAND2X1 U1523 ( .A(\mem<23><2> ), .B(n406), .Y(n1815) );
  OAI21X1 U1524 ( .A(n1600), .B(n1653), .C(n1815), .Y(n2433) );
  NAND2X1 U1525 ( .A(\mem<23><3> ), .B(n406), .Y(n1816) );
  OAI21X1 U1526 ( .A(n1600), .B(n1655), .C(n1816), .Y(n2432) );
  NAND2X1 U1527 ( .A(\mem<23><4> ), .B(n406), .Y(n1817) );
  OAI21X1 U1528 ( .A(n1600), .B(n1657), .C(n1817), .Y(n2431) );
  NAND2X1 U1529 ( .A(\mem<23><5> ), .B(n406), .Y(n1818) );
  OAI21X1 U1530 ( .A(n1600), .B(n1659), .C(n1818), .Y(n2430) );
  NAND2X1 U1531 ( .A(\mem<23><6> ), .B(n406), .Y(n1819) );
  OAI21X1 U1532 ( .A(n1600), .B(n1661), .C(n1819), .Y(n2429) );
  NAND2X1 U1533 ( .A(\mem<23><7> ), .B(n406), .Y(n1820) );
  OAI21X1 U1534 ( .A(n1600), .B(n1663), .C(n1820), .Y(n2428) );
  NAND2X1 U1535 ( .A(\mem<23><8> ), .B(n406), .Y(n1821) );
  OAI21X1 U1536 ( .A(n1601), .B(n1665), .C(n1821), .Y(n2427) );
  NAND2X1 U1537 ( .A(\mem<23><9> ), .B(n406), .Y(n1822) );
  OAI21X1 U1538 ( .A(n1601), .B(n1667), .C(n1822), .Y(n2426) );
  NAND2X1 U1539 ( .A(\mem<23><10> ), .B(n406), .Y(n1823) );
  OAI21X1 U1540 ( .A(n1601), .B(n1669), .C(n1823), .Y(n2425) );
  NAND2X1 U1541 ( .A(\mem<23><11> ), .B(n406), .Y(n1824) );
  OAI21X1 U1542 ( .A(n1601), .B(n1671), .C(n1824), .Y(n2424) );
  NAND2X1 U1543 ( .A(\mem<23><12> ), .B(n406), .Y(n1825) );
  OAI21X1 U1544 ( .A(n1601), .B(n1673), .C(n1825), .Y(n2423) );
  NAND2X1 U1545 ( .A(\mem<23><13> ), .B(n406), .Y(n1826) );
  OAI21X1 U1546 ( .A(n1601), .B(n1675), .C(n1826), .Y(n2422) );
  NAND2X1 U1547 ( .A(\mem<23><14> ), .B(n406), .Y(n1827) );
  OAI21X1 U1548 ( .A(n1601), .B(n1677), .C(n1827), .Y(n2421) );
  NAND2X1 U1549 ( .A(\mem<23><15> ), .B(n406), .Y(n1828) );
  OAI21X1 U1550 ( .A(n1601), .B(n1679), .C(n1828), .Y(n2420) );
  NAND2X1 U1551 ( .A(\mem<22><0> ), .B(n408), .Y(n1829) );
  OAI21X1 U1552 ( .A(n1602), .B(n1648), .C(n1829), .Y(n2419) );
  NAND2X1 U1553 ( .A(\mem<22><1> ), .B(n408), .Y(n1830) );
  OAI21X1 U1554 ( .A(n1602), .B(n1651), .C(n1830), .Y(n2418) );
  NAND2X1 U1555 ( .A(\mem<22><2> ), .B(n408), .Y(n1831) );
  OAI21X1 U1556 ( .A(n1602), .B(n1653), .C(n1831), .Y(n2417) );
  NAND2X1 U1557 ( .A(\mem<22><3> ), .B(n408), .Y(n1832) );
  OAI21X1 U1558 ( .A(n1602), .B(n1655), .C(n1832), .Y(n2416) );
  NAND2X1 U1559 ( .A(\mem<22><4> ), .B(n408), .Y(n1833) );
  OAI21X1 U1560 ( .A(n1602), .B(n1657), .C(n1833), .Y(n2415) );
  NAND2X1 U1561 ( .A(\mem<22><5> ), .B(n408), .Y(n1834) );
  OAI21X1 U1562 ( .A(n1602), .B(n1659), .C(n1834), .Y(n2414) );
  NAND2X1 U1563 ( .A(\mem<22><6> ), .B(n408), .Y(n1835) );
  OAI21X1 U1564 ( .A(n1602), .B(n1661), .C(n1835), .Y(n2413) );
  NAND2X1 U1565 ( .A(\mem<22><7> ), .B(n408), .Y(n1836) );
  OAI21X1 U1566 ( .A(n1602), .B(n1663), .C(n1836), .Y(n2412) );
  NAND2X1 U1567 ( .A(\mem<22><8> ), .B(n408), .Y(n1837) );
  OAI21X1 U1568 ( .A(n1603), .B(n1665), .C(n1837), .Y(n2411) );
  NAND2X1 U1569 ( .A(\mem<22><9> ), .B(n408), .Y(n1838) );
  OAI21X1 U1570 ( .A(n1603), .B(n1667), .C(n1838), .Y(n2410) );
  NAND2X1 U1571 ( .A(\mem<22><10> ), .B(n408), .Y(n1839) );
  OAI21X1 U1572 ( .A(n1603), .B(n1669), .C(n1839), .Y(n2409) );
  NAND2X1 U1573 ( .A(\mem<22><11> ), .B(n408), .Y(n1840) );
  OAI21X1 U1574 ( .A(n1603), .B(n1671), .C(n1840), .Y(n2408) );
  NAND2X1 U1575 ( .A(\mem<22><12> ), .B(n408), .Y(n1841) );
  OAI21X1 U1576 ( .A(n1603), .B(n1673), .C(n1841), .Y(n2407) );
  NAND2X1 U1577 ( .A(\mem<22><13> ), .B(n408), .Y(n1842) );
  OAI21X1 U1578 ( .A(n1603), .B(n1675), .C(n1842), .Y(n2406) );
  NAND2X1 U1579 ( .A(\mem<22><14> ), .B(n408), .Y(n1843) );
  OAI21X1 U1580 ( .A(n1603), .B(n1677), .C(n1843), .Y(n2405) );
  NAND2X1 U1581 ( .A(\mem<22><15> ), .B(n408), .Y(n1844) );
  OAI21X1 U1582 ( .A(n1603), .B(n1679), .C(n1844), .Y(n2404) );
  NAND2X1 U1583 ( .A(\mem<21><0> ), .B(n302), .Y(n1845) );
  OAI21X1 U1584 ( .A(n1604), .B(n1648), .C(n1845), .Y(n2403) );
  NAND2X1 U1585 ( .A(\mem<21><1> ), .B(n302), .Y(n1846) );
  OAI21X1 U1586 ( .A(n1604), .B(n1651), .C(n1846), .Y(n2402) );
  NAND2X1 U1587 ( .A(\mem<21><2> ), .B(n302), .Y(n1847) );
  OAI21X1 U1588 ( .A(n1604), .B(n1653), .C(n1847), .Y(n2401) );
  NAND2X1 U1589 ( .A(\mem<21><3> ), .B(n302), .Y(n1848) );
  OAI21X1 U1590 ( .A(n1604), .B(n1655), .C(n1848), .Y(n2400) );
  NAND2X1 U1591 ( .A(\mem<21><4> ), .B(n302), .Y(n1849) );
  OAI21X1 U1592 ( .A(n1604), .B(n1657), .C(n1849), .Y(n2399) );
  NAND2X1 U1593 ( .A(\mem<21><5> ), .B(n302), .Y(n1850) );
  OAI21X1 U1594 ( .A(n1604), .B(n1659), .C(n1850), .Y(n2398) );
  NAND2X1 U1595 ( .A(\mem<21><6> ), .B(n302), .Y(n1851) );
  OAI21X1 U1596 ( .A(n1604), .B(n1661), .C(n1851), .Y(n2397) );
  NAND2X1 U1597 ( .A(\mem<21><7> ), .B(n302), .Y(n1852) );
  OAI21X1 U1598 ( .A(n1604), .B(n1663), .C(n1852), .Y(n2396) );
  NAND2X1 U1599 ( .A(\mem<21><8> ), .B(n302), .Y(n1853) );
  OAI21X1 U1600 ( .A(n1605), .B(n1665), .C(n1853), .Y(n2395) );
  NAND2X1 U1601 ( .A(\mem<21><9> ), .B(n302), .Y(n1854) );
  OAI21X1 U1602 ( .A(n1605), .B(n1667), .C(n1854), .Y(n2394) );
  NAND2X1 U1603 ( .A(\mem<21><10> ), .B(n302), .Y(n1855) );
  OAI21X1 U1604 ( .A(n1605), .B(n1669), .C(n1855), .Y(n2393) );
  NAND2X1 U1605 ( .A(\mem<21><11> ), .B(n302), .Y(n1856) );
  OAI21X1 U1606 ( .A(n1605), .B(n1671), .C(n1856), .Y(n2392) );
  NAND2X1 U1607 ( .A(\mem<21><12> ), .B(n302), .Y(n1857) );
  OAI21X1 U1608 ( .A(n1605), .B(n1673), .C(n1857), .Y(n2391) );
  NAND2X1 U1609 ( .A(\mem<21><13> ), .B(n302), .Y(n1858) );
  OAI21X1 U1610 ( .A(n1605), .B(n1675), .C(n1858), .Y(n2390) );
  NAND2X1 U1611 ( .A(\mem<21><14> ), .B(n302), .Y(n1859) );
  OAI21X1 U1612 ( .A(n1605), .B(n1677), .C(n1859), .Y(n2389) );
  NAND2X1 U1613 ( .A(\mem<21><15> ), .B(n302), .Y(n1860) );
  OAI21X1 U1614 ( .A(n1605), .B(n1679), .C(n1860), .Y(n2388) );
  NAND2X1 U1615 ( .A(\mem<20><0> ), .B(n332), .Y(n1861) );
  OAI21X1 U1616 ( .A(n1606), .B(n1648), .C(n1861), .Y(n2387) );
  NAND2X1 U1617 ( .A(\mem<20><1> ), .B(n332), .Y(n1862) );
  OAI21X1 U1618 ( .A(n1606), .B(n1651), .C(n1862), .Y(n2386) );
  NAND2X1 U1619 ( .A(\mem<20><2> ), .B(n332), .Y(n1863) );
  OAI21X1 U1620 ( .A(n1606), .B(n1653), .C(n1863), .Y(n2385) );
  NAND2X1 U1621 ( .A(\mem<20><3> ), .B(n332), .Y(n1864) );
  OAI21X1 U1622 ( .A(n1606), .B(n1655), .C(n1864), .Y(n2384) );
  NAND2X1 U1623 ( .A(\mem<20><4> ), .B(n332), .Y(n1865) );
  OAI21X1 U1624 ( .A(n1606), .B(n1657), .C(n1865), .Y(n2383) );
  NAND2X1 U1625 ( .A(\mem<20><5> ), .B(n332), .Y(n1866) );
  OAI21X1 U1626 ( .A(n1606), .B(n1659), .C(n1866), .Y(n2382) );
  NAND2X1 U1627 ( .A(\mem<20><6> ), .B(n332), .Y(n1867) );
  OAI21X1 U1628 ( .A(n1606), .B(n1661), .C(n1867), .Y(n2381) );
  NAND2X1 U1629 ( .A(\mem<20><7> ), .B(n332), .Y(n1868) );
  OAI21X1 U1630 ( .A(n1606), .B(n1663), .C(n1868), .Y(n2380) );
  OAI21X1 U1631 ( .A(n1607), .B(n1665), .C(n87), .Y(n2379) );
  OAI21X1 U1632 ( .A(n1607), .B(n1667), .C(n89), .Y(n2378) );
  OAI21X1 U1633 ( .A(n1607), .B(n1669), .C(n91), .Y(n2377) );
  OAI21X1 U1634 ( .A(n1607), .B(n1671), .C(n93), .Y(n2376) );
  OAI21X1 U1635 ( .A(n1607), .B(n1673), .C(n95), .Y(n2375) );
  OAI21X1 U1636 ( .A(n1607), .B(n1675), .C(n97), .Y(n2374) );
  OAI21X1 U1637 ( .A(n1607), .B(n1677), .C(n99), .Y(n2373) );
  NAND2X1 U1638 ( .A(\mem<20><15> ), .B(n332), .Y(n1869) );
  OAI21X1 U1639 ( .A(n1607), .B(n1679), .C(n1869), .Y(n2372) );
  NAND2X1 U1640 ( .A(\mem<19><0> ), .B(n41), .Y(n1870) );
  OAI21X1 U1641 ( .A(n1608), .B(n1648), .C(n1870), .Y(n2371) );
  NAND2X1 U1642 ( .A(\mem<19><1> ), .B(n40), .Y(n1871) );
  OAI21X1 U1643 ( .A(n1608), .B(n1651), .C(n1871), .Y(n2370) );
  NAND2X1 U1644 ( .A(\mem<19><2> ), .B(n41), .Y(n1872) );
  OAI21X1 U1645 ( .A(n1608), .B(n1653), .C(n1872), .Y(n2369) );
  NAND2X1 U1646 ( .A(\mem<19><3> ), .B(n41), .Y(n1873) );
  OAI21X1 U1647 ( .A(n1608), .B(n1655), .C(n1873), .Y(n2368) );
  NAND2X1 U1648 ( .A(\mem<19><4> ), .B(n40), .Y(n1874) );
  OAI21X1 U1649 ( .A(n1608), .B(n1657), .C(n1874), .Y(n2367) );
  NAND2X1 U1650 ( .A(\mem<19><5> ), .B(n41), .Y(n1875) );
  OAI21X1 U1651 ( .A(n1608), .B(n1659), .C(n1875), .Y(n2366) );
  NAND2X1 U1652 ( .A(\mem<19><6> ), .B(n40), .Y(n1876) );
  OAI21X1 U1653 ( .A(n1608), .B(n1661), .C(n1876), .Y(n2365) );
  NAND2X1 U1654 ( .A(\mem<19><7> ), .B(n41), .Y(n1877) );
  OAI21X1 U1655 ( .A(n1608), .B(n1663), .C(n1877), .Y(n2364) );
  OAI21X1 U1656 ( .A(n1609), .B(n1665), .C(n101), .Y(n2363) );
  OAI21X1 U1657 ( .A(n1609), .B(n1667), .C(n103), .Y(n2362) );
  OAI21X1 U1658 ( .A(n1609), .B(n1669), .C(n105), .Y(n2361) );
  OAI21X1 U1659 ( .A(n1609), .B(n1671), .C(n107), .Y(n2360) );
  OAI21X1 U1660 ( .A(n1609), .B(n1673), .C(n109), .Y(n2359) );
  OAI21X1 U1661 ( .A(n1609), .B(n1675), .C(n111), .Y(n2358) );
  OAI21X1 U1662 ( .A(n1609), .B(n1677), .C(n113), .Y(n2357) );
  NAND2X1 U1663 ( .A(\mem<19><15> ), .B(n40), .Y(n1878) );
  OAI21X1 U1664 ( .A(n1609), .B(n1679), .C(n1878), .Y(n2356) );
  NAND2X1 U1665 ( .A(\mem<18><0> ), .B(n39), .Y(n1879) );
  OAI21X1 U1666 ( .A(n1610), .B(n1649), .C(n1879), .Y(n2355) );
  NAND2X1 U1667 ( .A(\mem<18><1> ), .B(n38), .Y(n1880) );
  OAI21X1 U1668 ( .A(n1610), .B(n1651), .C(n1880), .Y(n2354) );
  NAND2X1 U1669 ( .A(\mem<18><2> ), .B(n39), .Y(n1881) );
  OAI21X1 U1670 ( .A(n1610), .B(n1653), .C(n1881), .Y(n2353) );
  NAND2X1 U1671 ( .A(\mem<18><3> ), .B(n39), .Y(n1882) );
  OAI21X1 U1672 ( .A(n1610), .B(n1655), .C(n1882), .Y(n2352) );
  NAND2X1 U1673 ( .A(\mem<18><4> ), .B(n38), .Y(n1883) );
  OAI21X1 U1674 ( .A(n1610), .B(n1657), .C(n1883), .Y(n2351) );
  NAND2X1 U1675 ( .A(\mem<18><5> ), .B(n39), .Y(n1884) );
  OAI21X1 U1676 ( .A(n1610), .B(n1659), .C(n1884), .Y(n2350) );
  NAND2X1 U1677 ( .A(\mem<18><6> ), .B(n38), .Y(n1885) );
  OAI21X1 U1678 ( .A(n1610), .B(n1661), .C(n1885), .Y(n2349) );
  NAND2X1 U1679 ( .A(\mem<18><7> ), .B(n39), .Y(n1886) );
  OAI21X1 U1680 ( .A(n1610), .B(n1663), .C(n1886), .Y(n2348) );
  OAI21X1 U1681 ( .A(n1611), .B(n1665), .C(n115), .Y(n2347) );
  OAI21X1 U1682 ( .A(n1611), .B(n1667), .C(n117), .Y(n2346) );
  OAI21X1 U1683 ( .A(n1611), .B(n1669), .C(n119), .Y(n2345) );
  OAI21X1 U1684 ( .A(n1611), .B(n5), .C(n121), .Y(n2344) );
  OAI21X1 U1685 ( .A(n1611), .B(n4), .C(n123), .Y(n2343) );
  OAI21X1 U1686 ( .A(n1611), .B(n3), .C(n125), .Y(n2342) );
  OAI21X1 U1687 ( .A(n1611), .B(n1677), .C(n127), .Y(n2341) );
  NAND2X1 U1688 ( .A(\mem<18><15> ), .B(n38), .Y(n1887) );
  OAI21X1 U1689 ( .A(n1611), .B(n1679), .C(n1887), .Y(n2340) );
  NAND2X1 U1690 ( .A(\mem<17><0> ), .B(n37), .Y(n1888) );
  OAI21X1 U1691 ( .A(n1612), .B(n1648), .C(n1888), .Y(n2339) );
  NAND2X1 U1692 ( .A(\mem<17><1> ), .B(n36), .Y(n1889) );
  OAI21X1 U1693 ( .A(n1612), .B(n1651), .C(n1889), .Y(n2338) );
  NAND2X1 U1694 ( .A(\mem<17><2> ), .B(n37), .Y(n1890) );
  OAI21X1 U1695 ( .A(n1612), .B(n1653), .C(n1890), .Y(n2337) );
  NAND2X1 U1696 ( .A(\mem<17><3> ), .B(n37), .Y(n1891) );
  OAI21X1 U1697 ( .A(n1612), .B(n1655), .C(n1891), .Y(n2336) );
  NAND2X1 U1698 ( .A(\mem<17><4> ), .B(n36), .Y(n1892) );
  OAI21X1 U1699 ( .A(n1612), .B(n1657), .C(n1892), .Y(n2335) );
  NAND2X1 U1700 ( .A(\mem<17><5> ), .B(n37), .Y(n1893) );
  OAI21X1 U1701 ( .A(n1612), .B(n1659), .C(n1893), .Y(n2334) );
  NAND2X1 U1702 ( .A(\mem<17><6> ), .B(n36), .Y(n1894) );
  OAI21X1 U1703 ( .A(n1612), .B(n1661), .C(n1894), .Y(n2333) );
  NAND2X1 U1704 ( .A(\mem<17><7> ), .B(n37), .Y(n1895) );
  OAI21X1 U1705 ( .A(n1612), .B(n1663), .C(n1895), .Y(n2332) );
  OAI21X1 U1706 ( .A(n1613), .B(n1665), .C(n129), .Y(n2331) );
  OAI21X1 U1707 ( .A(n1613), .B(n1667), .C(n131), .Y(n2330) );
  OAI21X1 U1708 ( .A(n1613), .B(n1669), .C(n133), .Y(n2329) );
  OAI21X1 U1709 ( .A(n1613), .B(n5), .C(n135), .Y(n2328) );
  OAI21X1 U1710 ( .A(n1613), .B(n4), .C(n137), .Y(n2327) );
  OAI21X1 U1711 ( .A(n1613), .B(n3), .C(n139), .Y(n2326) );
  OAI21X1 U1712 ( .A(n1613), .B(n1677), .C(n141), .Y(n2325) );
  NAND2X1 U1713 ( .A(\mem<17><15> ), .B(n36), .Y(n1896) );
  OAI21X1 U1714 ( .A(n1613), .B(n1679), .C(n1896), .Y(n2324) );
  NAND2X1 U1715 ( .A(\mem<16><0> ), .B(n340), .Y(n1897) );
  OAI21X1 U1716 ( .A(n1614), .B(n1649), .C(n1897), .Y(n2323) );
  NAND2X1 U1717 ( .A(\mem<16><1> ), .B(n340), .Y(n1898) );
  OAI21X1 U1718 ( .A(n1614), .B(n1651), .C(n1898), .Y(n2322) );
  NAND2X1 U1719 ( .A(\mem<16><2> ), .B(n340), .Y(n1899) );
  OAI21X1 U1720 ( .A(n1614), .B(n1653), .C(n1899), .Y(n2321) );
  NAND2X1 U1721 ( .A(\mem<16><3> ), .B(n340), .Y(n1900) );
  OAI21X1 U1722 ( .A(n1614), .B(n1655), .C(n1900), .Y(n2320) );
  NAND2X1 U1723 ( .A(\mem<16><4> ), .B(n340), .Y(n1901) );
  OAI21X1 U1724 ( .A(n1614), .B(n1657), .C(n1901), .Y(n2319) );
  NAND2X1 U1725 ( .A(\mem<16><5> ), .B(n340), .Y(n1902) );
  OAI21X1 U1726 ( .A(n1614), .B(n1659), .C(n1902), .Y(n2318) );
  NAND2X1 U1727 ( .A(\mem<16><6> ), .B(n340), .Y(n1903) );
  OAI21X1 U1728 ( .A(n1614), .B(n1661), .C(n1903), .Y(n2317) );
  NAND2X1 U1729 ( .A(\mem<16><7> ), .B(n340), .Y(n1904) );
  OAI21X1 U1730 ( .A(n1614), .B(n1663), .C(n1904), .Y(n2316) );
  OAI21X1 U1731 ( .A(n1614), .B(n1665), .C(n143), .Y(n2315) );
  OAI21X1 U1732 ( .A(n1614), .B(n1667), .C(n145), .Y(n2314) );
  OAI21X1 U1733 ( .A(n1614), .B(n1669), .C(n147), .Y(n2313) );
  OAI21X1 U1734 ( .A(n1614), .B(n1671), .C(n149), .Y(n2312) );
  OAI21X1 U1735 ( .A(n1614), .B(n1673), .C(n151), .Y(n2311) );
  OAI21X1 U1736 ( .A(n1614), .B(n1675), .C(n153), .Y(n2310) );
  NAND2X1 U1737 ( .A(\mem<16><14> ), .B(n340), .Y(n1905) );
  OAI21X1 U1738 ( .A(n1614), .B(n1677), .C(n1905), .Y(n2309) );
  OAI21X1 U1739 ( .A(n1614), .B(n1679), .C(n155), .Y(n2308) );
  NAND3X1 U1740 ( .A(net89383), .B(n2564), .C(net89253), .Y(n1906) );
  NAND2X1 U1741 ( .A(\mem<15><0> ), .B(n35), .Y(n1907) );
  OAI21X1 U1742 ( .A(n1615), .B(n1649), .C(n1907), .Y(n2307) );
  NAND2X1 U1743 ( .A(\mem<15><1> ), .B(n34), .Y(n1908) );
  OAI21X1 U1744 ( .A(n1615), .B(n1651), .C(n1908), .Y(n2306) );
  NAND2X1 U1745 ( .A(\mem<15><2> ), .B(n35), .Y(n1909) );
  OAI21X1 U1746 ( .A(n1615), .B(n1653), .C(n1909), .Y(n2305) );
  NAND2X1 U1747 ( .A(\mem<15><3> ), .B(n35), .Y(n1910) );
  OAI21X1 U1748 ( .A(n1615), .B(n1655), .C(n1910), .Y(n2304) );
  NAND2X1 U1749 ( .A(\mem<15><4> ), .B(n34), .Y(n1911) );
  OAI21X1 U1750 ( .A(n1615), .B(n1657), .C(n1911), .Y(n2303) );
  NAND2X1 U1751 ( .A(\mem<15><5> ), .B(n35), .Y(n1912) );
  OAI21X1 U1752 ( .A(n1615), .B(n1659), .C(n1912), .Y(n2302) );
  NAND2X1 U1753 ( .A(\mem<15><6> ), .B(n34), .Y(n1913) );
  OAI21X1 U1754 ( .A(n1615), .B(n1661), .C(n1913), .Y(n2301) );
  NAND2X1 U1755 ( .A(\mem<15><7> ), .B(n35), .Y(n1914) );
  OAI21X1 U1756 ( .A(n1615), .B(n1663), .C(n1914), .Y(n2300) );
  OAI21X1 U1757 ( .A(n1616), .B(n1665), .C(n157), .Y(n2299) );
  OAI21X1 U1758 ( .A(n1616), .B(n1667), .C(n159), .Y(n2298) );
  OAI21X1 U1759 ( .A(n1616), .B(n1669), .C(n161), .Y(n2297) );
  OAI21X1 U1760 ( .A(n1616), .B(n5), .C(n163), .Y(n2296) );
  OAI21X1 U1761 ( .A(n1616), .B(n4), .C(n165), .Y(n2295) );
  OAI21X1 U1762 ( .A(n1616), .B(n3), .C(n167), .Y(n2294) );
  OAI21X1 U1763 ( .A(n1616), .B(n1677), .C(n169), .Y(n2293) );
  NAND2X1 U1764 ( .A(\mem<15><15> ), .B(n34), .Y(n1915) );
  OAI21X1 U1765 ( .A(n1616), .B(n1679), .C(n1915), .Y(n2292) );
  NAND2X1 U1766 ( .A(\mem<14><0> ), .B(n33), .Y(n1916) );
  OAI21X1 U1767 ( .A(n1617), .B(n1648), .C(n1916), .Y(n2291) );
  NAND2X1 U1768 ( .A(\mem<14><1> ), .B(n32), .Y(n1917) );
  OAI21X1 U1769 ( .A(n1617), .B(n1651), .C(n1917), .Y(n2290) );
  NAND2X1 U1770 ( .A(\mem<14><2> ), .B(n33), .Y(n1918) );
  OAI21X1 U1771 ( .A(n1617), .B(n1653), .C(n1918), .Y(n2289) );
  NAND2X1 U1772 ( .A(\mem<14><3> ), .B(n33), .Y(n1919) );
  OAI21X1 U1773 ( .A(n1617), .B(n1655), .C(n1919), .Y(n2288) );
  NAND2X1 U1774 ( .A(\mem<14><4> ), .B(n32), .Y(n1920) );
  OAI21X1 U1775 ( .A(n1617), .B(n1657), .C(n1920), .Y(n2287) );
  NAND2X1 U1776 ( .A(\mem<14><5> ), .B(n33), .Y(n1921) );
  OAI21X1 U1777 ( .A(n1617), .B(n1659), .C(n1921), .Y(n2286) );
  NAND2X1 U1778 ( .A(\mem<14><6> ), .B(n32), .Y(n1922) );
  OAI21X1 U1779 ( .A(n1617), .B(n1661), .C(n1922), .Y(n2285) );
  NAND2X1 U1780 ( .A(\mem<14><7> ), .B(n33), .Y(n1923) );
  OAI21X1 U1781 ( .A(n1617), .B(n1663), .C(n1923), .Y(n2284) );
  OAI21X1 U1782 ( .A(n1618), .B(n1665), .C(n171), .Y(n2283) );
  OAI21X1 U1783 ( .A(n1618), .B(n1667), .C(n173), .Y(n2282) );
  OAI21X1 U1784 ( .A(n1618), .B(n1669), .C(n175), .Y(n2281) );
  OAI21X1 U1785 ( .A(n1618), .B(n47), .C(n177), .Y(n2280) );
  OAI21X1 U1786 ( .A(n1618), .B(n46), .C(n179), .Y(n2279) );
  OAI21X1 U1787 ( .A(n1618), .B(n45), .C(n181), .Y(n2278) );
  OAI21X1 U1788 ( .A(n1618), .B(n44), .C(n183), .Y(n2277) );
  NAND2X1 U1789 ( .A(\mem<14><15> ), .B(n32), .Y(n1924) );
  OAI21X1 U1790 ( .A(n1618), .B(n1679), .C(n1924), .Y(n2276) );
  NAND2X1 U1791 ( .A(\mem<13><0> ), .B(n31), .Y(n1925) );
  OAI21X1 U1792 ( .A(n1619), .B(n1649), .C(n1925), .Y(n2275) );
  NAND2X1 U1793 ( .A(\mem<13><1> ), .B(n30), .Y(n1926) );
  OAI21X1 U1794 ( .A(n1619), .B(n1651), .C(n1926), .Y(n2274) );
  NAND2X1 U1795 ( .A(\mem<13><2> ), .B(n31), .Y(n1927) );
  OAI21X1 U1796 ( .A(n1619), .B(n1653), .C(n1927), .Y(n2273) );
  NAND2X1 U1797 ( .A(\mem<13><3> ), .B(n31), .Y(n1928) );
  OAI21X1 U1798 ( .A(n1619), .B(n1655), .C(n1928), .Y(n2272) );
  NAND2X1 U1799 ( .A(\mem<13><4> ), .B(n30), .Y(n1929) );
  OAI21X1 U1800 ( .A(n1619), .B(n1657), .C(n1929), .Y(n2271) );
  NAND2X1 U1801 ( .A(\mem<13><5> ), .B(n31), .Y(n1930) );
  OAI21X1 U1802 ( .A(n1619), .B(n1659), .C(n1930), .Y(n2270) );
  NAND2X1 U1803 ( .A(\mem<13><6> ), .B(n30), .Y(n1931) );
  OAI21X1 U1804 ( .A(n1619), .B(n1661), .C(n1931), .Y(n2269) );
  NAND2X1 U1805 ( .A(\mem<13><7> ), .B(n31), .Y(n1932) );
  OAI21X1 U1806 ( .A(n1619), .B(n1663), .C(n1932), .Y(n2268) );
  OAI21X1 U1807 ( .A(n1620), .B(n1665), .C(n185), .Y(n2267) );
  OAI21X1 U1808 ( .A(n1620), .B(n1667), .C(n187), .Y(n2266) );
  OAI21X1 U1809 ( .A(n1620), .B(n1669), .C(n189), .Y(n2265) );
  OAI21X1 U1810 ( .A(n1620), .B(n47), .C(n191), .Y(n2264) );
  OAI21X1 U1811 ( .A(n1620), .B(n46), .C(n193), .Y(n2263) );
  OAI21X1 U1812 ( .A(n1620), .B(n45), .C(n195), .Y(n2262) );
  OAI21X1 U1813 ( .A(n1620), .B(n44), .C(n197), .Y(n2261) );
  NAND2X1 U1814 ( .A(\mem<13><15> ), .B(n30), .Y(n1933) );
  OAI21X1 U1815 ( .A(n1620), .B(n1679), .C(n1933), .Y(n2260) );
  NAND2X1 U1816 ( .A(\mem<12><0> ), .B(n29), .Y(n1934) );
  OAI21X1 U1817 ( .A(n1621), .B(n1648), .C(n1934), .Y(n2259) );
  NAND2X1 U1818 ( .A(\mem<12><1> ), .B(n28), .Y(n1935) );
  OAI21X1 U1819 ( .A(n1621), .B(n1651), .C(n1935), .Y(n2258) );
  NAND2X1 U1820 ( .A(\mem<12><2> ), .B(n29), .Y(n1936) );
  OAI21X1 U1821 ( .A(n1621), .B(n1653), .C(n1936), .Y(n2257) );
  NAND2X1 U1822 ( .A(\mem<12><3> ), .B(n29), .Y(n1937) );
  OAI21X1 U1823 ( .A(n1621), .B(n1655), .C(n1937), .Y(n2256) );
  NAND2X1 U1824 ( .A(\mem<12><4> ), .B(n28), .Y(n1938) );
  OAI21X1 U1825 ( .A(n1621), .B(n1657), .C(n1938), .Y(n2255) );
  NAND2X1 U1826 ( .A(\mem<12><5> ), .B(n29), .Y(n1939) );
  OAI21X1 U1827 ( .A(n1621), .B(n1659), .C(n1939), .Y(n2254) );
  NAND2X1 U1828 ( .A(\mem<12><6> ), .B(n28), .Y(n1940) );
  OAI21X1 U1829 ( .A(n1621), .B(n1661), .C(n1940), .Y(n2253) );
  NAND2X1 U1830 ( .A(\mem<12><7> ), .B(n29), .Y(n1941) );
  OAI21X1 U1831 ( .A(n1621), .B(n1663), .C(n1941), .Y(n2252) );
  OAI21X1 U1832 ( .A(n1622), .B(n1665), .C(n199), .Y(n2251) );
  OAI21X1 U1833 ( .A(n1622), .B(n1667), .C(n201), .Y(n2250) );
  OAI21X1 U1834 ( .A(n1622), .B(n1669), .C(n203), .Y(n2249) );
  OAI21X1 U1835 ( .A(n1622), .B(n47), .C(n205), .Y(n2248) );
  OAI21X1 U1836 ( .A(n1622), .B(n46), .C(n207), .Y(n2247) );
  OAI21X1 U1837 ( .A(n1622), .B(n45), .C(n209), .Y(n2246) );
  OAI21X1 U1838 ( .A(n1622), .B(n44), .C(n211), .Y(n2245) );
  NAND2X1 U1839 ( .A(\mem<12><15> ), .B(n28), .Y(n1942) );
  OAI21X1 U1840 ( .A(n1622), .B(n1679), .C(n1942), .Y(n2244) );
  NAND2X1 U1841 ( .A(\mem<11><0> ), .B(n27), .Y(n1943) );
  OAI21X1 U1842 ( .A(n1623), .B(n1649), .C(n1943), .Y(n2243) );
  NAND2X1 U1843 ( .A(\mem<11><1> ), .B(n26), .Y(n1944) );
  OAI21X1 U1844 ( .A(n1623), .B(n1650), .C(n1944), .Y(n2242) );
  NAND2X1 U1845 ( .A(\mem<11><2> ), .B(n27), .Y(n1945) );
  OAI21X1 U1846 ( .A(n1623), .B(n1652), .C(n1945), .Y(n2241) );
  NAND2X1 U1847 ( .A(\mem<11><3> ), .B(n27), .Y(n1946) );
  OAI21X1 U1848 ( .A(n1623), .B(n1654), .C(n1946), .Y(n2240) );
  NAND2X1 U1849 ( .A(\mem<11><4> ), .B(n26), .Y(n1947) );
  OAI21X1 U1850 ( .A(n1623), .B(n1656), .C(n1947), .Y(n2239) );
  NAND2X1 U1851 ( .A(\mem<11><5> ), .B(n27), .Y(n1948) );
  OAI21X1 U1852 ( .A(n1623), .B(n1658), .C(n1948), .Y(n2238) );
  NAND2X1 U1853 ( .A(\mem<11><6> ), .B(n26), .Y(n1949) );
  OAI21X1 U1854 ( .A(n1623), .B(n1660), .C(n1949), .Y(n2237) );
  NAND2X1 U1855 ( .A(\mem<11><7> ), .B(n27), .Y(n1950) );
  OAI21X1 U1856 ( .A(n1623), .B(n1662), .C(n1950), .Y(n2236) );
  OAI21X1 U1857 ( .A(n1624), .B(n1664), .C(n213), .Y(n2235) );
  OAI21X1 U1858 ( .A(n1624), .B(n1666), .C(n216), .Y(n2234) );
  OAI21X1 U1859 ( .A(n1624), .B(n1668), .C(n218), .Y(n2233) );
  OAI21X1 U1860 ( .A(n1624), .B(n1671), .C(n220), .Y(n2232) );
  OAI21X1 U1861 ( .A(n1624), .B(n1673), .C(n222), .Y(n2231) );
  OAI21X1 U1862 ( .A(n1624), .B(n1675), .C(n224), .Y(n2230) );
  OAI21X1 U1863 ( .A(n1624), .B(n1677), .C(n226), .Y(n2229) );
  NAND2X1 U1864 ( .A(\mem<11><15> ), .B(n26), .Y(n1951) );
  OAI21X1 U1865 ( .A(n1624), .B(n7), .C(n1951), .Y(n2228) );
  NAND2X1 U1866 ( .A(\mem<10><0> ), .B(n25), .Y(n1952) );
  OAI21X1 U1867 ( .A(n1625), .B(n1649), .C(n1952), .Y(n2227) );
  NAND2X1 U1868 ( .A(\mem<10><1> ), .B(n24), .Y(n1953) );
  OAI21X1 U1869 ( .A(n1625), .B(n1650), .C(n1953), .Y(n2226) );
  NAND2X1 U1870 ( .A(\mem<10><2> ), .B(n25), .Y(n1954) );
  OAI21X1 U1871 ( .A(n1625), .B(n1652), .C(n1954), .Y(n2225) );
  NAND2X1 U1872 ( .A(\mem<10><3> ), .B(n25), .Y(n1955) );
  OAI21X1 U1873 ( .A(n1625), .B(n1654), .C(n1955), .Y(n2224) );
  NAND2X1 U1874 ( .A(\mem<10><4> ), .B(n24), .Y(n1956) );
  OAI21X1 U1875 ( .A(n1625), .B(n1656), .C(n1956), .Y(n2223) );
  NAND2X1 U1876 ( .A(\mem<10><5> ), .B(n25), .Y(n1957) );
  OAI21X1 U1877 ( .A(n1625), .B(n1658), .C(n1957), .Y(n2222) );
  NAND2X1 U1878 ( .A(\mem<10><6> ), .B(n24), .Y(n1958) );
  OAI21X1 U1879 ( .A(n1625), .B(n1660), .C(n1958), .Y(n2221) );
  NAND2X1 U1880 ( .A(\mem<10><7> ), .B(n25), .Y(n1959) );
  OAI21X1 U1881 ( .A(n1625), .B(n1662), .C(n1959), .Y(n2220) );
  OAI21X1 U1882 ( .A(n1626), .B(n1664), .C(n228), .Y(n2219) );
  OAI21X1 U1883 ( .A(n1626), .B(n1666), .C(n230), .Y(n2218) );
  OAI21X1 U1884 ( .A(n1626), .B(n1668), .C(n232), .Y(n2217) );
  OAI21X1 U1885 ( .A(n1626), .B(n1671), .C(n234), .Y(n2216) );
  OAI21X1 U1886 ( .A(n1626), .B(n1673), .C(n236), .Y(n2215) );
  OAI21X1 U1887 ( .A(n1626), .B(n1675), .C(n238), .Y(n2214) );
  OAI21X1 U1888 ( .A(n1626), .B(n1677), .C(n240), .Y(n2213) );
  NAND2X1 U1889 ( .A(\mem<10><15> ), .B(n24), .Y(n1960) );
  OAI21X1 U1890 ( .A(n1626), .B(n1678), .C(n1960), .Y(n2212) );
  NAND2X1 U1891 ( .A(\mem<9><0> ), .B(n23), .Y(n1961) );
  OAI21X1 U1892 ( .A(n1627), .B(n1649), .C(n1961), .Y(n2211) );
  NAND2X1 U1893 ( .A(\mem<9><1> ), .B(n22), .Y(n1962) );
  OAI21X1 U1894 ( .A(n1627), .B(n1650), .C(n1962), .Y(n2210) );
  NAND2X1 U1895 ( .A(\mem<9><2> ), .B(n23), .Y(n1963) );
  OAI21X1 U1896 ( .A(n1627), .B(n1652), .C(n1963), .Y(n2209) );
  NAND2X1 U1897 ( .A(\mem<9><3> ), .B(n23), .Y(n1964) );
  OAI21X1 U1898 ( .A(n1627), .B(n1654), .C(n1964), .Y(n2208) );
  NAND2X1 U1899 ( .A(\mem<9><4> ), .B(n22), .Y(n1965) );
  OAI21X1 U1900 ( .A(n1627), .B(n1656), .C(n1965), .Y(n2207) );
  NAND2X1 U1901 ( .A(\mem<9><5> ), .B(n23), .Y(n1966) );
  OAI21X1 U1902 ( .A(n1627), .B(n1658), .C(n1966), .Y(n2206) );
  NAND2X1 U1903 ( .A(\mem<9><6> ), .B(n22), .Y(n1967) );
  OAI21X1 U1904 ( .A(n1627), .B(n1660), .C(n1967), .Y(n2205) );
  NAND2X1 U1905 ( .A(\mem<9><7> ), .B(n23), .Y(n1968) );
  OAI21X1 U1906 ( .A(n1627), .B(n1662), .C(n1968), .Y(n2204) );
  OAI21X1 U1907 ( .A(n1628), .B(n1664), .C(n242), .Y(n2203) );
  OAI21X1 U1908 ( .A(n1628), .B(n1666), .C(n244), .Y(n2202) );
  OAI21X1 U1909 ( .A(n1628), .B(n1668), .C(n246), .Y(n2201) );
  OAI21X1 U1910 ( .A(n1628), .B(n1671), .C(n248), .Y(n2200) );
  OAI21X1 U1911 ( .A(n1628), .B(n1673), .C(n250), .Y(n2199) );
  OAI21X1 U1912 ( .A(n1628), .B(n1675), .C(n252), .Y(n2198) );
  OAI21X1 U1913 ( .A(n1628), .B(n1677), .C(n254), .Y(n2197) );
  NAND2X1 U1914 ( .A(\mem<9><15> ), .B(n22), .Y(n1969) );
  OAI21X1 U1915 ( .A(n1628), .B(n7), .C(n1969), .Y(n2196) );
  NAND2X1 U1916 ( .A(\mem<8><0> ), .B(n43), .Y(n1971) );
  OAI21X1 U1917 ( .A(n1629), .B(n1649), .C(n1971), .Y(n2195) );
  NAND2X1 U1918 ( .A(\mem<8><1> ), .B(n356), .Y(n1972) );
  OAI21X1 U1919 ( .A(n1629), .B(n1650), .C(n1972), .Y(n2194) );
  NAND2X1 U1920 ( .A(\mem<8><2> ), .B(n42), .Y(n1973) );
  OAI21X1 U1921 ( .A(n1629), .B(n1652), .C(n1973), .Y(n2193) );
  NAND2X1 U1922 ( .A(\mem<8><3> ), .B(n356), .Y(n1974) );
  OAI21X1 U1923 ( .A(n1629), .B(n1654), .C(n1974), .Y(n2192) );
  NAND2X1 U1924 ( .A(\mem<8><4> ), .B(n42), .Y(n1975) );
  OAI21X1 U1925 ( .A(n1629), .B(n1656), .C(n1975), .Y(n2191) );
  NAND2X1 U1926 ( .A(\mem<8><5> ), .B(n43), .Y(n1976) );
  OAI21X1 U1927 ( .A(n1629), .B(n1658), .C(n1976), .Y(n2190) );
  NAND2X1 U1928 ( .A(\mem<8><6> ), .B(n42), .Y(n1977) );
  OAI21X1 U1929 ( .A(n1629), .B(n1660), .C(n1977), .Y(n2189) );
  NAND2X1 U1930 ( .A(\mem<8><7> ), .B(n356), .Y(n1978) );
  OAI21X1 U1931 ( .A(n1629), .B(n1662), .C(n1978), .Y(n2188) );
  OAI21X1 U1932 ( .A(n1629), .B(n1664), .C(n256), .Y(n2187) );
  OAI21X1 U1933 ( .A(n1629), .B(n1666), .C(n258), .Y(n2186) );
  OAI21X1 U1934 ( .A(n1629), .B(n1668), .C(n374), .Y(n2185) );
  OAI21X1 U1935 ( .A(n1629), .B(n1670), .C(n426), .Y(n2184) );
  OAI21X1 U1936 ( .A(n1629), .B(n1672), .C(n428), .Y(n2183) );
  OAI21X1 U1937 ( .A(n1629), .B(n1674), .C(n430), .Y(n2182) );
  OAI21X1 U1938 ( .A(n1629), .B(n1676), .C(n432), .Y(n2181) );
  OAI21X1 U1939 ( .A(n1629), .B(n1678), .C(n434), .Y(n2180) );
  NAND3X1 U1940 ( .A(net89385), .B(n2564), .C(net89253), .Y(n1979) );
  NAND2X1 U1941 ( .A(\mem<7><0> ), .B(n20), .Y(n1980) );
  OAI21X1 U1942 ( .A(n1630), .B(n1649), .C(n1980), .Y(n2179) );
  NAND2X1 U1943 ( .A(\mem<7><1> ), .B(n21), .Y(n1981) );
  OAI21X1 U1944 ( .A(n1630), .B(n1650), .C(n1981), .Y(n2178) );
  NAND2X1 U1945 ( .A(\mem<7><2> ), .B(n21), .Y(n1982) );
  OAI21X1 U1946 ( .A(n1630), .B(n1652), .C(n1982), .Y(n2177) );
  NAND2X1 U1947 ( .A(\mem<7><3> ), .B(n21), .Y(n1983) );
  OAI21X1 U1948 ( .A(n1630), .B(n1654), .C(n1983), .Y(n2176) );
  NAND2X1 U1949 ( .A(\mem<7><4> ), .B(n20), .Y(n1984) );
  OAI21X1 U1950 ( .A(n1630), .B(n1656), .C(n1984), .Y(n2175) );
  NAND2X1 U1951 ( .A(\mem<7><5> ), .B(n20), .Y(n1985) );
  OAI21X1 U1952 ( .A(n1630), .B(n1658), .C(n1985), .Y(n2174) );
  NAND2X1 U1953 ( .A(\mem<7><6> ), .B(n21), .Y(n1986) );
  OAI21X1 U1954 ( .A(n1630), .B(n1660), .C(n1986), .Y(n2173) );
  NAND2X1 U1955 ( .A(\mem<7><7> ), .B(n20), .Y(n1987) );
  OAI21X1 U1956 ( .A(n1630), .B(n1662), .C(n1987), .Y(n2172) );
  OAI21X1 U1957 ( .A(n1631), .B(n1664), .C(n260), .Y(n2171) );
  OAI21X1 U1958 ( .A(n1631), .B(n1666), .C(n262), .Y(n2170) );
  OAI21X1 U1959 ( .A(n1631), .B(n1668), .C(n376), .Y(n2169) );
  OAI21X1 U1960 ( .A(n1631), .B(n1671), .C(n436), .Y(n2168) );
  OAI21X1 U1961 ( .A(n1631), .B(n1673), .C(n438), .Y(n2167) );
  OAI21X1 U1962 ( .A(n1631), .B(n1675), .C(n440), .Y(n2166) );
  OAI21X1 U1963 ( .A(n1631), .B(n1677), .C(n442), .Y(n2165) );
  OAI21X1 U1964 ( .A(n1631), .B(n1678), .C(n444), .Y(n2164) );
  NAND2X1 U1965 ( .A(\mem<6><0> ), .B(n18), .Y(n1988) );
  OAI21X1 U1966 ( .A(n1632), .B(n1649), .C(n1988), .Y(n2163) );
  NAND2X1 U1967 ( .A(\mem<6><1> ), .B(n19), .Y(n1989) );
  OAI21X1 U1968 ( .A(n1632), .B(n1650), .C(n1989), .Y(n2162) );
  NAND2X1 U1969 ( .A(\mem<6><2> ), .B(n19), .Y(n1990) );
  OAI21X1 U1970 ( .A(n1632), .B(n1652), .C(n1990), .Y(n2161) );
  NAND2X1 U1971 ( .A(\mem<6><3> ), .B(n19), .Y(n1991) );
  OAI21X1 U1972 ( .A(n1632), .B(n1654), .C(n1991), .Y(n2160) );
  NAND2X1 U1973 ( .A(\mem<6><4> ), .B(n18), .Y(n1992) );
  OAI21X1 U1974 ( .A(n1632), .B(n1656), .C(n1992), .Y(n2159) );
  NAND2X1 U1975 ( .A(\mem<6><5> ), .B(n18), .Y(n1993) );
  OAI21X1 U1976 ( .A(n1632), .B(n1658), .C(n1993), .Y(n2158) );
  NAND2X1 U1977 ( .A(\mem<6><6> ), .B(n19), .Y(n1994) );
  OAI21X1 U1978 ( .A(n1632), .B(n1660), .C(n1994), .Y(n2157) );
  NAND2X1 U1979 ( .A(\mem<6><7> ), .B(n18), .Y(n1995) );
  OAI21X1 U1980 ( .A(n1632), .B(n1662), .C(n1995), .Y(n2156) );
  OAI21X1 U1981 ( .A(n1633), .B(n1664), .C(n264), .Y(n2155) );
  OAI21X1 U1982 ( .A(n1633), .B(n1666), .C(n266), .Y(n2154) );
  OAI21X1 U1983 ( .A(n1633), .B(n1668), .C(n378), .Y(n2153) );
  OAI21X1 U1984 ( .A(n1633), .B(n1671), .C(n446), .Y(n2152) );
  OAI21X1 U1985 ( .A(n1633), .B(n1673), .C(n448), .Y(n2151) );
  OAI21X1 U1986 ( .A(n1633), .B(n1675), .C(n450), .Y(n2150) );
  OAI21X1 U1987 ( .A(n1633), .B(n1677), .C(n452), .Y(n2149) );
  OAI21X1 U1988 ( .A(n1633), .B(n7), .C(n454), .Y(n2148) );
  NAND2X1 U1989 ( .A(\mem<5><0> ), .B(n16), .Y(n1997) );
  OAI21X1 U1990 ( .A(n1634), .B(n1649), .C(n1997), .Y(n2147) );
  NAND2X1 U1991 ( .A(\mem<5><1> ), .B(n17), .Y(n1998) );
  OAI21X1 U1992 ( .A(n1634), .B(n1650), .C(n1998), .Y(n2146) );
  NAND2X1 U1993 ( .A(\mem<5><2> ), .B(n17), .Y(n1999) );
  OAI21X1 U1994 ( .A(n1634), .B(n1652), .C(n1999), .Y(n2145) );
  NAND2X1 U1995 ( .A(\mem<5><3> ), .B(n17), .Y(n2000) );
  OAI21X1 U1996 ( .A(n1634), .B(n1654), .C(n2000), .Y(n2144) );
  NAND2X1 U1997 ( .A(\mem<5><4> ), .B(n16), .Y(n2001) );
  OAI21X1 U1998 ( .A(n1634), .B(n1656), .C(n2001), .Y(n2143) );
  NAND2X1 U1999 ( .A(\mem<5><5> ), .B(n16), .Y(n2002) );
  OAI21X1 U2000 ( .A(n1634), .B(n1658), .C(n2002), .Y(n2142) );
  NAND2X1 U2001 ( .A(\mem<5><6> ), .B(n17), .Y(n2003) );
  OAI21X1 U2002 ( .A(n1634), .B(n1660), .C(n2003), .Y(n2141) );
  NAND2X1 U2003 ( .A(\mem<5><7> ), .B(n16), .Y(n2004) );
  OAI21X1 U2004 ( .A(n1634), .B(n1662), .C(n2004), .Y(n2140) );
  OAI21X1 U2005 ( .A(n1635), .B(n1664), .C(n268), .Y(n2139) );
  OAI21X1 U2006 ( .A(n1635), .B(n1666), .C(n270), .Y(n2138) );
  OAI21X1 U2007 ( .A(n1635), .B(n1668), .C(n380), .Y(n2137) );
  OAI21X1 U2008 ( .A(n1635), .B(n1671), .C(n456), .Y(n2136) );
  OAI21X1 U2009 ( .A(n1635), .B(n1673), .C(n458), .Y(n2135) );
  OAI21X1 U2010 ( .A(n1635), .B(n1675), .C(n460), .Y(n2134) );
  OAI21X1 U2011 ( .A(n1635), .B(n1677), .C(n462), .Y(n2133) );
  OAI21X1 U2012 ( .A(n1635), .B(n7), .C(n464), .Y(n2132) );
  NAND2X1 U2013 ( .A(\mem<4><0> ), .B(n14), .Y(n2006) );
  OAI21X1 U2014 ( .A(n1636), .B(n1649), .C(n2006), .Y(n2131) );
  NAND2X1 U2015 ( .A(\mem<4><1> ), .B(n15), .Y(n2007) );
  OAI21X1 U2016 ( .A(n1636), .B(n1650), .C(n2007), .Y(n2130) );
  NAND2X1 U2017 ( .A(\mem<4><2> ), .B(n15), .Y(n2008) );
  OAI21X1 U2018 ( .A(n1636), .B(n1652), .C(n2008), .Y(n2129) );
  NAND2X1 U2019 ( .A(\mem<4><3> ), .B(n15), .Y(n2009) );
  OAI21X1 U2020 ( .A(n1636), .B(n1654), .C(n2009), .Y(n2128) );
  NAND2X1 U2021 ( .A(\mem<4><4> ), .B(n14), .Y(n2010) );
  OAI21X1 U2022 ( .A(n1636), .B(n1656), .C(n2010), .Y(n2127) );
  NAND2X1 U2023 ( .A(\mem<4><5> ), .B(n14), .Y(n2011) );
  OAI21X1 U2024 ( .A(n1636), .B(n1658), .C(n2011), .Y(n2126) );
  NAND2X1 U2025 ( .A(\mem<4><6> ), .B(n15), .Y(n2012) );
  OAI21X1 U2026 ( .A(n1636), .B(n1660), .C(n2012), .Y(n2125) );
  NAND2X1 U2027 ( .A(\mem<4><7> ), .B(n14), .Y(n2013) );
  OAI21X1 U2028 ( .A(n1636), .B(n1662), .C(n2013), .Y(n2124) );
  OAI21X1 U2029 ( .A(n1637), .B(n1664), .C(n272), .Y(n2123) );
  OAI21X1 U2030 ( .A(n1637), .B(n1666), .C(n274), .Y(n2122) );
  OAI21X1 U2031 ( .A(n1637), .B(n1668), .C(n382), .Y(n2121) );
  OAI21X1 U2032 ( .A(n1637), .B(n1671), .C(n466), .Y(n2120) );
  OAI21X1 U2033 ( .A(n1637), .B(n1673), .C(n468), .Y(n2119) );
  OAI21X1 U2034 ( .A(n1637), .B(n1675), .C(n470), .Y(n2118) );
  OAI21X1 U2035 ( .A(n1637), .B(n1677), .C(n472), .Y(n2117) );
  OAI21X1 U2036 ( .A(n1637), .B(n7), .C(n474), .Y(n2116) );
  NAND2X1 U2037 ( .A(\mem<3><0> ), .B(n12), .Y(n2015) );
  OAI21X1 U2038 ( .A(n1638), .B(n1649), .C(n2015), .Y(n2115) );
  NAND2X1 U2039 ( .A(\mem<3><1> ), .B(n13), .Y(n2016) );
  OAI21X1 U2040 ( .A(n1638), .B(n1650), .C(n2016), .Y(n2114) );
  NAND2X1 U2041 ( .A(\mem<3><2> ), .B(n13), .Y(n2017) );
  OAI21X1 U2042 ( .A(n1638), .B(n1652), .C(n2017), .Y(n2113) );
  NAND2X1 U2043 ( .A(\mem<3><3> ), .B(n13), .Y(n2018) );
  OAI21X1 U2044 ( .A(n1638), .B(n1654), .C(n2018), .Y(n2112) );
  NAND2X1 U2045 ( .A(\mem<3><4> ), .B(n12), .Y(n2019) );
  OAI21X1 U2046 ( .A(n1638), .B(n1656), .C(n2019), .Y(n2111) );
  NAND2X1 U2047 ( .A(\mem<3><5> ), .B(n12), .Y(n2020) );
  OAI21X1 U2048 ( .A(n1638), .B(n1658), .C(n2020), .Y(n2110) );
  NAND2X1 U2049 ( .A(\mem<3><6> ), .B(n13), .Y(n2021) );
  OAI21X1 U2050 ( .A(n1638), .B(n1660), .C(n2021), .Y(n2109) );
  NAND2X1 U2051 ( .A(\mem<3><7> ), .B(n12), .Y(n2022) );
  OAI21X1 U2052 ( .A(n1638), .B(n1662), .C(n2022), .Y(n2108) );
  OAI21X1 U2053 ( .A(n1639), .B(n1664), .C(n276), .Y(n2107) );
  OAI21X1 U2054 ( .A(n1639), .B(n1666), .C(n278), .Y(n2106) );
  OAI21X1 U2055 ( .A(n1639), .B(n1668), .C(n384), .Y(n2105) );
  OAI21X1 U2056 ( .A(n1639), .B(n1671), .C(n476), .Y(n2104) );
  OAI21X1 U2057 ( .A(n1639), .B(n1673), .C(n478), .Y(n2103) );
  OAI21X1 U2058 ( .A(n1639), .B(n1675), .C(n480), .Y(n2102) );
  OAI21X1 U2059 ( .A(n1639), .B(n1677), .C(n482), .Y(n2101) );
  OAI21X1 U2060 ( .A(n1639), .B(n7), .C(n484), .Y(n2100) );
  NAND2X1 U2061 ( .A(\mem<2><0> ), .B(n10), .Y(n2024) );
  OAI21X1 U2062 ( .A(n1640), .B(n1649), .C(n2024), .Y(n2099) );
  NAND2X1 U2063 ( .A(\mem<2><1> ), .B(n11), .Y(n2025) );
  OAI21X1 U2064 ( .A(n1640), .B(n1650), .C(n2025), .Y(n2098) );
  NAND2X1 U2065 ( .A(\mem<2><2> ), .B(n11), .Y(n2026) );
  OAI21X1 U2066 ( .A(n1640), .B(n1652), .C(n2026), .Y(n2097) );
  NAND2X1 U2067 ( .A(\mem<2><3> ), .B(n11), .Y(n2027) );
  OAI21X1 U2068 ( .A(n1640), .B(n1654), .C(n2027), .Y(n2096) );
  NAND2X1 U2069 ( .A(\mem<2><4> ), .B(n10), .Y(n2028) );
  OAI21X1 U2070 ( .A(n1640), .B(n1656), .C(n2028), .Y(n2095) );
  NAND2X1 U2071 ( .A(\mem<2><5> ), .B(n10), .Y(n2029) );
  OAI21X1 U2072 ( .A(n1640), .B(n1658), .C(n2029), .Y(n2094) );
  NAND2X1 U2073 ( .A(\mem<2><6> ), .B(n11), .Y(n2030) );
  OAI21X1 U2074 ( .A(n1640), .B(n1660), .C(n2030), .Y(n2093) );
  NAND2X1 U2075 ( .A(\mem<2><7> ), .B(n10), .Y(n2031) );
  OAI21X1 U2076 ( .A(n1640), .B(n1662), .C(n2031), .Y(n2092) );
  OAI21X1 U2077 ( .A(n1641), .B(n1664), .C(n280), .Y(n2091) );
  OAI21X1 U2078 ( .A(n1641), .B(n1666), .C(n282), .Y(n2090) );
  OAI21X1 U2079 ( .A(n1641), .B(n1668), .C(n386), .Y(n2089) );
  OAI21X1 U2080 ( .A(n1641), .B(n1671), .C(n486), .Y(n2088) );
  OAI21X1 U2081 ( .A(n1641), .B(n1673), .C(n488), .Y(n2087) );
  OAI21X1 U2082 ( .A(n1641), .B(n1675), .C(n490), .Y(n2086) );
  OAI21X1 U2083 ( .A(n1641), .B(n1677), .C(n492), .Y(n2085) );
  OAI21X1 U2084 ( .A(n1641), .B(n7), .C(n494), .Y(n2084) );
  NAND2X1 U2085 ( .A(\mem<1><0> ), .B(n8), .Y(n2033) );
  OAI21X1 U2086 ( .A(n1642), .B(n1649), .C(n2033), .Y(n2083) );
  NAND2X1 U2087 ( .A(\mem<1><1> ), .B(n9), .Y(n2034) );
  OAI21X1 U2088 ( .A(n1642), .B(n1650), .C(n2034), .Y(n2082) );
  NAND2X1 U2089 ( .A(\mem<1><2> ), .B(n9), .Y(n2035) );
  OAI21X1 U2090 ( .A(n1642), .B(n1652), .C(n2035), .Y(n2081) );
  NAND2X1 U2091 ( .A(\mem<1><3> ), .B(n9), .Y(n2036) );
  OAI21X1 U2092 ( .A(n1642), .B(n1654), .C(n2036), .Y(n2080) );
  NAND2X1 U2093 ( .A(\mem<1><4> ), .B(n8), .Y(n2037) );
  OAI21X1 U2094 ( .A(n1642), .B(n1656), .C(n2037), .Y(n2079) );
  NAND2X1 U2095 ( .A(\mem<1><5> ), .B(n8), .Y(n2038) );
  OAI21X1 U2096 ( .A(n1642), .B(n1658), .C(n2038), .Y(n2078) );
  NAND2X1 U2097 ( .A(\mem<1><6> ), .B(n9), .Y(n2039) );
  OAI21X1 U2098 ( .A(n1642), .B(n1660), .C(n2039), .Y(n2077) );
  NAND2X1 U2099 ( .A(\mem<1><7> ), .B(n8), .Y(n2040) );
  OAI21X1 U2100 ( .A(n1642), .B(n1662), .C(n2040), .Y(n2076) );
  OAI21X1 U2101 ( .A(n1643), .B(n1664), .C(n284), .Y(n2075) );
  OAI21X1 U2102 ( .A(n1643), .B(n1666), .C(n286), .Y(n2074) );
  OAI21X1 U2103 ( .A(n1643), .B(n1668), .C(n388), .Y(n2073) );
  OAI21X1 U2104 ( .A(n1643), .B(n1670), .C(n496), .Y(n2072) );
  OAI21X1 U2105 ( .A(n1643), .B(n1672), .C(n498), .Y(n2071) );
  OAI21X1 U2106 ( .A(n1643), .B(n1674), .C(n500), .Y(n2070) );
  OAI21X1 U2107 ( .A(n1643), .B(n1676), .C(n502), .Y(n2069) );
  OAI21X1 U2108 ( .A(n1643), .B(n7), .C(n504), .Y(n2068) );
  NAND2X1 U2109 ( .A(\mem<0><0> ), .B(n48), .Y(n2043) );
  OAI21X1 U2110 ( .A(n1644), .B(n1649), .C(n2043), .Y(n2067) );
  NAND2X1 U2111 ( .A(\mem<0><1> ), .B(n48), .Y(n2044) );
  OAI21X1 U2112 ( .A(n1644), .B(n1650), .C(n2044), .Y(n2066) );
  NAND2X1 U2113 ( .A(\mem<0><2> ), .B(n49), .Y(n2045) );
  OAI21X1 U2114 ( .A(n1644), .B(n1652), .C(n2045), .Y(n2065) );
  NAND2X1 U2115 ( .A(\mem<0><3> ), .B(n49), .Y(n2046) );
  OAI21X1 U2116 ( .A(n1644), .B(n1654), .C(n2046), .Y(n2064) );
  NAND2X1 U2117 ( .A(\mem<0><4> ), .B(n49), .Y(n2047) );
  OAI21X1 U2118 ( .A(n1644), .B(n1656), .C(n2047), .Y(n2063) );
  NAND2X1 U2119 ( .A(\mem<0><5> ), .B(n49), .Y(n2048) );
  OAI21X1 U2120 ( .A(n1644), .B(n1658), .C(n2048), .Y(n2062) );
  NAND2X1 U2121 ( .A(\mem<0><6> ), .B(n48), .Y(n2049) );
  OAI21X1 U2122 ( .A(n1644), .B(n1660), .C(n2049), .Y(n2061) );
  NAND2X1 U2123 ( .A(\mem<0><7> ), .B(n48), .Y(n2050) );
  OAI21X1 U2124 ( .A(n1644), .B(n1662), .C(n2050), .Y(n2060) );
  OAI21X1 U2125 ( .A(n1644), .B(n1664), .C(n288), .Y(n2059) );
  OAI21X1 U2126 ( .A(n1644), .B(n1666), .C(n290), .Y(n2058) );
  OAI21X1 U2127 ( .A(n1644), .B(n1668), .C(n292), .Y(n2057) );
  OAI21X1 U2128 ( .A(n1644), .B(n1670), .C(n294), .Y(n2056) );
  OAI21X1 U2129 ( .A(n1644), .B(n1672), .C(n296), .Y(n2055) );
  OAI21X1 U2130 ( .A(n1644), .B(n1674), .C(n298), .Y(n2054) );
  NAND2X1 U2131 ( .A(\mem<0><14> ), .B(n48), .Y(n2051) );
  OAI21X1 U2132 ( .A(n1644), .B(n1676), .C(n2051), .Y(n2053) );
  OAI21X1 U2133 ( .A(n1644), .B(n1678), .C(n300), .Y(n2052) );
endmodule


module memc_Size16_4 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n112, n114, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n126, n128, n130, n132, n134, n136, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2223), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2224), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2225), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2226), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2227), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2228), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2229), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2230), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2231), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2232), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2233), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2234), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2235), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2236), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2237), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2238), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2239), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2240), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2241), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2242), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2243), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2244), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2245), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2246), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2247), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2248), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2249), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2250), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2251), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2252), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2253), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2254), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2255), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2256), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2257), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2258), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2259), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2260), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2261), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2262), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2263), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2264), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2265), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2266), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2267), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2268), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2269), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2270), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2271), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2272), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2273), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2274), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2275), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2276), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2277), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2278), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2279), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2280), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2281), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2282), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2283), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2284), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2285), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2286), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2287), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2288), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2289), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2290), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2291), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2292), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2293), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2294), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2295), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2296), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2297), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2298), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2299), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2300), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2301), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2302), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2303), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2304), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2305), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2306), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2307), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2308), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2309), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2310), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2311), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2312), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2313), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2314), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2315), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2316), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2317), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2318), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2319), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2320), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2321), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2322), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2323), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2324), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2325), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2326), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2327), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2328), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2329), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2330), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2331), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2332), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2333), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2334), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2335), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2336), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2337), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2338), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2339), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2340), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2341), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2342), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2343), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2344), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2345), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2346), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2347), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2348), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2349), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2350), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2351), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2352), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2353), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2354), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2355), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2356), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2357), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2358), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2359), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2360), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2361), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2362), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2363), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2364), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2365), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2366), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2367), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2368), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2369), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2370), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2371), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2372), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2373), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2374), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2375), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2376), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2377), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2378), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2379), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2380), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2381), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2382), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2383), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2384), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2385), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2386), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2387), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2388), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2389), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2390), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2391), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2392), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2393), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2394), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2395), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2396), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2397), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2398), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2399), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2400), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2401), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2402), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2403), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2404), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2405), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2406), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2407), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2408), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2409), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2410), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2411), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2412), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2413), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2414), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2415), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2416), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2417), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2418), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2419), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2420), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2421), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2422), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2423), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2424), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2425), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2426), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2427), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2428), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2429), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2430), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2431), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2432), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2433), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2434), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2435), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2436), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2437), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2438), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2439), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2440), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2441), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2442), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2443), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2444), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2445), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2446), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2447), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2448), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2449), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2450), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2451), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2452), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2453), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2454), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2455), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2456), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2457), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2458), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2459), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2460), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2461), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2462), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2463), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2464), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2465), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2466), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2467), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2468), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2469), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2470), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2471), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2472), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2473), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2474), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2475), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2476), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2477), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2478), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2479), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2480), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2481), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2482), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2483), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2484), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2485), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2486), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2487), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2488), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2489), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2490), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2491), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2492), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2493), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2494), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2495), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2496), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2497), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2498), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2499), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2500), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2501), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2502), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2503), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2504), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2505), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2506), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2507), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2508), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2509), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2510), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2511), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2512), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2513), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2514), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2515), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2516), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2517), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2518), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2519), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2520), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2521), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2522), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2523), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2524), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2525), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2526), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2527), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2528), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2529), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2530), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2531), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2532), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2533), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2534), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2535), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2536), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2537), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2538), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2539), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2540), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2541), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2542), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2543), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2544), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2545), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2546), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2547), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2548), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2549), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2550), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2551), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2552), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2553), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2554), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2555), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2556), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2557), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2558), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2559), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2560), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2561), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2562), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2563), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2564), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2565), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2566), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2567), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2568), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2569), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2570), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2571), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2572), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2573), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2574), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2575), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2576), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2577), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2578), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2579), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2580), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2581), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2582), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2583), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2584), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2585), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2586), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2587), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2588), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2589), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2590), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2591), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2592), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2593), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2594), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2595), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2596), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2597), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2598), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2599), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2600), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2601), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2602), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2603), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2604), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2605), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2606), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2607), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2608), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2609), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2610), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2611), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2612), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2613), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2614), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2615), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2616), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2617), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2618), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2619), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2620), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2621), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2622), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2623), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2624), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2625), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2626), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2627), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2628), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2629), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2630), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2631), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2632), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2633), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2634), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2635), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2636), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2637), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2638), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2639), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2640), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2641), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2642), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2643), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2644), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2645), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2646), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2647), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2648), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2649), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2650), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2651), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2652), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2653), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2654), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2655), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2656), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2657), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2658), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2659), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2660), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2661), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2662), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2663), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2664), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2665), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2666), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2667), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2668), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2669), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2670), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2671), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2672), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2673), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2674), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2675), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2676), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2677), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2678), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2679), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2680), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2681), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2682), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2683), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2684), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2685), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2686), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2687), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2688), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2689), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2690), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2691), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2692), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2693), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2694), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2695), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2696), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2697), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2698), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2699), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2700), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2701), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2702), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2703), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2704), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2705), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2706), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2707), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2708), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2709), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2710), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2711), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2712), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2713), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2714), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2715), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2716), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2717), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2718), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2719), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2720), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2721), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2722), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2723), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2724), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2725), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2726), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2727), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2728), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2729), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2730), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2731), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2732), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2733), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2734), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2735) );
  INVX1 U2 ( .A(write), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n33), .Y(n3) );
  AND2X2 U5 ( .A(n34), .B(n1216), .Y(\data_out<7> ) );
  INVX4 U6 ( .A(n185), .Y(n1916) );
  AND2X2 U7 ( .A(N25), .B(n1953), .Y(n1216) );
  INVX2 U8 ( .A(n1802), .Y(n1803) );
  INVX1 U9 ( .A(n1961), .Y(n1800) );
  INVX1 U10 ( .A(n1963), .Y(n1799) );
  INVX1 U11 ( .A(n1963), .Y(n1798) );
  INVX2 U12 ( .A(n1820), .Y(n1821) );
  INVX1 U13 ( .A(n1956), .Y(n1820) );
  INVX2 U14 ( .A(n1820), .Y(n1815) );
  INVX2 U15 ( .A(n1820), .Y(n1816) );
  INVX1 U16 ( .A(n1786), .Y(N28) );
  INVX1 U17 ( .A(n1789), .Y(N25) );
  INVX2 U18 ( .A(n1802), .Y(n1804) );
  INVX1 U19 ( .A(n1795), .Y(N19) );
  INVX1 U20 ( .A(n1797), .Y(N17) );
  INVX1 U21 ( .A(n1782), .Y(N32) );
  INVX1 U22 ( .A(n1783), .Y(N31) );
  INVX1 U23 ( .A(n1784), .Y(N30) );
  INVX1 U24 ( .A(n1785), .Y(N29) );
  INVX1 U25 ( .A(n1787), .Y(N27) );
  INVX1 U26 ( .A(n1788), .Y(N26) );
  INVX1 U27 ( .A(n1790), .Y(N24) );
  INVX1 U28 ( .A(n1792), .Y(N22) );
  INVX1 U29 ( .A(n1793), .Y(N21) );
  INVX1 U30 ( .A(n1794), .Y(N20) );
  INVX1 U31 ( .A(n1796), .Y(N18) );
  INVX1 U32 ( .A(n1791), .Y(N23) );
  INVX2 U33 ( .A(n196), .Y(n1935) );
  INVX2 U34 ( .A(n198), .Y(n1938) );
  BUFX2 U35 ( .A(n1247), .Y(n1851) );
  BUFX2 U36 ( .A(n1249), .Y(n1853) );
  BUFX2 U37 ( .A(n1251), .Y(n1856) );
  BUFX2 U38 ( .A(n1253), .Y(n1858) );
  BUFX2 U39 ( .A(n1255), .Y(n1860) );
  BUFX2 U40 ( .A(n1257), .Y(n1862) );
  BUFX2 U41 ( .A(n1259), .Y(n1864) );
  BUFX2 U42 ( .A(n1261), .Y(n1867) );
  BUFX2 U43 ( .A(n1263), .Y(n1869) );
  BUFX2 U44 ( .A(n1265), .Y(n1871) );
  BUFX2 U45 ( .A(n1267), .Y(n1873) );
  BUFX2 U46 ( .A(n1269), .Y(n1875) );
  BUFX2 U47 ( .A(n1271), .Y(n1877) );
  BUFX2 U48 ( .A(n1273), .Y(n1879) );
  BUFX2 U49 ( .A(n1275), .Y(n1882) );
  BUFX2 U50 ( .A(n1277), .Y(n1884) );
  BUFX2 U51 ( .A(n1279), .Y(n1886) );
  BUFX2 U52 ( .A(n1281), .Y(n1888) );
  BUFX2 U53 ( .A(n1283), .Y(n1890) );
  BUFX2 U54 ( .A(n1285), .Y(n1892) );
  BUFX2 U55 ( .A(n1287), .Y(n1894) );
  BUFX2 U56 ( .A(n1289), .Y(n1897) );
  BUFX2 U57 ( .A(n1291), .Y(n1899) );
  BUFX2 U58 ( .A(n1293), .Y(n1901) );
  BUFX2 U59 ( .A(n1295), .Y(n1903) );
  BUFX2 U60 ( .A(n1297), .Y(n1905) );
  BUFX2 U61 ( .A(n1299), .Y(n1907) );
  BUFX2 U62 ( .A(n1301), .Y(n1909) );
  INVX4 U63 ( .A(n1850), .Y(n1828) );
  INVX4 U64 ( .A(n1850), .Y(n1826) );
  INVX1 U65 ( .A(N12), .Y(n1959) );
  INVX2 U66 ( .A(n1954), .Y(n1849) );
  INVX2 U67 ( .A(n1961), .Y(n1801) );
  INVX2 U68 ( .A(n1959), .Y(n1805) );
  INVX2 U69 ( .A(n1959), .Y(n1806) );
  INVX1 U70 ( .A(rst), .Y(n1953) );
  INVX1 U71 ( .A(n1963), .Y(n1962) );
  INVX1 U72 ( .A(N14), .Y(n1963) );
  INVX1 U73 ( .A(n1958), .Y(n1802) );
  INVX4 U74 ( .A(n202), .Y(n1945) );
  INVX4 U75 ( .A(n202), .Y(n1946) );
  INVX1 U76 ( .A(n1244), .Y(n1896) );
  INVX1 U77 ( .A(n1245), .Y(n1911) );
  BUFX2 U78 ( .A(n1263), .Y(n1870) );
  BUFX2 U79 ( .A(n1265), .Y(n1872) );
  BUFX2 U80 ( .A(n1267), .Y(n1874) );
  BUFX2 U81 ( .A(n1269), .Y(n1876) );
  BUFX2 U82 ( .A(n1271), .Y(n1878) );
  BUFX2 U83 ( .A(n1273), .Y(n1880) );
  BUFX2 U84 ( .A(n1275), .Y(n1883) );
  BUFX2 U85 ( .A(n1277), .Y(n1885) );
  BUFX2 U86 ( .A(n1279), .Y(n1887) );
  BUFX2 U87 ( .A(n1281), .Y(n1889) );
  BUFX2 U88 ( .A(n1283), .Y(n1891) );
  BUFX2 U89 ( .A(n1285), .Y(n1893) );
  BUFX2 U90 ( .A(n1287), .Y(n1895) );
  INVX1 U91 ( .A(n1961), .Y(n1960) );
  INVX1 U92 ( .A(N13), .Y(n1961) );
  BUFX2 U93 ( .A(n1247), .Y(n1852) );
  BUFX2 U94 ( .A(n1289), .Y(n1898) );
  BUFX2 U95 ( .A(n1291), .Y(n1900) );
  BUFX2 U96 ( .A(n1293), .Y(n1902) );
  BUFX2 U97 ( .A(n1295), .Y(n1904) );
  BUFX2 U98 ( .A(n1297), .Y(n1906) );
  BUFX2 U99 ( .A(n1299), .Y(n1908) );
  BUFX2 U100 ( .A(n1301), .Y(n1910) );
  BUFX2 U101 ( .A(n1251), .Y(n1857) );
  BUFX2 U102 ( .A(n1253), .Y(n1859) );
  BUFX2 U103 ( .A(n1255), .Y(n1861) );
  BUFX2 U104 ( .A(n1257), .Y(n1863) );
  BUFX2 U105 ( .A(n1259), .Y(n1865) );
  BUFX2 U106 ( .A(n1261), .Y(n1868) );
  BUFX2 U107 ( .A(n1249), .Y(n1854) );
  INVX1 U108 ( .A(n1242), .Y(n1866) );
  INVX1 U109 ( .A(n1243), .Y(n1881) );
  INVX4 U110 ( .A(n202), .Y(n12) );
  INVX1 U111 ( .A(n195), .Y(n5) );
  INVX1 U112 ( .A(n1935), .Y(n1933) );
  INVX1 U113 ( .A(n197), .Y(n6) );
  INVX1 U114 ( .A(n1938), .Y(n16) );
  INVX1 U115 ( .A(n1935), .Y(n7) );
  INVX1 U116 ( .A(n1927), .Y(n8) );
  INVX1 U117 ( .A(n1930), .Y(n9) );
  INVX1 U118 ( .A(n1920), .Y(n10) );
  INVX1 U119 ( .A(n1938), .Y(n11) );
  INVX8 U120 ( .A(n1920), .Y(n13) );
  INVX8 U121 ( .A(n1927), .Y(n14) );
  INVX8 U122 ( .A(n1930), .Y(n15) );
  INVX8 U123 ( .A(n1935), .Y(n17) );
  INVX4 U124 ( .A(n1915), .Y(n1913) );
  INVX1 U125 ( .A(n34), .Y(n18) );
  INVX2 U126 ( .A(n157), .Y(n19) );
  INVX2 U127 ( .A(n151), .Y(n20) );
  INVX2 U128 ( .A(n148), .Y(n21) );
  INVX2 U129 ( .A(n145), .Y(n22) );
  INVX2 U130 ( .A(n142), .Y(n23) );
  INVX2 U131 ( .A(n139), .Y(n24) );
  INVX2 U132 ( .A(n154), .Y(n25) );
  INVX4 U133 ( .A(n108), .Y(n109) );
  INVX4 U134 ( .A(n180), .Y(n181) );
  INVX4 U135 ( .A(n178), .Y(n179) );
  INVX4 U136 ( .A(n176), .Y(n177) );
  INVX4 U137 ( .A(n174), .Y(n175) );
  INVX4 U138 ( .A(n172), .Y(n173) );
  INVX4 U139 ( .A(n170), .Y(n171) );
  INVX4 U140 ( .A(n168), .Y(n169) );
  INVX4 U141 ( .A(n164), .Y(n165) );
  INVX4 U142 ( .A(n162), .Y(n163) );
  INVX4 U143 ( .A(n160), .Y(n161) );
  INVX4 U144 ( .A(n166), .Y(n167) );
  INVX4 U145 ( .A(n106), .Y(n107) );
  INVX4 U146 ( .A(n104), .Y(n105) );
  INVX4 U147 ( .A(n102), .Y(n103) );
  AND2X2 U148 ( .A(n35), .B(n1224), .Y(\data_out<12> ) );
  AND2X2 U149 ( .A(n35), .B(n1215), .Y(\data_out<6> ) );
  AND2X2 U150 ( .A(n33), .B(n1227), .Y(\data_out<14> ) );
  AND2X2 U151 ( .A(n33), .B(n1219), .Y(\data_out<9> ) );
  INVX4 U152 ( .A(n100), .Y(n101) );
  INVX4 U153 ( .A(n98), .Y(n99) );
  INVX4 U154 ( .A(n96), .Y(n97) );
  INVX4 U155 ( .A(n94), .Y(n95) );
  INVX4 U156 ( .A(n92), .Y(n93) );
  INVX1 U157 ( .A(write), .Y(n30) );
  INVX1 U158 ( .A(n30), .Y(n31) );
  INVX1 U159 ( .A(n35), .Y(n32) );
  INVX1 U160 ( .A(write), .Y(n33) );
  INVX1 U161 ( .A(write), .Y(n34) );
  INVX1 U162 ( .A(write), .Y(n35) );
  AND2X2 U163 ( .A(\mem<31><1> ), .B(n117), .Y(n36) );
  INVX1 U164 ( .A(n36), .Y(n37) );
  AND2X2 U165 ( .A(\mem<31><2> ), .B(n117), .Y(n38) );
  INVX1 U166 ( .A(n38), .Y(n39) );
  AND2X2 U167 ( .A(\mem<31><3> ), .B(n117), .Y(n40) );
  INVX1 U168 ( .A(n40), .Y(n41) );
  AND2X2 U169 ( .A(\mem<31><4> ), .B(n117), .Y(n42) );
  INVX1 U170 ( .A(n42), .Y(n43) );
  AND2X2 U171 ( .A(\mem<31><5> ), .B(n117), .Y(n44) );
  INVX1 U172 ( .A(n44), .Y(n45) );
  AND2X2 U173 ( .A(\mem<31><6> ), .B(n117), .Y(n46) );
  INVX1 U174 ( .A(n46), .Y(n47) );
  AND2X2 U175 ( .A(\mem<31><7> ), .B(n117), .Y(n48) );
  INVX1 U176 ( .A(n48), .Y(n49) );
  AND2X2 U177 ( .A(\mem<22><8> ), .B(n119), .Y(n50) );
  INVX1 U178 ( .A(n50), .Y(n51) );
  AND2X2 U179 ( .A(\mem<22><9> ), .B(n119), .Y(n52) );
  INVX1 U180 ( .A(n52), .Y(n53) );
  AND2X2 U181 ( .A(\mem<22><10> ), .B(n119), .Y(n54) );
  INVX1 U182 ( .A(n54), .Y(n55) );
  AND2X2 U183 ( .A(\mem<22><11> ), .B(n119), .Y(n56) );
  INVX1 U184 ( .A(n56), .Y(n57) );
  AND2X2 U185 ( .A(\mem<22><12> ), .B(n119), .Y(n58) );
  INVX1 U186 ( .A(n58), .Y(n59) );
  AND2X2 U187 ( .A(\mem<22><13> ), .B(n119), .Y(n60) );
  INVX1 U188 ( .A(n60), .Y(n61) );
  AND2X2 U189 ( .A(\mem<22><14> ), .B(n119), .Y(n62) );
  INVX1 U190 ( .A(n62), .Y(n63) );
  AND2X2 U191 ( .A(\mem<21><8> ), .B(n121), .Y(n64) );
  INVX1 U192 ( .A(n64), .Y(n65) );
  AND2X2 U193 ( .A(\mem<21><9> ), .B(n121), .Y(n66) );
  INVX1 U194 ( .A(n66), .Y(n67) );
  AND2X2 U195 ( .A(\mem<21><10> ), .B(n121), .Y(n68) );
  INVX1 U196 ( .A(n68), .Y(n69) );
  AND2X2 U197 ( .A(\mem<21><11> ), .B(n121), .Y(n70) );
  INVX1 U198 ( .A(n70), .Y(n71) );
  AND2X2 U199 ( .A(\mem<21><12> ), .B(n121), .Y(n72) );
  INVX1 U200 ( .A(n72), .Y(n73) );
  AND2X2 U201 ( .A(\mem<21><13> ), .B(n121), .Y(n74) );
  INVX1 U202 ( .A(n74), .Y(n75) );
  AND2X2 U203 ( .A(\mem<21><14> ), .B(n121), .Y(n76) );
  INVX1 U204 ( .A(n76), .Y(n77) );
  AND2X2 U205 ( .A(\mem<20><8> ), .B(n123), .Y(n78) );
  INVX1 U206 ( .A(n78), .Y(n79) );
  AND2X2 U207 ( .A(\mem<20><9> ), .B(n123), .Y(n80) );
  INVX1 U208 ( .A(n80), .Y(n81) );
  AND2X2 U209 ( .A(\mem<20><10> ), .B(n123), .Y(n82) );
  INVX1 U210 ( .A(n82), .Y(n83) );
  AND2X2 U211 ( .A(\mem<20><11> ), .B(n123), .Y(n84) );
  INVX1 U212 ( .A(n84), .Y(n85) );
  AND2X2 U213 ( .A(\mem<20><12> ), .B(n123), .Y(n86) );
  INVX1 U214 ( .A(n86), .Y(n87) );
  AND2X2 U215 ( .A(\mem<20><13> ), .B(n123), .Y(n88) );
  INVX1 U216 ( .A(n88), .Y(n89) );
  AND2X2 U217 ( .A(\mem<20><14> ), .B(n123), .Y(n90) );
  INVX1 U218 ( .A(n90), .Y(n91) );
  INVX4 U219 ( .A(n118), .Y(n119) );
  INVX4 U220 ( .A(n120), .Y(n121) );
  INVX4 U221 ( .A(n122), .Y(n123) );
  INVX4 U222 ( .A(n116), .Y(n117) );
  AND2X2 U223 ( .A(n1913), .B(n1244), .Y(n92) );
  AND2X2 U224 ( .A(n1914), .B(n1288), .Y(n94) );
  AND2X2 U225 ( .A(n1912), .B(n1290), .Y(n96) );
  AND2X2 U226 ( .A(n1914), .B(n1292), .Y(n98) );
  AND2X2 U227 ( .A(n1912), .B(n1294), .Y(n100) );
  AND2X2 U228 ( .A(n1913), .B(n1296), .Y(n102) );
  AND2X2 U229 ( .A(n1914), .B(n1298), .Y(n104) );
  AND2X2 U230 ( .A(n1912), .B(n1300), .Y(n106) );
  AND2X2 U231 ( .A(n1914), .B(n1245), .Y(n108) );
  OR2X2 U232 ( .A(n2), .B(n1218), .Y(n110) );
  INVX1 U233 ( .A(n110), .Y(\data_out<8> ) );
  OR2X2 U234 ( .A(write), .B(n1221), .Y(n112) );
  INVX1 U235 ( .A(n112), .Y(\data_out<10> ) );
  OR2X2 U236 ( .A(n31), .B(n1229), .Y(n114) );
  INVX1 U237 ( .A(n114), .Y(\data_out<15> ) );
  AND2X2 U238 ( .A(n1914), .B(n1246), .Y(n116) );
  AND2X2 U239 ( .A(n1914), .B(n1262), .Y(n118) );
  AND2X2 U240 ( .A(n1912), .B(n1264), .Y(n120) );
  AND2X2 U241 ( .A(n1914), .B(n1266), .Y(n122) );
  OR2X2 U242 ( .A(write), .B(n1204), .Y(n124) );
  INVX1 U243 ( .A(n124), .Y(\data_out<0> ) );
  OR2X2 U244 ( .A(write), .B(n1206), .Y(n126) );
  INVX1 U245 ( .A(n126), .Y(\data_out<1> ) );
  OR2X2 U246 ( .A(n18), .B(n1208), .Y(n128) );
  INVX1 U247 ( .A(n128), .Y(\data_out<2> ) );
  OR2X2 U248 ( .A(write), .B(n1210), .Y(n130) );
  INVX1 U249 ( .A(n130), .Y(\data_out<3> ) );
  OR2X2 U250 ( .A(write), .B(n1214), .Y(n132) );
  INVX1 U251 ( .A(n132), .Y(\data_out<5> ) );
  OR2X2 U252 ( .A(write), .B(n1223), .Y(n134) );
  INVX1 U253 ( .A(n134), .Y(\data_out<11> ) );
  OR2X2 U254 ( .A(n32), .B(n1226), .Y(n136) );
  INVX1 U255 ( .A(n136), .Y(\data_out<13> ) );
  AND2X2 U256 ( .A(n3), .B(n1953), .Y(n138) );
  AND2X2 U257 ( .A(n1912), .B(n1250), .Y(n139) );
  INVX1 U258 ( .A(n139), .Y(n140) );
  INVX1 U259 ( .A(n139), .Y(n141) );
  AND2X2 U260 ( .A(n1914), .B(n1252), .Y(n142) );
  INVX1 U261 ( .A(n142), .Y(n143) );
  INVX1 U262 ( .A(n142), .Y(n144) );
  AND2X2 U263 ( .A(n1912), .B(n1254), .Y(n145) );
  INVX1 U264 ( .A(n145), .Y(n146) );
  INVX1 U265 ( .A(n145), .Y(n147) );
  AND2X2 U266 ( .A(n1914), .B(n1256), .Y(n148) );
  INVX1 U267 ( .A(n148), .Y(n149) );
  INVX1 U268 ( .A(n148), .Y(n150) );
  AND2X2 U269 ( .A(n1913), .B(n1258), .Y(n151) );
  INVX1 U270 ( .A(n151), .Y(n152) );
  INVX1 U271 ( .A(n151), .Y(n153) );
  AND2X2 U272 ( .A(n1914), .B(n1242), .Y(n154) );
  INVX1 U273 ( .A(n154), .Y(n155) );
  INVX1 U274 ( .A(n154), .Y(n156) );
  AND2X2 U275 ( .A(n1912), .B(n1260), .Y(n157) );
  INVX1 U276 ( .A(n157), .Y(n158) );
  INVX1 U277 ( .A(n157), .Y(n159) );
  AND2X2 U278 ( .A(n1912), .B(n1268), .Y(n160) );
  AND2X2 U279 ( .A(n1914), .B(n1270), .Y(n162) );
  AND2X2 U280 ( .A(n1912), .B(n1272), .Y(n164) );
  AND2X2 U281 ( .A(n1912), .B(n1243), .Y(n166) );
  AND2X2 U282 ( .A(n1912), .B(n1274), .Y(n168) );
  AND2X2 U283 ( .A(n1913), .B(n1276), .Y(n170) );
  AND2X2 U284 ( .A(n1912), .B(n1278), .Y(n172) );
  AND2X2 U285 ( .A(n1912), .B(n1280), .Y(n174) );
  AND2X2 U286 ( .A(n1914), .B(n1282), .Y(n176) );
  AND2X2 U287 ( .A(n1912), .B(n1284), .Y(n178) );
  AND2X2 U288 ( .A(n1912), .B(n1286), .Y(n180) );
  AND2X2 U289 ( .A(n1913), .B(n1248), .Y(n182) );
  INVX1 U290 ( .A(n182), .Y(n183) );
  INVX1 U291 ( .A(n182), .Y(n184) );
  AND2X2 U292 ( .A(\data_in<0> ), .B(n1912), .Y(n185) );
  AND2X2 U293 ( .A(\data_in<1> ), .B(n1914), .Y(n186) );
  INVX1 U294 ( .A(n186), .Y(n187) );
  AND2X2 U295 ( .A(\data_in<2> ), .B(n1914), .Y(n188) );
  AND2X2 U296 ( .A(\data_in<3> ), .B(n1914), .Y(n189) );
  AND2X2 U297 ( .A(\data_in<4> ), .B(n1914), .Y(n190) );
  INVX1 U298 ( .A(n190), .Y(n191) );
  AND2X2 U299 ( .A(\data_in<5> ), .B(n1914), .Y(n192) );
  INVX1 U300 ( .A(n192), .Y(n193) );
  AND2X2 U301 ( .A(\data_in<6> ), .B(n1914), .Y(n194) );
  AND2X2 U302 ( .A(\data_in<7> ), .B(n1914), .Y(n195) );
  INVX1 U303 ( .A(n195), .Y(n196) );
  AND2X2 U304 ( .A(\data_in<8> ), .B(n1914), .Y(n197) );
  INVX1 U305 ( .A(n197), .Y(n198) );
  AND2X2 U306 ( .A(\data_in<9> ), .B(n1914), .Y(n199) );
  AND2X2 U307 ( .A(\data_in<10> ), .B(n1912), .Y(n200) );
  AND2X2 U308 ( .A(\data_in<11> ), .B(n1913), .Y(n201) );
  AND2X2 U309 ( .A(\data_in<12> ), .B(n1913), .Y(n202) );
  AND2X2 U310 ( .A(\data_in<13> ), .B(n1913), .Y(n203) );
  AND2X2 U311 ( .A(\data_in<14> ), .B(n1913), .Y(n204) );
  AND2X2 U312 ( .A(\data_in<15> ), .B(n1914), .Y(n205) );
  OR2X2 U313 ( .A(write), .B(n1212), .Y(n206) );
  AND2X2 U314 ( .A(\mem<19><1> ), .B(n161), .Y(n207) );
  INVX1 U315 ( .A(n207), .Y(n208) );
  AND2X2 U316 ( .A(\mem<19><2> ), .B(n161), .Y(n209) );
  INVX1 U317 ( .A(n209), .Y(n210) );
  AND2X2 U318 ( .A(\mem<19><3> ), .B(n161), .Y(n211) );
  INVX1 U319 ( .A(n211), .Y(n212) );
  AND2X2 U320 ( .A(\mem<19><4> ), .B(n161), .Y(n213) );
  INVX1 U321 ( .A(n213), .Y(n215) );
  AND2X2 U322 ( .A(\mem<19><5> ), .B(n161), .Y(n216) );
  INVX1 U323 ( .A(n216), .Y(n217) );
  AND2X2 U324 ( .A(\mem<19><6> ), .B(n161), .Y(n218) );
  INVX1 U325 ( .A(n218), .Y(n219) );
  AND2X2 U326 ( .A(\mem<19><7> ), .B(n161), .Y(n220) );
  INVX1 U327 ( .A(n220), .Y(n221) );
  AND2X2 U328 ( .A(\mem<18><1> ), .B(n163), .Y(n222) );
  INVX1 U329 ( .A(n222), .Y(n223) );
  AND2X2 U330 ( .A(\mem<18><2> ), .B(n163), .Y(n224) );
  INVX1 U331 ( .A(n224), .Y(n225) );
  AND2X2 U332 ( .A(\mem<18><3> ), .B(n163), .Y(n226) );
  INVX1 U333 ( .A(n226), .Y(n227) );
  AND2X2 U334 ( .A(\mem<18><4> ), .B(n163), .Y(n228) );
  INVX1 U335 ( .A(n228), .Y(n229) );
  AND2X2 U336 ( .A(\mem<18><5> ), .B(n163), .Y(n230) );
  INVX1 U337 ( .A(n230), .Y(n231) );
  AND2X2 U338 ( .A(\mem<18><6> ), .B(n163), .Y(n232) );
  INVX1 U339 ( .A(n232), .Y(n233) );
  AND2X2 U340 ( .A(\mem<18><7> ), .B(n163), .Y(n234) );
  INVX1 U341 ( .A(n234), .Y(n235) );
  AND2X2 U342 ( .A(\mem<17><1> ), .B(n165), .Y(n236) );
  INVX1 U343 ( .A(n236), .Y(n237) );
  AND2X2 U344 ( .A(\mem<17><2> ), .B(n165), .Y(n238) );
  INVX1 U345 ( .A(n238), .Y(n239) );
  AND2X2 U346 ( .A(\mem<17><3> ), .B(n165), .Y(n240) );
  INVX1 U347 ( .A(n240), .Y(n241) );
  AND2X2 U348 ( .A(\mem<17><4> ), .B(n165), .Y(n242) );
  INVX1 U349 ( .A(n242), .Y(n243) );
  AND2X2 U350 ( .A(\mem<17><5> ), .B(n165), .Y(n244) );
  INVX1 U351 ( .A(n244), .Y(n245) );
  AND2X2 U352 ( .A(\mem<17><6> ), .B(n165), .Y(n246) );
  INVX1 U353 ( .A(n246), .Y(n247) );
  AND2X2 U354 ( .A(\mem<17><7> ), .B(n165), .Y(n248) );
  INVX1 U355 ( .A(n248), .Y(n249) );
  AND2X2 U356 ( .A(\mem<16><1> ), .B(n167), .Y(n250) );
  INVX1 U357 ( .A(n250), .Y(n251) );
  AND2X2 U358 ( .A(\mem<16><2> ), .B(n167), .Y(n252) );
  INVX1 U359 ( .A(n252), .Y(n253) );
  AND2X2 U360 ( .A(\mem<16><3> ), .B(n167), .Y(n254) );
  INVX1 U361 ( .A(n254), .Y(n255) );
  AND2X2 U362 ( .A(\mem<16><4> ), .B(n167), .Y(n256) );
  INVX1 U363 ( .A(n256), .Y(n257) );
  AND2X2 U364 ( .A(\mem<16><5> ), .B(n167), .Y(n258) );
  INVX1 U365 ( .A(n258), .Y(n259) );
  AND2X2 U366 ( .A(\mem<16><6> ), .B(n167), .Y(n260) );
  INVX1 U367 ( .A(n260), .Y(n261) );
  AND2X2 U368 ( .A(\mem<16><7> ), .B(n167), .Y(n262) );
  INVX1 U369 ( .A(n262), .Y(n263) );
  AND2X2 U370 ( .A(\mem<15><1> ), .B(n169), .Y(n264) );
  INVX1 U371 ( .A(n264), .Y(n265) );
  AND2X2 U372 ( .A(\mem<15><2> ), .B(n169), .Y(n266) );
  INVX1 U373 ( .A(n266), .Y(n267) );
  AND2X2 U374 ( .A(\mem<15><3> ), .B(n169), .Y(n268) );
  INVX1 U375 ( .A(n268), .Y(n269) );
  AND2X2 U376 ( .A(\mem<15><4> ), .B(n169), .Y(n270) );
  INVX1 U377 ( .A(n270), .Y(n271) );
  AND2X2 U378 ( .A(\mem<15><5> ), .B(n169), .Y(n272) );
  INVX1 U379 ( .A(n272), .Y(n273) );
  AND2X2 U380 ( .A(\mem<15><6> ), .B(n169), .Y(n274) );
  INVX1 U381 ( .A(n274), .Y(n275) );
  AND2X2 U382 ( .A(\mem<15><7> ), .B(n169), .Y(n276) );
  INVX1 U383 ( .A(n276), .Y(n277) );
  AND2X2 U384 ( .A(\mem<14><1> ), .B(n171), .Y(n278) );
  INVX1 U385 ( .A(n278), .Y(n279) );
  AND2X2 U386 ( .A(\mem<14><2> ), .B(n171), .Y(n280) );
  INVX1 U387 ( .A(n280), .Y(n281) );
  AND2X2 U388 ( .A(\mem<14><3> ), .B(n171), .Y(n282) );
  INVX1 U389 ( .A(n282), .Y(n283) );
  AND2X2 U390 ( .A(\mem<14><4> ), .B(n171), .Y(n284) );
  INVX1 U391 ( .A(n284), .Y(n285) );
  AND2X2 U392 ( .A(\mem<14><5> ), .B(n171), .Y(n286) );
  INVX1 U393 ( .A(n286), .Y(n287) );
  AND2X2 U394 ( .A(\mem<14><6> ), .B(n171), .Y(n288) );
  INVX1 U395 ( .A(n288), .Y(n289) );
  AND2X2 U396 ( .A(\mem<14><7> ), .B(n171), .Y(n290) );
  INVX1 U397 ( .A(n290), .Y(n291) );
  AND2X2 U398 ( .A(\mem<13><1> ), .B(n173), .Y(n292) );
  INVX1 U399 ( .A(n292), .Y(n293) );
  AND2X2 U400 ( .A(\mem<13><2> ), .B(n173), .Y(n294) );
  INVX1 U401 ( .A(n294), .Y(n295) );
  AND2X2 U402 ( .A(\mem<13><3> ), .B(n173), .Y(n296) );
  INVX1 U403 ( .A(n296), .Y(n297) );
  AND2X2 U404 ( .A(\mem<13><4> ), .B(n173), .Y(n298) );
  INVX1 U405 ( .A(n298), .Y(n299) );
  AND2X2 U406 ( .A(\mem<13><5> ), .B(n173), .Y(n300) );
  INVX1 U407 ( .A(n300), .Y(n301) );
  AND2X2 U408 ( .A(\mem<13><6> ), .B(n173), .Y(n302) );
  INVX1 U409 ( .A(n302), .Y(n303) );
  AND2X2 U410 ( .A(\mem<13><7> ), .B(n173), .Y(n304) );
  INVX1 U411 ( .A(n304), .Y(n305) );
  AND2X2 U412 ( .A(\mem<12><1> ), .B(n175), .Y(n306) );
  INVX1 U413 ( .A(n306), .Y(n307) );
  AND2X2 U414 ( .A(\mem<12><2> ), .B(n175), .Y(n308) );
  INVX1 U415 ( .A(n308), .Y(n309) );
  AND2X2 U416 ( .A(\mem<12><3> ), .B(n175), .Y(n310) );
  INVX1 U417 ( .A(n310), .Y(n311) );
  AND2X2 U418 ( .A(\mem<12><4> ), .B(n175), .Y(n312) );
  INVX1 U419 ( .A(n312), .Y(n313) );
  AND2X2 U420 ( .A(\mem<12><5> ), .B(n175), .Y(n314) );
  INVX1 U421 ( .A(n314), .Y(n315) );
  AND2X2 U422 ( .A(\mem<12><6> ), .B(n175), .Y(n316) );
  INVX1 U423 ( .A(n316), .Y(n317) );
  AND2X2 U424 ( .A(\mem<12><7> ), .B(n175), .Y(n318) );
  INVX1 U425 ( .A(n318), .Y(n319) );
  AND2X2 U426 ( .A(\mem<11><1> ), .B(n177), .Y(n320) );
  INVX1 U427 ( .A(n320), .Y(n321) );
  AND2X2 U428 ( .A(\mem<11><2> ), .B(n177), .Y(n322) );
  INVX1 U429 ( .A(n322), .Y(n323) );
  AND2X2 U430 ( .A(\mem<11><3> ), .B(n177), .Y(n324) );
  INVX1 U431 ( .A(n324), .Y(n325) );
  AND2X2 U432 ( .A(\mem<11><4> ), .B(n177), .Y(n326) );
  INVX1 U433 ( .A(n326), .Y(n327) );
  AND2X2 U434 ( .A(\mem<11><5> ), .B(n177), .Y(n328) );
  INVX1 U435 ( .A(n328), .Y(n329) );
  AND2X2 U436 ( .A(\mem<11><6> ), .B(n177), .Y(n330) );
  INVX1 U437 ( .A(n330), .Y(n331) );
  AND2X2 U438 ( .A(\mem<11><7> ), .B(n177), .Y(n332) );
  INVX1 U439 ( .A(n332), .Y(n333) );
  AND2X2 U440 ( .A(\mem<10><1> ), .B(n179), .Y(n334) );
  INVX1 U441 ( .A(n334), .Y(n335) );
  AND2X2 U442 ( .A(\mem<10><2> ), .B(n179), .Y(n336) );
  INVX1 U443 ( .A(n336), .Y(n337) );
  AND2X2 U444 ( .A(\mem<10><3> ), .B(n179), .Y(n338) );
  INVX1 U445 ( .A(n338), .Y(n339) );
  AND2X2 U446 ( .A(\mem<10><4> ), .B(n179), .Y(n340) );
  INVX1 U447 ( .A(n340), .Y(n341) );
  AND2X2 U448 ( .A(\mem<10><5> ), .B(n179), .Y(n342) );
  INVX1 U449 ( .A(n342), .Y(n343) );
  AND2X2 U450 ( .A(\mem<10><6> ), .B(n179), .Y(n344) );
  INVX1 U451 ( .A(n344), .Y(n345) );
  AND2X2 U452 ( .A(\mem<10><7> ), .B(n179), .Y(n346) );
  INVX1 U453 ( .A(n346), .Y(n347) );
  AND2X2 U454 ( .A(\mem<9><1> ), .B(n181), .Y(n348) );
  INVX1 U455 ( .A(n348), .Y(n349) );
  AND2X2 U456 ( .A(\mem<9><2> ), .B(n181), .Y(n350) );
  INVX1 U457 ( .A(n350), .Y(n351) );
  AND2X2 U458 ( .A(\mem<9><3> ), .B(n181), .Y(n352) );
  INVX1 U459 ( .A(n352), .Y(n353) );
  AND2X2 U460 ( .A(\mem<9><4> ), .B(n181), .Y(n354) );
  INVX1 U461 ( .A(n354), .Y(n355) );
  AND2X2 U462 ( .A(\mem<9><5> ), .B(n181), .Y(n356) );
  INVX1 U463 ( .A(n356), .Y(n357) );
  AND2X2 U464 ( .A(\mem<9><6> ), .B(n181), .Y(n358) );
  INVX1 U465 ( .A(n358), .Y(n359) );
  AND2X2 U466 ( .A(\mem<9><7> ), .B(n181), .Y(n360) );
  INVX1 U467 ( .A(n360), .Y(n361) );
  AND2X2 U468 ( .A(\mem<8><8> ), .B(n93), .Y(n362) );
  INVX1 U469 ( .A(n362), .Y(n363) );
  AND2X2 U470 ( .A(\mem<8><9> ), .B(n93), .Y(n364) );
  INVX1 U471 ( .A(n364), .Y(n365) );
  AND2X2 U472 ( .A(\mem<8><10> ), .B(n93), .Y(n366) );
  INVX1 U473 ( .A(n366), .Y(n367) );
  AND2X2 U474 ( .A(\mem<8><11> ), .B(n93), .Y(n368) );
  INVX1 U475 ( .A(n368), .Y(n369) );
  AND2X2 U476 ( .A(\mem<8><12> ), .B(n93), .Y(n370) );
  INVX1 U477 ( .A(n370), .Y(n371) );
  AND2X2 U478 ( .A(\mem<8><13> ), .B(n93), .Y(n372) );
  INVX1 U479 ( .A(n372), .Y(n373) );
  AND2X2 U480 ( .A(\mem<8><14> ), .B(n93), .Y(n374) );
  INVX1 U481 ( .A(n374), .Y(n375) );
  AND2X2 U482 ( .A(\mem<8><15> ), .B(n93), .Y(n376) );
  INVX1 U483 ( .A(n376), .Y(n377) );
  AND2X2 U484 ( .A(\mem<7><8> ), .B(n95), .Y(n378) );
  INVX1 U485 ( .A(n378), .Y(n379) );
  AND2X2 U486 ( .A(\mem<7><9> ), .B(n95), .Y(n380) );
  INVX1 U487 ( .A(n380), .Y(n381) );
  AND2X2 U488 ( .A(\mem<7><10> ), .B(n95), .Y(n382) );
  INVX1 U489 ( .A(n382), .Y(n383) );
  AND2X2 U490 ( .A(\mem<7><11> ), .B(n95), .Y(n384) );
  INVX1 U491 ( .A(n384), .Y(n385) );
  AND2X2 U492 ( .A(\mem<7><12> ), .B(n95), .Y(n386) );
  INVX1 U493 ( .A(n386), .Y(n387) );
  AND2X2 U494 ( .A(\mem<7><13> ), .B(n95), .Y(n388) );
  INVX1 U495 ( .A(n388), .Y(n389) );
  AND2X2 U496 ( .A(\mem<7><14> ), .B(n95), .Y(n390) );
  INVX1 U497 ( .A(n390), .Y(n391) );
  AND2X2 U498 ( .A(\mem<7><15> ), .B(n95), .Y(n392) );
  INVX1 U499 ( .A(n392), .Y(n393) );
  AND2X2 U500 ( .A(\mem<6><8> ), .B(n97), .Y(n394) );
  INVX1 U501 ( .A(n394), .Y(n395) );
  AND2X2 U502 ( .A(\mem<6><9> ), .B(n97), .Y(n396) );
  INVX1 U503 ( .A(n396), .Y(n397) );
  AND2X2 U504 ( .A(\mem<6><10> ), .B(n97), .Y(n398) );
  INVX1 U505 ( .A(n398), .Y(n399) );
  AND2X2 U506 ( .A(\mem<6><11> ), .B(n97), .Y(n400) );
  INVX1 U507 ( .A(n400), .Y(n401) );
  AND2X2 U508 ( .A(\mem<6><12> ), .B(n97), .Y(n402) );
  INVX1 U509 ( .A(n402), .Y(n403) );
  AND2X2 U510 ( .A(\mem<6><13> ), .B(n97), .Y(n404) );
  INVX1 U511 ( .A(n404), .Y(n405) );
  AND2X2 U512 ( .A(\mem<6><14> ), .B(n97), .Y(n406) );
  INVX1 U513 ( .A(n406), .Y(n407) );
  AND2X2 U514 ( .A(\mem<6><15> ), .B(n97), .Y(n408) );
  INVX1 U515 ( .A(n408), .Y(n409) );
  AND2X2 U516 ( .A(\mem<5><8> ), .B(n99), .Y(n410) );
  INVX1 U517 ( .A(n410), .Y(n411) );
  AND2X2 U518 ( .A(\mem<5><9> ), .B(n99), .Y(n412) );
  INVX1 U519 ( .A(n412), .Y(n413) );
  AND2X2 U520 ( .A(\mem<5><10> ), .B(n99), .Y(n414) );
  INVX1 U521 ( .A(n414), .Y(n415) );
  AND2X2 U522 ( .A(\mem<5><11> ), .B(n99), .Y(n416) );
  INVX1 U523 ( .A(n416), .Y(n417) );
  AND2X2 U524 ( .A(\mem<5><12> ), .B(n99), .Y(n418) );
  INVX1 U525 ( .A(n418), .Y(n419) );
  AND2X2 U526 ( .A(\mem<5><13> ), .B(n99), .Y(n420) );
  INVX1 U527 ( .A(n420), .Y(n421) );
  AND2X2 U528 ( .A(\mem<5><14> ), .B(n99), .Y(n422) );
  INVX1 U529 ( .A(n422), .Y(n423) );
  AND2X2 U530 ( .A(\mem<5><15> ), .B(n99), .Y(n424) );
  INVX1 U531 ( .A(n424), .Y(n425) );
  AND2X2 U532 ( .A(\mem<4><8> ), .B(n101), .Y(n426) );
  INVX1 U533 ( .A(n426), .Y(n427) );
  AND2X2 U534 ( .A(\mem<4><9> ), .B(n101), .Y(n428) );
  INVX1 U535 ( .A(n428), .Y(n429) );
  AND2X2 U536 ( .A(\mem<4><10> ), .B(n101), .Y(n430) );
  INVX1 U537 ( .A(n430), .Y(n431) );
  AND2X2 U538 ( .A(\mem<4><11> ), .B(n101), .Y(n432) );
  INVX1 U539 ( .A(n432), .Y(n433) );
  AND2X2 U540 ( .A(\mem<4><12> ), .B(n101), .Y(n434) );
  INVX1 U541 ( .A(n434), .Y(n435) );
  AND2X2 U542 ( .A(\mem<4><13> ), .B(n101), .Y(n436) );
  INVX1 U543 ( .A(n436), .Y(n437) );
  AND2X2 U544 ( .A(\mem<4><14> ), .B(n101), .Y(n438) );
  INVX1 U545 ( .A(n438), .Y(n439) );
  AND2X2 U546 ( .A(\mem<4><15> ), .B(n101), .Y(n440) );
  INVX1 U547 ( .A(n440), .Y(n441) );
  AND2X2 U548 ( .A(\mem<3><8> ), .B(n103), .Y(n442) );
  INVX1 U549 ( .A(n442), .Y(n443) );
  AND2X2 U550 ( .A(\mem<3><9> ), .B(n103), .Y(n444) );
  INVX1 U551 ( .A(n444), .Y(n445) );
  AND2X2 U552 ( .A(\mem<3><10> ), .B(n103), .Y(n446) );
  INVX1 U553 ( .A(n446), .Y(n447) );
  AND2X2 U554 ( .A(\mem<3><11> ), .B(n103), .Y(n448) );
  INVX1 U555 ( .A(n448), .Y(n449) );
  AND2X2 U556 ( .A(\mem<3><12> ), .B(n103), .Y(n450) );
  INVX1 U557 ( .A(n450), .Y(n451) );
  AND2X2 U558 ( .A(\mem<3><13> ), .B(n103), .Y(n452) );
  INVX1 U559 ( .A(n452), .Y(n453) );
  AND2X2 U560 ( .A(\mem<3><14> ), .B(n103), .Y(n454) );
  INVX1 U561 ( .A(n454), .Y(n455) );
  AND2X2 U562 ( .A(\mem<3><15> ), .B(n103), .Y(n456) );
  INVX1 U563 ( .A(n456), .Y(n457) );
  AND2X2 U564 ( .A(\mem<2><8> ), .B(n105), .Y(n458) );
  INVX1 U565 ( .A(n458), .Y(n459) );
  AND2X2 U566 ( .A(\mem<2><9> ), .B(n105), .Y(n460) );
  INVX1 U567 ( .A(n460), .Y(n461) );
  AND2X2 U568 ( .A(\mem<2><10> ), .B(n105), .Y(n462) );
  INVX1 U569 ( .A(n462), .Y(n463) );
  AND2X2 U570 ( .A(\mem<2><11> ), .B(n105), .Y(n464) );
  INVX1 U571 ( .A(n464), .Y(n465) );
  AND2X2 U572 ( .A(\mem<2><12> ), .B(n105), .Y(n466) );
  INVX1 U573 ( .A(n466), .Y(n467) );
  AND2X2 U574 ( .A(\mem<2><13> ), .B(n105), .Y(n468) );
  INVX1 U575 ( .A(n468), .Y(n469) );
  AND2X2 U576 ( .A(\mem<2><14> ), .B(n105), .Y(n470) );
  INVX1 U577 ( .A(n470), .Y(n471) );
  AND2X2 U578 ( .A(\mem<2><15> ), .B(n105), .Y(n472) );
  INVX1 U579 ( .A(n472), .Y(n473) );
  AND2X2 U580 ( .A(\mem<1><8> ), .B(n107), .Y(n474) );
  INVX1 U581 ( .A(n474), .Y(n475) );
  AND2X2 U582 ( .A(\mem<1><9> ), .B(n107), .Y(n476) );
  INVX1 U583 ( .A(n476), .Y(n477) );
  AND2X2 U584 ( .A(\mem<1><10> ), .B(n107), .Y(n478) );
  INVX1 U585 ( .A(n478), .Y(n479) );
  AND2X2 U586 ( .A(\mem<1><11> ), .B(n107), .Y(n480) );
  INVX1 U587 ( .A(n480), .Y(n481) );
  AND2X2 U588 ( .A(\mem<1><12> ), .B(n107), .Y(n482) );
  INVX1 U589 ( .A(n482), .Y(n483) );
  AND2X2 U590 ( .A(\mem<1><13> ), .B(n107), .Y(n484) );
  INVX1 U591 ( .A(n484), .Y(n485) );
  AND2X2 U592 ( .A(\mem<1><14> ), .B(n107), .Y(n486) );
  INVX1 U593 ( .A(n486), .Y(n487) );
  AND2X2 U594 ( .A(\mem<1><15> ), .B(n107), .Y(n488) );
  INVX1 U595 ( .A(n488), .Y(n489) );
  BUFX2 U596 ( .A(n184), .Y(n490) );
  INVX1 U597 ( .A(n1959), .Y(n1958) );
  INVX1 U598 ( .A(n1955), .Y(n1954) );
  AND2X1 U599 ( .A(n1958), .B(n1956), .Y(n491) );
  INVX1 U600 ( .A(n1957), .Y(n1956) );
  AND2X1 U601 ( .A(n2735), .B(n1962), .Y(n492) );
  AND2X2 U602 ( .A(\mem<19><0> ), .B(n161), .Y(n493) );
  INVX1 U603 ( .A(n493), .Y(n494) );
  AND2X2 U604 ( .A(\mem<19><8> ), .B(n161), .Y(n495) );
  INVX1 U605 ( .A(n495), .Y(n496) );
  AND2X2 U606 ( .A(\mem<19><9> ), .B(n161), .Y(n497) );
  INVX1 U607 ( .A(n497), .Y(n498) );
  AND2X2 U608 ( .A(\mem<19><10> ), .B(n161), .Y(n499) );
  INVX1 U609 ( .A(n499), .Y(n500) );
  AND2X2 U610 ( .A(\mem<19><11> ), .B(n161), .Y(n501) );
  INVX1 U611 ( .A(n501), .Y(n502) );
  AND2X2 U612 ( .A(\mem<19><12> ), .B(n161), .Y(n503) );
  INVX1 U613 ( .A(n503), .Y(n504) );
  AND2X2 U614 ( .A(\mem<19><13> ), .B(n161), .Y(n505) );
  INVX1 U615 ( .A(n505), .Y(n506) );
  AND2X2 U616 ( .A(\mem<19><14> ), .B(n161), .Y(n507) );
  INVX1 U617 ( .A(n507), .Y(n508) );
  AND2X2 U618 ( .A(\mem<19><15> ), .B(n161), .Y(n509) );
  INVX1 U619 ( .A(n509), .Y(n510) );
  AND2X2 U620 ( .A(\mem<18><0> ), .B(n163), .Y(n511) );
  INVX1 U621 ( .A(n511), .Y(n512) );
  AND2X2 U622 ( .A(\mem<18><8> ), .B(n163), .Y(n513) );
  INVX1 U623 ( .A(n513), .Y(n514) );
  AND2X2 U624 ( .A(\mem<18><9> ), .B(n163), .Y(n515) );
  INVX1 U625 ( .A(n515), .Y(n516) );
  AND2X2 U626 ( .A(\mem<18><10> ), .B(n163), .Y(n517) );
  INVX1 U627 ( .A(n517), .Y(n518) );
  AND2X2 U628 ( .A(\mem<18><11> ), .B(n163), .Y(n519) );
  INVX1 U629 ( .A(n519), .Y(n520) );
  AND2X2 U630 ( .A(\mem<18><12> ), .B(n163), .Y(n521) );
  INVX1 U631 ( .A(n521), .Y(n522) );
  AND2X2 U632 ( .A(\mem<18><13> ), .B(n163), .Y(n523) );
  INVX1 U633 ( .A(n523), .Y(n524) );
  AND2X2 U634 ( .A(\mem<18><14> ), .B(n163), .Y(n525) );
  INVX1 U635 ( .A(n525), .Y(n526) );
  AND2X2 U636 ( .A(\mem<18><15> ), .B(n163), .Y(n527) );
  INVX1 U637 ( .A(n527), .Y(n528) );
  AND2X2 U638 ( .A(\mem<17><0> ), .B(n165), .Y(n529) );
  INVX1 U639 ( .A(n529), .Y(n530) );
  AND2X2 U640 ( .A(\mem<17><8> ), .B(n165), .Y(n531) );
  INVX1 U641 ( .A(n531), .Y(n532) );
  AND2X2 U642 ( .A(\mem<17><9> ), .B(n165), .Y(n533) );
  INVX1 U643 ( .A(n533), .Y(n534) );
  AND2X2 U644 ( .A(\mem<17><10> ), .B(n165), .Y(n535) );
  INVX1 U645 ( .A(n535), .Y(n536) );
  AND2X2 U646 ( .A(\mem<17><11> ), .B(n165), .Y(n537) );
  INVX1 U647 ( .A(n537), .Y(n538) );
  AND2X2 U648 ( .A(\mem<17><12> ), .B(n165), .Y(n539) );
  INVX1 U649 ( .A(n539), .Y(n540) );
  AND2X2 U650 ( .A(\mem<17><13> ), .B(n165), .Y(n541) );
  INVX1 U651 ( .A(n541), .Y(n542) );
  AND2X2 U652 ( .A(\mem<17><14> ), .B(n165), .Y(n543) );
  INVX1 U653 ( .A(n543), .Y(n544) );
  AND2X2 U654 ( .A(\mem<17><15> ), .B(n165), .Y(n545) );
  INVX1 U655 ( .A(n545), .Y(n546) );
  AND2X2 U656 ( .A(\mem<16><0> ), .B(n167), .Y(n547) );
  INVX1 U657 ( .A(n547), .Y(n548) );
  AND2X2 U658 ( .A(\mem<16><8> ), .B(n167), .Y(n549) );
  INVX1 U659 ( .A(n549), .Y(n550) );
  AND2X2 U660 ( .A(\mem<16><9> ), .B(n167), .Y(n551) );
  INVX1 U661 ( .A(n551), .Y(n552) );
  AND2X2 U662 ( .A(\mem<16><10> ), .B(n167), .Y(n553) );
  INVX1 U663 ( .A(n553), .Y(n554) );
  AND2X2 U664 ( .A(\mem<16><11> ), .B(n167), .Y(n555) );
  INVX1 U665 ( .A(n555), .Y(n556) );
  AND2X2 U666 ( .A(\mem<16><12> ), .B(n167), .Y(n557) );
  INVX1 U667 ( .A(n557), .Y(n558) );
  AND2X2 U668 ( .A(\mem<16><13> ), .B(n167), .Y(n559) );
  INVX1 U669 ( .A(n559), .Y(n560) );
  AND2X2 U670 ( .A(\mem<16><14> ), .B(n167), .Y(n561) );
  INVX1 U671 ( .A(n561), .Y(n562) );
  AND2X2 U672 ( .A(\mem<16><15> ), .B(n167), .Y(n563) );
  INVX1 U673 ( .A(n563), .Y(n564) );
  AND2X2 U674 ( .A(\mem<15><0> ), .B(n169), .Y(n565) );
  INVX1 U675 ( .A(n565), .Y(n566) );
  AND2X2 U676 ( .A(\mem<15><8> ), .B(n169), .Y(n567) );
  INVX1 U677 ( .A(n567), .Y(n568) );
  AND2X2 U678 ( .A(\mem<15><9> ), .B(n169), .Y(n569) );
  INVX1 U679 ( .A(n569), .Y(n570) );
  AND2X2 U680 ( .A(\mem<15><10> ), .B(n169), .Y(n571) );
  INVX1 U681 ( .A(n571), .Y(n572) );
  AND2X2 U682 ( .A(\mem<15><11> ), .B(n169), .Y(n573) );
  INVX1 U683 ( .A(n573), .Y(n574) );
  AND2X2 U684 ( .A(\mem<15><12> ), .B(n169), .Y(n575) );
  INVX1 U685 ( .A(n575), .Y(n576) );
  AND2X2 U686 ( .A(\mem<15><13> ), .B(n169), .Y(n577) );
  INVX1 U687 ( .A(n577), .Y(n578) );
  AND2X2 U688 ( .A(\mem<15><14> ), .B(n169), .Y(n579) );
  INVX1 U689 ( .A(n579), .Y(n580) );
  AND2X2 U690 ( .A(\mem<15><15> ), .B(n169), .Y(n581) );
  INVX1 U691 ( .A(n581), .Y(n582) );
  AND2X2 U692 ( .A(\mem<14><0> ), .B(n171), .Y(n583) );
  INVX1 U693 ( .A(n583), .Y(n584) );
  AND2X2 U694 ( .A(\mem<14><8> ), .B(n171), .Y(n585) );
  INVX1 U695 ( .A(n585), .Y(n586) );
  AND2X2 U696 ( .A(\mem<14><9> ), .B(n171), .Y(n587) );
  INVX1 U697 ( .A(n587), .Y(n588) );
  AND2X2 U698 ( .A(\mem<14><10> ), .B(n171), .Y(n589) );
  INVX1 U699 ( .A(n589), .Y(n590) );
  AND2X2 U700 ( .A(\mem<14><11> ), .B(n171), .Y(n591) );
  INVX1 U701 ( .A(n591), .Y(n592) );
  AND2X2 U702 ( .A(\mem<14><12> ), .B(n171), .Y(n593) );
  INVX1 U703 ( .A(n593), .Y(n594) );
  AND2X2 U704 ( .A(\mem<14><13> ), .B(n171), .Y(n595) );
  INVX1 U705 ( .A(n595), .Y(n596) );
  AND2X2 U706 ( .A(\mem<14><14> ), .B(n171), .Y(n597) );
  INVX1 U707 ( .A(n597), .Y(n598) );
  AND2X2 U708 ( .A(\mem<14><15> ), .B(n171), .Y(n599) );
  INVX1 U709 ( .A(n599), .Y(n600) );
  AND2X2 U710 ( .A(\mem<13><0> ), .B(n173), .Y(n601) );
  INVX1 U711 ( .A(n601), .Y(n602) );
  AND2X2 U712 ( .A(\mem<13><8> ), .B(n173), .Y(n603) );
  INVX1 U713 ( .A(n603), .Y(n604) );
  AND2X2 U714 ( .A(\mem<13><9> ), .B(n173), .Y(n605) );
  INVX1 U715 ( .A(n605), .Y(n606) );
  AND2X2 U716 ( .A(\mem<13><10> ), .B(n173), .Y(n607) );
  INVX1 U717 ( .A(n607), .Y(n608) );
  AND2X2 U718 ( .A(\mem<13><11> ), .B(n173), .Y(n609) );
  INVX1 U719 ( .A(n609), .Y(n610) );
  AND2X2 U720 ( .A(\mem<13><12> ), .B(n173), .Y(n611) );
  INVX1 U721 ( .A(n611), .Y(n612) );
  AND2X2 U722 ( .A(\mem<13><13> ), .B(n173), .Y(n613) );
  INVX1 U723 ( .A(n613), .Y(n614) );
  AND2X2 U724 ( .A(\mem<13><14> ), .B(n173), .Y(n615) );
  INVX1 U725 ( .A(n615), .Y(n616) );
  AND2X2 U726 ( .A(\mem<13><15> ), .B(n173), .Y(n617) );
  INVX1 U727 ( .A(n617), .Y(n618) );
  AND2X2 U728 ( .A(\mem<12><0> ), .B(n175), .Y(n619) );
  INVX1 U729 ( .A(n619), .Y(n620) );
  AND2X2 U730 ( .A(\mem<12><8> ), .B(n175), .Y(n621) );
  INVX1 U731 ( .A(n621), .Y(n622) );
  AND2X2 U732 ( .A(\mem<12><9> ), .B(n175), .Y(n623) );
  INVX1 U733 ( .A(n623), .Y(n624) );
  AND2X2 U734 ( .A(\mem<12><10> ), .B(n175), .Y(n625) );
  INVX1 U735 ( .A(n625), .Y(n626) );
  AND2X2 U736 ( .A(\mem<12><11> ), .B(n175), .Y(n627) );
  INVX1 U737 ( .A(n627), .Y(n628) );
  AND2X2 U738 ( .A(\mem<12><12> ), .B(n175), .Y(n629) );
  INVX1 U739 ( .A(n629), .Y(n630) );
  AND2X2 U740 ( .A(\mem<12><13> ), .B(n175), .Y(n631) );
  INVX1 U741 ( .A(n631), .Y(n632) );
  AND2X2 U742 ( .A(\mem<12><14> ), .B(n175), .Y(n633) );
  INVX1 U743 ( .A(n633), .Y(n634) );
  AND2X2 U744 ( .A(\mem<12><15> ), .B(n175), .Y(n635) );
  INVX1 U745 ( .A(n635), .Y(n636) );
  AND2X2 U746 ( .A(\mem<11><0> ), .B(n177), .Y(n637) );
  INVX1 U747 ( .A(n637), .Y(n638) );
  AND2X2 U748 ( .A(\mem<11><8> ), .B(n177), .Y(n639) );
  INVX1 U749 ( .A(n639), .Y(n640) );
  AND2X2 U750 ( .A(\mem<11><9> ), .B(n177), .Y(n641) );
  INVX1 U751 ( .A(n641), .Y(n642) );
  AND2X2 U752 ( .A(\mem<11><10> ), .B(n177), .Y(n643) );
  INVX1 U753 ( .A(n643), .Y(n644) );
  AND2X2 U754 ( .A(\mem<11><11> ), .B(n177), .Y(n645) );
  INVX1 U755 ( .A(n645), .Y(n646) );
  AND2X2 U756 ( .A(\mem<11><12> ), .B(n177), .Y(n647) );
  INVX1 U757 ( .A(n647), .Y(n648) );
  AND2X2 U758 ( .A(\mem<11><13> ), .B(n177), .Y(n649) );
  INVX1 U759 ( .A(n649), .Y(n650) );
  AND2X2 U760 ( .A(\mem<11><14> ), .B(n177), .Y(n1163) );
  INVX1 U761 ( .A(n1163), .Y(n1164) );
  AND2X2 U762 ( .A(\mem<11><15> ), .B(n177), .Y(n1165) );
  INVX1 U763 ( .A(n1165), .Y(n1166) );
  AND2X2 U764 ( .A(\mem<10><0> ), .B(n179), .Y(n1167) );
  INVX1 U765 ( .A(n1167), .Y(n1168) );
  AND2X2 U766 ( .A(\mem<10><8> ), .B(n179), .Y(n1169) );
  INVX1 U767 ( .A(n1169), .Y(n1170) );
  AND2X2 U768 ( .A(\mem<10><9> ), .B(n179), .Y(n1171) );
  INVX1 U769 ( .A(n1171), .Y(n1172) );
  AND2X2 U770 ( .A(\mem<10><10> ), .B(n179), .Y(n1173) );
  INVX1 U771 ( .A(n1173), .Y(n1174) );
  AND2X2 U772 ( .A(\mem<10><11> ), .B(n179), .Y(n1175) );
  INVX1 U773 ( .A(n1175), .Y(n1176) );
  AND2X2 U774 ( .A(\mem<10><12> ), .B(n179), .Y(n1177) );
  INVX1 U775 ( .A(n1177), .Y(n1178) );
  AND2X2 U776 ( .A(\mem<10><13> ), .B(n179), .Y(n1179) );
  INVX1 U777 ( .A(n1179), .Y(n1180) );
  AND2X2 U778 ( .A(\mem<10><14> ), .B(n179), .Y(n1181) );
  INVX1 U779 ( .A(n1181), .Y(n1182) );
  AND2X2 U780 ( .A(\mem<10><15> ), .B(n179), .Y(n1183) );
  INVX1 U781 ( .A(n1183), .Y(n1184) );
  AND2X2 U782 ( .A(\mem<9><0> ), .B(n181), .Y(n1185) );
  INVX1 U783 ( .A(n1185), .Y(n1186) );
  AND2X2 U784 ( .A(\mem<9><8> ), .B(n181), .Y(n1187) );
  INVX1 U785 ( .A(n1187), .Y(n1188) );
  AND2X2 U786 ( .A(\mem<9><9> ), .B(n181), .Y(n1189) );
  INVX1 U787 ( .A(n1189), .Y(n1190) );
  AND2X2 U788 ( .A(\mem<9><10> ), .B(n181), .Y(n1191) );
  INVX1 U789 ( .A(n1191), .Y(n1192) );
  AND2X2 U790 ( .A(\mem<9><11> ), .B(n181), .Y(n1193) );
  INVX1 U791 ( .A(n1193), .Y(n1194) );
  AND2X2 U792 ( .A(\mem<9><12> ), .B(n181), .Y(n1195) );
  INVX1 U793 ( .A(n1195), .Y(n1196) );
  AND2X2 U794 ( .A(\mem<9><13> ), .B(n181), .Y(n1197) );
  INVX1 U795 ( .A(n1197), .Y(n1198) );
  AND2X2 U796 ( .A(\mem<9><14> ), .B(n181), .Y(n1199) );
  INVX1 U797 ( .A(n1199), .Y(n1200) );
  AND2X2 U798 ( .A(\mem<9><15> ), .B(n181), .Y(n1201) );
  INVX1 U799 ( .A(n1201), .Y(n1202) );
  AND2X1 U800 ( .A(N32), .B(n1953), .Y(n1203) );
  INVX1 U801 ( .A(n1203), .Y(n1204) );
  AND2X1 U802 ( .A(N31), .B(n1953), .Y(n1205) );
  INVX1 U803 ( .A(n1205), .Y(n1206) );
  AND2X1 U804 ( .A(N30), .B(n1953), .Y(n1207) );
  INVX1 U805 ( .A(n1207), .Y(n1208) );
  AND2X1 U806 ( .A(N29), .B(n1953), .Y(n1209) );
  INVX1 U807 ( .A(n1209), .Y(n1210) );
  AND2X1 U808 ( .A(N28), .B(n1953), .Y(n1211) );
  INVX1 U809 ( .A(n1211), .Y(n1212) );
  AND2X1 U810 ( .A(N27), .B(n1953), .Y(n1213) );
  INVX1 U811 ( .A(n1213), .Y(n1214) );
  AND2X1 U812 ( .A(N26), .B(n1953), .Y(n1215) );
  AND2X1 U813 ( .A(N24), .B(n1953), .Y(n1217) );
  INVX1 U814 ( .A(n1217), .Y(n1218) );
  AND2X1 U815 ( .A(N23), .B(n1953), .Y(n1219) );
  AND2X1 U816 ( .A(N22), .B(n1953), .Y(n1220) );
  INVX1 U817 ( .A(n1220), .Y(n1221) );
  AND2X1 U818 ( .A(N21), .B(n1953), .Y(n1222) );
  INVX1 U819 ( .A(n1222), .Y(n1223) );
  AND2X1 U820 ( .A(N20), .B(n1953), .Y(n1224) );
  AND2X1 U821 ( .A(N19), .B(n1953), .Y(n1225) );
  INVX1 U822 ( .A(n1225), .Y(n1226) );
  AND2X1 U823 ( .A(N18), .B(n1953), .Y(n1227) );
  AND2X1 U824 ( .A(N17), .B(n1953), .Y(n1228) );
  INVX1 U825 ( .A(n1228), .Y(n1229) );
  BUFX2 U826 ( .A(n1989), .Y(n1230) );
  INVX1 U827 ( .A(n1230), .Y(n2160) );
  BUFX2 U828 ( .A(n2006), .Y(n1231) );
  INVX1 U829 ( .A(n1231), .Y(n2169) );
  BUFX2 U830 ( .A(n2023), .Y(n1232) );
  INVX1 U831 ( .A(n1232), .Y(n2178) );
  BUFX2 U832 ( .A(n2040), .Y(n1233) );
  INVX1 U833 ( .A(n1233), .Y(n2187) );
  BUFX2 U834 ( .A(n2057), .Y(n1234) );
  INVX1 U835 ( .A(n1234), .Y(n2196) );
  BUFX2 U836 ( .A(n2133), .Y(n1235) );
  INVX1 U837 ( .A(n1235), .Y(n2134) );
  BUFX2 U838 ( .A(n2143), .Y(n1236) );
  INVX1 U839 ( .A(n1236), .Y(n2205) );
  AND2X1 U840 ( .A(n1954), .B(n491), .Y(n1237) );
  AND2X1 U841 ( .A(n1960), .B(n492), .Y(n1238) );
  AND2X1 U842 ( .A(n1955), .B(n491), .Y(n1239) );
  AND2X1 U843 ( .A(n1961), .B(n492), .Y(n1240) );
  INVX1 U844 ( .A(n206), .Y(\data_out<4> ) );
  AND2X1 U845 ( .A(n1238), .B(n2206), .Y(n1242) );
  AND2X1 U846 ( .A(n2206), .B(n1240), .Y(n1243) );
  AND2X1 U847 ( .A(n2206), .B(n2134), .Y(n1244) );
  AND2X1 U848 ( .A(n2206), .B(n2205), .Y(n1245) );
  AND2X1 U849 ( .A(n1237), .B(n1238), .Y(n1246) );
  INVX1 U850 ( .A(n1246), .Y(n1247) );
  AND2X1 U851 ( .A(n1238), .B(n1239), .Y(n1248) );
  INVX1 U852 ( .A(n1248), .Y(n1249) );
  BUFX2 U853 ( .A(n184), .Y(n1855) );
  AND2X1 U854 ( .A(n1238), .B(n2160), .Y(n1250) );
  INVX1 U855 ( .A(n1250), .Y(n1251) );
  AND2X1 U856 ( .A(n1238), .B(n2169), .Y(n1252) );
  INVX1 U857 ( .A(n1252), .Y(n1253) );
  AND2X1 U858 ( .A(n1238), .B(n2178), .Y(n1254) );
  INVX1 U859 ( .A(n1254), .Y(n1255) );
  AND2X1 U860 ( .A(n1238), .B(n2187), .Y(n1256) );
  INVX1 U861 ( .A(n1256), .Y(n1257) );
  AND2X1 U862 ( .A(n1238), .B(n2196), .Y(n1258) );
  INVX1 U863 ( .A(n1258), .Y(n1259) );
  AND2X1 U864 ( .A(n1237), .B(n1240), .Y(n1260) );
  INVX1 U865 ( .A(n1260), .Y(n1261) );
  AND2X1 U866 ( .A(n1239), .B(n1240), .Y(n1262) );
  INVX1 U867 ( .A(n1262), .Y(n1263) );
  AND2X1 U868 ( .A(n2160), .B(n1240), .Y(n1264) );
  INVX1 U869 ( .A(n1264), .Y(n1265) );
  AND2X1 U870 ( .A(n2169), .B(n1240), .Y(n1266) );
  INVX1 U871 ( .A(n1266), .Y(n1267) );
  AND2X1 U872 ( .A(n2178), .B(n1240), .Y(n1268) );
  INVX1 U873 ( .A(n1268), .Y(n1269) );
  AND2X1 U874 ( .A(n2187), .B(n1240), .Y(n1270) );
  INVX1 U875 ( .A(n1270), .Y(n1271) );
  AND2X1 U876 ( .A(n2196), .B(n1240), .Y(n1272) );
  INVX1 U877 ( .A(n1272), .Y(n1273) );
  AND2X1 U878 ( .A(n1237), .B(n2134), .Y(n1274) );
  INVX1 U879 ( .A(n1274), .Y(n1275) );
  AND2X1 U880 ( .A(n1239), .B(n2134), .Y(n1276) );
  INVX1 U881 ( .A(n1276), .Y(n1277) );
  AND2X1 U882 ( .A(n2160), .B(n2134), .Y(n1278) );
  INVX1 U883 ( .A(n1278), .Y(n1279) );
  AND2X1 U884 ( .A(n2169), .B(n2134), .Y(n1280) );
  INVX1 U885 ( .A(n1280), .Y(n1281) );
  AND2X1 U886 ( .A(n2178), .B(n2134), .Y(n1282) );
  INVX1 U887 ( .A(n1282), .Y(n1283) );
  AND2X1 U888 ( .A(n2187), .B(n2134), .Y(n1284) );
  INVX1 U889 ( .A(n1284), .Y(n1285) );
  AND2X1 U890 ( .A(n2196), .B(n2134), .Y(n1286) );
  INVX1 U891 ( .A(n1286), .Y(n1287) );
  AND2X1 U892 ( .A(n1237), .B(n2205), .Y(n1288) );
  INVX1 U893 ( .A(n1288), .Y(n1289) );
  AND2X1 U894 ( .A(n1239), .B(n2205), .Y(n1290) );
  INVX1 U895 ( .A(n1290), .Y(n1291) );
  AND2X1 U896 ( .A(n2160), .B(n2205), .Y(n1292) );
  INVX1 U897 ( .A(n1292), .Y(n1293) );
  AND2X1 U898 ( .A(n2169), .B(n2205), .Y(n1294) );
  INVX1 U899 ( .A(n1294), .Y(n1295) );
  AND2X1 U900 ( .A(n2178), .B(n2205), .Y(n1296) );
  INVX1 U901 ( .A(n1296), .Y(n1297) );
  AND2X1 U902 ( .A(n2187), .B(n2205), .Y(n1298) );
  INVX1 U903 ( .A(n1298), .Y(n1299) );
  AND2X1 U904 ( .A(n2196), .B(n2205), .Y(n1300) );
  INVX1 U905 ( .A(n1300), .Y(n1301) );
  INVX8 U906 ( .A(n1915), .Y(n1912) );
  INVX1 U907 ( .A(N11), .Y(n1957) );
  MUX2X1 U908 ( .B(n1303), .A(n1304), .S(n1809), .Y(n1302) );
  MUX2X1 U909 ( .B(n1306), .A(n1307), .S(n1809), .Y(n1305) );
  MUX2X1 U910 ( .B(n1309), .A(n1310), .S(n1809), .Y(n1308) );
  MUX2X1 U911 ( .B(n1312), .A(n1313), .S(n1809), .Y(n1311) );
  MUX2X1 U912 ( .B(n1315), .A(n1316), .S(n1801), .Y(n1314) );
  MUX2X1 U913 ( .B(n1318), .A(n1319), .S(n1809), .Y(n1317) );
  MUX2X1 U914 ( .B(n1321), .A(n1322), .S(n1809), .Y(n1320) );
  MUX2X1 U915 ( .B(n1324), .A(n1325), .S(n1809), .Y(n1323) );
  MUX2X1 U916 ( .B(n1327), .A(n1328), .S(n1809), .Y(n1326) );
  MUX2X1 U917 ( .B(n1330), .A(n1331), .S(n1801), .Y(n1329) );
  MUX2X1 U918 ( .B(n1333), .A(n1334), .S(n1810), .Y(n1332) );
  MUX2X1 U919 ( .B(n1336), .A(n1337), .S(n1810), .Y(n1335) );
  MUX2X1 U920 ( .B(n1339), .A(n1340), .S(n1810), .Y(n1338) );
  MUX2X1 U921 ( .B(n1342), .A(n1343), .S(n1810), .Y(n1341) );
  MUX2X1 U922 ( .B(n1345), .A(n1346), .S(n1801), .Y(n1344) );
  MUX2X1 U923 ( .B(n1348), .A(n1349), .S(n1810), .Y(n1347) );
  MUX2X1 U924 ( .B(n1351), .A(n1352), .S(n1810), .Y(n1350) );
  MUX2X1 U925 ( .B(n1354), .A(n1355), .S(n1810), .Y(n1353) );
  MUX2X1 U926 ( .B(n1357), .A(n1358), .S(n1810), .Y(n1356) );
  MUX2X1 U927 ( .B(n1360), .A(n1361), .S(n1801), .Y(n1359) );
  MUX2X1 U928 ( .B(n1363), .A(n1364), .S(n1810), .Y(n1362) );
  MUX2X1 U929 ( .B(n1366), .A(n1367), .S(n1810), .Y(n1365) );
  MUX2X1 U930 ( .B(n1369), .A(n1370), .S(n1810), .Y(n1368) );
  MUX2X1 U931 ( .B(n1372), .A(n1373), .S(n1810), .Y(n1371) );
  MUX2X1 U932 ( .B(n1375), .A(n1376), .S(n1801), .Y(n1374) );
  MUX2X1 U933 ( .B(n1378), .A(n1379), .S(n1811), .Y(n1377) );
  MUX2X1 U934 ( .B(n1381), .A(n1382), .S(n1811), .Y(n1380) );
  MUX2X1 U935 ( .B(n1384), .A(n1385), .S(n1811), .Y(n1383) );
  MUX2X1 U936 ( .B(n1387), .A(n1388), .S(n1811), .Y(n1386) );
  MUX2X1 U937 ( .B(n1390), .A(n1391), .S(n1801), .Y(n1389) );
  MUX2X1 U938 ( .B(n1393), .A(n1394), .S(n1811), .Y(n1392) );
  MUX2X1 U939 ( .B(n1396), .A(n1397), .S(n1811), .Y(n1395) );
  MUX2X1 U940 ( .B(n1399), .A(n1400), .S(n1811), .Y(n1398) );
  MUX2X1 U941 ( .B(n1402), .A(n1403), .S(n1811), .Y(n1401) );
  MUX2X1 U942 ( .B(n1405), .A(n1406), .S(n1801), .Y(n1404) );
  MUX2X1 U943 ( .B(n1408), .A(n1409), .S(n1811), .Y(n1407) );
  MUX2X1 U944 ( .B(n1411), .A(n1412), .S(n1811), .Y(n1410) );
  MUX2X1 U945 ( .B(n1414), .A(n1415), .S(n1811), .Y(n1413) );
  MUX2X1 U946 ( .B(n1417), .A(n1418), .S(n1811), .Y(n1416) );
  MUX2X1 U947 ( .B(n1420), .A(n1421), .S(n1801), .Y(n1419) );
  MUX2X1 U948 ( .B(n1423), .A(n1424), .S(n1812), .Y(n1422) );
  MUX2X1 U949 ( .B(n1426), .A(n1427), .S(n1812), .Y(n1425) );
  MUX2X1 U950 ( .B(n1429), .A(n1430), .S(n1812), .Y(n1428) );
  MUX2X1 U951 ( .B(n1432), .A(n1433), .S(n1812), .Y(n1431) );
  MUX2X1 U952 ( .B(n1435), .A(n1436), .S(n1801), .Y(n1434) );
  MUX2X1 U953 ( .B(n1438), .A(n1439), .S(n1812), .Y(n1437) );
  MUX2X1 U954 ( .B(n1441), .A(n1442), .S(n1812), .Y(n1440) );
  MUX2X1 U955 ( .B(n1444), .A(n1445), .S(n1812), .Y(n1443) );
  MUX2X1 U956 ( .B(n1447), .A(n1448), .S(n1812), .Y(n1446) );
  MUX2X1 U957 ( .B(n1450), .A(n1451), .S(n1801), .Y(n1449) );
  MUX2X1 U958 ( .B(n1453), .A(n1454), .S(n1812), .Y(n1452) );
  MUX2X1 U959 ( .B(n1456), .A(n1457), .S(n1812), .Y(n1455) );
  MUX2X1 U960 ( .B(n1459), .A(n1460), .S(n1812), .Y(n1458) );
  MUX2X1 U961 ( .B(n1462), .A(n1463), .S(n1812), .Y(n1461) );
  MUX2X1 U962 ( .B(n1465), .A(n1466), .S(n1801), .Y(n1464) );
  MUX2X1 U963 ( .B(n1468), .A(n1469), .S(n1813), .Y(n1467) );
  MUX2X1 U964 ( .B(n1471), .A(n1472), .S(n1813), .Y(n1470) );
  MUX2X1 U965 ( .B(n1474), .A(n1475), .S(n1813), .Y(n1473) );
  MUX2X1 U966 ( .B(n1477), .A(n1478), .S(n1813), .Y(n1476) );
  MUX2X1 U967 ( .B(n1480), .A(n1481), .S(n1801), .Y(n1479) );
  MUX2X1 U968 ( .B(n1483), .A(n1484), .S(n1813), .Y(n1482) );
  MUX2X1 U969 ( .B(n1486), .A(n1487), .S(n1813), .Y(n1485) );
  MUX2X1 U970 ( .B(n1489), .A(n1490), .S(n1813), .Y(n1488) );
  MUX2X1 U971 ( .B(n1492), .A(n1493), .S(n1813), .Y(n1491) );
  MUX2X1 U972 ( .B(n1495), .A(n1496), .S(n1800), .Y(n1494) );
  MUX2X1 U973 ( .B(n1498), .A(n1499), .S(n1813), .Y(n1497) );
  MUX2X1 U974 ( .B(n1501), .A(n1502), .S(n1813), .Y(n1500) );
  MUX2X1 U975 ( .B(n1504), .A(n1505), .S(n1813), .Y(n1503) );
  MUX2X1 U976 ( .B(n1507), .A(n1508), .S(n1813), .Y(n1506) );
  MUX2X1 U977 ( .B(n1510), .A(n1511), .S(n1800), .Y(n1509) );
  MUX2X1 U978 ( .B(n1513), .A(n1514), .S(n1814), .Y(n1512) );
  MUX2X1 U979 ( .B(n1516), .A(n1517), .S(n1814), .Y(n1515) );
  MUX2X1 U980 ( .B(n1519), .A(n1520), .S(n1814), .Y(n1518) );
  MUX2X1 U981 ( .B(n1522), .A(n1523), .S(n1814), .Y(n1521) );
  MUX2X1 U982 ( .B(n1525), .A(n1526), .S(n1800), .Y(n1524) );
  MUX2X1 U983 ( .B(n1528), .A(n1529), .S(n1814), .Y(n1527) );
  MUX2X1 U984 ( .B(n1531), .A(n1532), .S(n1814), .Y(n1530) );
  MUX2X1 U985 ( .B(n1534), .A(n1535), .S(n1814), .Y(n1533) );
  MUX2X1 U986 ( .B(n1537), .A(n1538), .S(n1814), .Y(n1536) );
  MUX2X1 U987 ( .B(n1540), .A(n1541), .S(n1800), .Y(n1539) );
  MUX2X1 U988 ( .B(n1543), .A(n1544), .S(n1814), .Y(n1542) );
  MUX2X1 U989 ( .B(n1546), .A(n1547), .S(n1814), .Y(n1545) );
  MUX2X1 U990 ( .B(n1549), .A(n1550), .S(n1814), .Y(n1548) );
  MUX2X1 U991 ( .B(n1552), .A(n1553), .S(n1814), .Y(n1551) );
  MUX2X1 U992 ( .B(n1555), .A(n1556), .S(n1800), .Y(n1554) );
  MUX2X1 U993 ( .B(n1558), .A(n1559), .S(n1815), .Y(n1557) );
  MUX2X1 U994 ( .B(n1561), .A(n1562), .S(n1815), .Y(n1560) );
  MUX2X1 U995 ( .B(n1564), .A(n1565), .S(n1815), .Y(n1563) );
  MUX2X1 U996 ( .B(n1567), .A(n1568), .S(n1815), .Y(n1566) );
  MUX2X1 U997 ( .B(n1570), .A(n1571), .S(n1800), .Y(n1569) );
  MUX2X1 U998 ( .B(n1573), .A(n1574), .S(n1815), .Y(n1572) );
  MUX2X1 U999 ( .B(n1576), .A(n1577), .S(n1815), .Y(n1575) );
  MUX2X1 U1000 ( .B(n1579), .A(n1580), .S(n1815), .Y(n1578) );
  MUX2X1 U1001 ( .B(n1582), .A(n1583), .S(n1815), .Y(n1581) );
  MUX2X1 U1002 ( .B(n1585), .A(n1586), .S(n1800), .Y(n1584) );
  MUX2X1 U1003 ( .B(n1588), .A(n1589), .S(n1815), .Y(n1587) );
  MUX2X1 U1004 ( .B(n1591), .A(n1592), .S(n1815), .Y(n1590) );
  MUX2X1 U1005 ( .B(n1594), .A(n1595), .S(n1815), .Y(n1593) );
  MUX2X1 U1006 ( .B(n1597), .A(n1598), .S(n1815), .Y(n1596) );
  MUX2X1 U1007 ( .B(n1600), .A(n1601), .S(n1800), .Y(n1599) );
  MUX2X1 U1008 ( .B(n1603), .A(n1604), .S(n1816), .Y(n1602) );
  MUX2X1 U1009 ( .B(n1606), .A(n1607), .S(n1816), .Y(n1605) );
  MUX2X1 U1010 ( .B(n1609), .A(n1610), .S(n1816), .Y(n1608) );
  MUX2X1 U1011 ( .B(n1612), .A(n1613), .S(n1816), .Y(n1611) );
  MUX2X1 U1012 ( .B(n1615), .A(n1616), .S(n1800), .Y(n1614) );
  MUX2X1 U1013 ( .B(n1618), .A(n1619), .S(n1816), .Y(n1617) );
  MUX2X1 U1014 ( .B(n1621), .A(n1622), .S(n1816), .Y(n1620) );
  MUX2X1 U1015 ( .B(n1624), .A(n1625), .S(n1816), .Y(n1623) );
  MUX2X1 U1016 ( .B(n1627), .A(n1628), .S(n1816), .Y(n1626) );
  MUX2X1 U1017 ( .B(n1630), .A(n1631), .S(n1800), .Y(n1629) );
  MUX2X1 U1018 ( .B(n1633), .A(n1634), .S(n1816), .Y(n1632) );
  MUX2X1 U1019 ( .B(n1636), .A(n1637), .S(n1816), .Y(n1635) );
  MUX2X1 U1020 ( .B(n1639), .A(n1640), .S(n1816), .Y(n1638) );
  MUX2X1 U1021 ( .B(n1642), .A(n1643), .S(n1816), .Y(n1641) );
  MUX2X1 U1022 ( .B(n1645), .A(n1646), .S(n1800), .Y(n1644) );
  MUX2X1 U1023 ( .B(n1648), .A(n1649), .S(n1817), .Y(n1647) );
  MUX2X1 U1024 ( .B(n1651), .A(n1652), .S(n1817), .Y(n1650) );
  MUX2X1 U1025 ( .B(n1654), .A(n1655), .S(n1817), .Y(n1653) );
  MUX2X1 U1026 ( .B(n1657), .A(n1658), .S(n1817), .Y(n1656) );
  MUX2X1 U1027 ( .B(n1660), .A(n1661), .S(n1800), .Y(n1659) );
  MUX2X1 U1028 ( .B(n1663), .A(n1664), .S(n1817), .Y(n1662) );
  MUX2X1 U1029 ( .B(n1666), .A(n1667), .S(n1817), .Y(n1665) );
  MUX2X1 U1030 ( .B(n1669), .A(n1670), .S(n1817), .Y(n1668) );
  MUX2X1 U1031 ( .B(n1672), .A(n1673), .S(n1817), .Y(n1671) );
  MUX2X1 U1032 ( .B(n1675), .A(n1676), .S(n1960), .Y(n1674) );
  MUX2X1 U1033 ( .B(n1678), .A(n1679), .S(n1817), .Y(n1677) );
  MUX2X1 U1034 ( .B(n1681), .A(n1682), .S(n1817), .Y(n1680) );
  MUX2X1 U1035 ( .B(n1684), .A(n1685), .S(n1817), .Y(n1683) );
  MUX2X1 U1036 ( .B(n1687), .A(n1688), .S(n1817), .Y(n1686) );
  MUX2X1 U1037 ( .B(n1690), .A(n1691), .S(n1801), .Y(n1689) );
  MUX2X1 U1038 ( .B(n1693), .A(n1694), .S(n1818), .Y(n1692) );
  MUX2X1 U1039 ( .B(n1696), .A(n1697), .S(n1818), .Y(n1695) );
  MUX2X1 U1040 ( .B(n1699), .A(n1700), .S(n1818), .Y(n1698) );
  MUX2X1 U1041 ( .B(n1702), .A(n1703), .S(n1818), .Y(n1701) );
  MUX2X1 U1042 ( .B(n1705), .A(n1706), .S(n1801), .Y(n1704) );
  MUX2X1 U1043 ( .B(n1708), .A(n1709), .S(n1818), .Y(n1707) );
  MUX2X1 U1044 ( .B(n1711), .A(n1712), .S(n1818), .Y(n1710) );
  MUX2X1 U1045 ( .B(n1714), .A(n1715), .S(n1818), .Y(n1713) );
  MUX2X1 U1046 ( .B(n1717), .A(n1718), .S(n1818), .Y(n1716) );
  MUX2X1 U1047 ( .B(n1720), .A(n1721), .S(n1960), .Y(n1719) );
  MUX2X1 U1048 ( .B(n1723), .A(n1724), .S(n1818), .Y(n1722) );
  MUX2X1 U1049 ( .B(n1726), .A(n1727), .S(n1818), .Y(n1725) );
  MUX2X1 U1050 ( .B(n1729), .A(n1730), .S(n1818), .Y(n1728) );
  MUX2X1 U1051 ( .B(n1732), .A(n1733), .S(n1818), .Y(n1731) );
  MUX2X1 U1052 ( .B(n1735), .A(n1736), .S(n1801), .Y(n1734) );
  MUX2X1 U1053 ( .B(n1738), .A(n1739), .S(n1819), .Y(n1737) );
  MUX2X1 U1054 ( .B(n1741), .A(n1742), .S(n1819), .Y(n1740) );
  MUX2X1 U1055 ( .B(n1744), .A(n1745), .S(n1819), .Y(n1743) );
  MUX2X1 U1056 ( .B(n1747), .A(n1748), .S(n1819), .Y(n1746) );
  MUX2X1 U1057 ( .B(n1750), .A(n1751), .S(n1801), .Y(n1749) );
  MUX2X1 U1058 ( .B(n1753), .A(n1754), .S(n1819), .Y(n1752) );
  MUX2X1 U1059 ( .B(n1756), .A(n1757), .S(n1819), .Y(n1755) );
  MUX2X1 U1060 ( .B(n1759), .A(n1760), .S(n1819), .Y(n1758) );
  MUX2X1 U1061 ( .B(n1762), .A(n1763), .S(n1819), .Y(n1761) );
  MUX2X1 U1062 ( .B(n1765), .A(n1766), .S(n1801), .Y(n1764) );
  MUX2X1 U1063 ( .B(n1768), .A(n1769), .S(n1819), .Y(n1767) );
  MUX2X1 U1064 ( .B(n1771), .A(n1772), .S(n1819), .Y(n1770) );
  MUX2X1 U1065 ( .B(n1774), .A(n1775), .S(n1819), .Y(n1773) );
  MUX2X1 U1066 ( .B(n1777), .A(n1778), .S(n1819), .Y(n1776) );
  MUX2X1 U1067 ( .B(n1780), .A(n1781), .S(n1801), .Y(n1779) );
  MUX2X1 U1068 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1829), .Y(n1304) );
  MUX2X1 U1069 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1829), .Y(n1303) );
  MUX2X1 U1070 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1829), .Y(n1307) );
  MUX2X1 U1071 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1829), .Y(n1306) );
  MUX2X1 U1072 ( .B(n1305), .A(n1302), .S(n1806), .Y(n1316) );
  MUX2X1 U1073 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1840), .Y(n1310) );
  MUX2X1 U1074 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1844), .Y(n1309) );
  MUX2X1 U1075 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1844), .Y(n1313) );
  MUX2X1 U1076 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1836), .Y(n1312) );
  MUX2X1 U1077 ( .B(n1311), .A(n1308), .S(n1806), .Y(n1315) );
  MUX2X1 U1078 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1832), .Y(n1319) );
  MUX2X1 U1079 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1832), .Y(n1318) );
  MUX2X1 U1080 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1829), .Y(n1322) );
  MUX2X1 U1081 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1829), .Y(n1321) );
  MUX2X1 U1082 ( .B(n1320), .A(n1317), .S(n1806), .Y(n1331) );
  MUX2X1 U1083 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1847), .Y(n1325) );
  MUX2X1 U1084 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1837), .Y(n1324) );
  MUX2X1 U1085 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1829), .Y(n1328) );
  MUX2X1 U1086 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1829), .Y(n1327) );
  MUX2X1 U1087 ( .B(n1326), .A(n1323), .S(n1806), .Y(n1330) );
  MUX2X1 U1088 ( .B(n1329), .A(n1314), .S(n1799), .Y(n1782) );
  MUX2X1 U1089 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1830), .Y(n1334) );
  MUX2X1 U1090 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1830), .Y(n1333) );
  MUX2X1 U1091 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1830), .Y(n1337) );
  MUX2X1 U1092 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1830), .Y(n1336) );
  MUX2X1 U1093 ( .B(n1335), .A(n1332), .S(n1806), .Y(n1346) );
  MUX2X1 U1094 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1830), .Y(n1340) );
  MUX2X1 U1095 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1830), .Y(n1339) );
  MUX2X1 U1096 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1830), .Y(n1343) );
  MUX2X1 U1097 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1830), .Y(n1342) );
  MUX2X1 U1098 ( .B(n1341), .A(n1338), .S(n1806), .Y(n1345) );
  MUX2X1 U1099 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1830), .Y(n1349) );
  MUX2X1 U1100 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1830), .Y(n1348) );
  MUX2X1 U1101 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1830), .Y(n1352) );
  MUX2X1 U1102 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1830), .Y(n1351) );
  MUX2X1 U1103 ( .B(n1350), .A(n1347), .S(n1806), .Y(n1361) );
  MUX2X1 U1104 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1831), .Y(n1355) );
  MUX2X1 U1105 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1831), .Y(n1354) );
  MUX2X1 U1106 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1831), .Y(n1358) );
  MUX2X1 U1107 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1831), .Y(n1357) );
  MUX2X1 U1108 ( .B(n1356), .A(n1353), .S(n1806), .Y(n1360) );
  MUX2X1 U1109 ( .B(n1359), .A(n1344), .S(n1799), .Y(n1783) );
  MUX2X1 U1110 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1831), .Y(n1364) );
  MUX2X1 U1111 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1831), .Y(n1363) );
  MUX2X1 U1112 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1831), .Y(n1367) );
  MUX2X1 U1113 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1831), .Y(n1366) );
  MUX2X1 U1114 ( .B(n1365), .A(n1362), .S(n1806), .Y(n1376) );
  MUX2X1 U1115 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1831), .Y(n1370) );
  MUX2X1 U1116 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1831), .Y(n1369) );
  MUX2X1 U1117 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1831), .Y(n1373) );
  MUX2X1 U1118 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1831), .Y(n1372) );
  MUX2X1 U1119 ( .B(n1371), .A(n1368), .S(n1806), .Y(n1375) );
  MUX2X1 U1120 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1832), .Y(n1379) );
  MUX2X1 U1121 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1832), .Y(n1378) );
  MUX2X1 U1122 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1832), .Y(n1382) );
  MUX2X1 U1123 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1832), .Y(n1381) );
  MUX2X1 U1124 ( .B(n1380), .A(n1377), .S(n1806), .Y(n1391) );
  MUX2X1 U1125 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1832), .Y(n1385) );
  MUX2X1 U1126 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1832), .Y(n1384) );
  MUX2X1 U1127 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1832), .Y(n1388) );
  MUX2X1 U1128 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1832), .Y(n1387) );
  MUX2X1 U1129 ( .B(n1386), .A(n1383), .S(n1806), .Y(n1390) );
  MUX2X1 U1130 ( .B(n1389), .A(n1374), .S(n1799), .Y(n1784) );
  MUX2X1 U1131 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1832), .Y(n1394) );
  MUX2X1 U1132 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1832), .Y(n1393) );
  MUX2X1 U1133 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1832), .Y(n1397) );
  MUX2X1 U1134 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1832), .Y(n1396) );
  MUX2X1 U1135 ( .B(n1395), .A(n1392), .S(n1805), .Y(n1406) );
  MUX2X1 U1136 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1833), .Y(n1400) );
  MUX2X1 U1137 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1833), .Y(n1399) );
  MUX2X1 U1138 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1833), .Y(n1403) );
  MUX2X1 U1139 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1833), .Y(n1402) );
  MUX2X1 U1140 ( .B(n1401), .A(n1398), .S(n1805), .Y(n1405) );
  MUX2X1 U1141 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1833), .Y(n1409) );
  MUX2X1 U1142 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1833), .Y(n1408) );
  MUX2X1 U1143 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1833), .Y(n1412) );
  MUX2X1 U1144 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1833), .Y(n1411) );
  MUX2X1 U1145 ( .B(n1410), .A(n1407), .S(n1805), .Y(n1421) );
  MUX2X1 U1146 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1833), .Y(n1415) );
  MUX2X1 U1147 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1833), .Y(n1414) );
  MUX2X1 U1148 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1833), .Y(n1418) );
  MUX2X1 U1149 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1833), .Y(n1417) );
  MUX2X1 U1150 ( .B(n1416), .A(n1413), .S(n1805), .Y(n1420) );
  MUX2X1 U1151 ( .B(n1419), .A(n1404), .S(n1799), .Y(n1785) );
  MUX2X1 U1152 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1834), .Y(n1424) );
  MUX2X1 U1153 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1834), .Y(n1423) );
  MUX2X1 U1154 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1834), .Y(n1427) );
  MUX2X1 U1155 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1834), .Y(n1426) );
  MUX2X1 U1156 ( .B(n1425), .A(n1422), .S(n1805), .Y(n1436) );
  MUX2X1 U1157 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1834), .Y(n1430) );
  MUX2X1 U1158 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1834), .Y(n1429) );
  MUX2X1 U1159 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1834), .Y(n1433) );
  MUX2X1 U1160 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1834), .Y(n1432) );
  MUX2X1 U1161 ( .B(n1431), .A(n1428), .S(n1805), .Y(n1435) );
  MUX2X1 U1162 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1834), .Y(n1439) );
  MUX2X1 U1163 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1834), .Y(n1438) );
  MUX2X1 U1164 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1834), .Y(n1442) );
  MUX2X1 U1165 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1834), .Y(n1441) );
  MUX2X1 U1166 ( .B(n1440), .A(n1437), .S(n1805), .Y(n1451) );
  MUX2X1 U1167 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1836), .Y(n1445) );
  MUX2X1 U1168 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1844), .Y(n1444) );
  MUX2X1 U1169 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1829), .Y(n1448) );
  MUX2X1 U1170 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1829), .Y(n1447) );
  MUX2X1 U1171 ( .B(n1446), .A(n1443), .S(n1805), .Y(n1450) );
  MUX2X1 U1172 ( .B(n1449), .A(n1434), .S(n1799), .Y(n1786) );
  MUX2X1 U1173 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1844), .Y(n1454) );
  MUX2X1 U1174 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1836), .Y(n1453) );
  MUX2X1 U1175 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1840), .Y(n1457) );
  MUX2X1 U1177 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1840), .Y(n1456) );
  MUX2X1 U1178 ( .B(n1455), .A(n1452), .S(n1805), .Y(n1466) );
  MUX2X1 U1179 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1840), .Y(n1460) );
  MUX2X1 U1180 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1837), .Y(n1459) );
  MUX2X1 U1181 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1844), .Y(n1463) );
  MUX2X1 U1182 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1837), .Y(n1462) );
  MUX2X1 U1183 ( .B(n1461), .A(n1458), .S(n1805), .Y(n1465) );
  MUX2X1 U1184 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1835), .Y(n1469) );
  MUX2X1 U1185 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1835), .Y(n1468) );
  MUX2X1 U1186 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1835), .Y(n1472) );
  MUX2X1 U1187 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1835), .Y(n1471) );
  MUX2X1 U1188 ( .B(n1470), .A(n1467), .S(n1805), .Y(n1481) );
  MUX2X1 U1189 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1835), .Y(n1475) );
  MUX2X1 U1190 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1835), .Y(n1474) );
  MUX2X1 U1191 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1835), .Y(n1478) );
  MUX2X1 U1192 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1835), .Y(n1477) );
  MUX2X1 U1193 ( .B(n1476), .A(n1473), .S(n1805), .Y(n1480) );
  MUX2X1 U1194 ( .B(n1479), .A(n1464), .S(n1799), .Y(n1787) );
  MUX2X1 U1195 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1835), .Y(n1484) );
  MUX2X1 U1196 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1835), .Y(n1483) );
  MUX2X1 U1197 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1835), .Y(n1487) );
  MUX2X1 U1198 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1835), .Y(n1486) );
  MUX2X1 U1199 ( .B(n1485), .A(n1482), .S(n1805), .Y(n1496) );
  MUX2X1 U1200 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1836), .Y(n1490) );
  MUX2X1 U1201 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1836), .Y(n1489) );
  MUX2X1 U1202 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1836), .Y(n1493) );
  MUX2X1 U1203 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1836), .Y(n1492) );
  MUX2X1 U1204 ( .B(n1491), .A(n1488), .S(n1806), .Y(n1495) );
  MUX2X1 U1205 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1836), .Y(n1499) );
  MUX2X1 U1206 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1836), .Y(n1498) );
  MUX2X1 U1207 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1836), .Y(n1502) );
  MUX2X1 U1208 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1836), .Y(n1501) );
  MUX2X1 U1209 ( .B(n1500), .A(n1497), .S(n1805), .Y(n1511) );
  MUX2X1 U1210 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1836), .Y(n1505) );
  MUX2X1 U1211 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1836), .Y(n1504) );
  MUX2X1 U1212 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1836), .Y(n1508) );
  MUX2X1 U1213 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1836), .Y(n1507) );
  MUX2X1 U1214 ( .B(n1506), .A(n1503), .S(n1806), .Y(n1510) );
  MUX2X1 U1215 ( .B(n1509), .A(n1494), .S(n1799), .Y(n1788) );
  MUX2X1 U1216 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1837), .Y(n1514) );
  MUX2X1 U1217 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1837), .Y(n1513) );
  MUX2X1 U1218 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1837), .Y(n1517) );
  MUX2X1 U1219 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1837), .Y(n1516) );
  MUX2X1 U1220 ( .B(n1515), .A(n1512), .S(n1805), .Y(n1526) );
  MUX2X1 U1221 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1837), .Y(n1520) );
  MUX2X1 U1222 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1837), .Y(n1519) );
  MUX2X1 U1223 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1837), .Y(n1523) );
  MUX2X1 U1224 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1837), .Y(n1522) );
  MUX2X1 U1225 ( .B(n1521), .A(n1518), .S(n1806), .Y(n1525) );
  MUX2X1 U1226 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1837), .Y(n1529) );
  MUX2X1 U1227 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1837), .Y(n1528) );
  MUX2X1 U1228 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1837), .Y(n1532) );
  MUX2X1 U1229 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1837), .Y(n1531) );
  MUX2X1 U1230 ( .B(n1530), .A(n1527), .S(n1805), .Y(n1541) );
  MUX2X1 U1231 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1838), .Y(n1535) );
  MUX2X1 U1232 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1838), .Y(n1534) );
  MUX2X1 U1233 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1838), .Y(n1538) );
  MUX2X1 U1234 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1838), .Y(n1537) );
  MUX2X1 U1235 ( .B(n1536), .A(n1533), .S(n1806), .Y(n1540) );
  MUX2X1 U1236 ( .B(n1539), .A(n1524), .S(n1799), .Y(n1789) );
  MUX2X1 U1237 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1838), .Y(n1544) );
  MUX2X1 U1238 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1838), .Y(n1543) );
  MUX2X1 U1239 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1838), .Y(n1547) );
  MUX2X1 U1240 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1838), .Y(n1546) );
  MUX2X1 U1241 ( .B(n1545), .A(n1542), .S(n1806), .Y(n1556) );
  MUX2X1 U1242 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1838), .Y(n1550) );
  MUX2X1 U1243 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1838), .Y(n1549) );
  MUX2X1 U1244 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1838), .Y(n1553) );
  MUX2X1 U1245 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1838), .Y(n1552) );
  MUX2X1 U1246 ( .B(n1551), .A(n1548), .S(n1806), .Y(n1555) );
  MUX2X1 U1247 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1839), .Y(n1559) );
  MUX2X1 U1248 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1839), .Y(n1558) );
  MUX2X1 U1249 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1839), .Y(n1562) );
  MUX2X1 U1250 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1839), .Y(n1561) );
  MUX2X1 U1251 ( .B(n1560), .A(n1557), .S(n1805), .Y(n1571) );
  MUX2X1 U1252 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1839), .Y(n1565) );
  MUX2X1 U1253 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1839), .Y(n1564) );
  MUX2X1 U1254 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1839), .Y(n1568) );
  MUX2X1 U1255 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1839), .Y(n1567) );
  MUX2X1 U1256 ( .B(n1566), .A(n1563), .S(n1806), .Y(n1570) );
  MUX2X1 U1257 ( .B(n1569), .A(n1554), .S(n1799), .Y(n1790) );
  MUX2X1 U1258 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1839), .Y(n1574) );
  MUX2X1 U1259 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1839), .Y(n1573) );
  MUX2X1 U1260 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1839), .Y(n1577) );
  MUX2X1 U1261 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1839), .Y(n1576) );
  MUX2X1 U1262 ( .B(n1575), .A(n1572), .S(n1804), .Y(n1586) );
  MUX2X1 U1263 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1840), .Y(n1580) );
  MUX2X1 U1264 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1840), .Y(n1579) );
  MUX2X1 U1265 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1840), .Y(n1583) );
  MUX2X1 U1266 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1840), .Y(n1582) );
  MUX2X1 U1267 ( .B(n1581), .A(n1578), .S(n1804), .Y(n1585) );
  MUX2X1 U1268 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1840), .Y(n1589) );
  MUX2X1 U1269 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1840), .Y(n1588) );
  MUX2X1 U1270 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1840), .Y(n1592) );
  MUX2X1 U1271 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1840), .Y(n1591) );
  MUX2X1 U1272 ( .B(n1590), .A(n1587), .S(n1804), .Y(n1601) );
  MUX2X1 U1273 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1840), .Y(n1595) );
  MUX2X1 U1274 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1840), .Y(n1594) );
  MUX2X1 U1275 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1840), .Y(n1598) );
  MUX2X1 U1276 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1840), .Y(n1597) );
  MUX2X1 U1277 ( .B(n1596), .A(n1593), .S(n1804), .Y(n1600) );
  MUX2X1 U1278 ( .B(n1599), .A(n1584), .S(n1799), .Y(n1791) );
  MUX2X1 U1279 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1841), .Y(n1604) );
  MUX2X1 U1280 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1841), .Y(n1603) );
  MUX2X1 U1281 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1841), .Y(n1607) );
  MUX2X1 U1282 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1841), .Y(n1606) );
  MUX2X1 U1283 ( .B(n1605), .A(n1602), .S(n1804), .Y(n1616) );
  MUX2X1 U1284 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1841), .Y(n1610) );
  MUX2X1 U1285 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1841), .Y(n1609) );
  MUX2X1 U1286 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1841), .Y(n1613) );
  MUX2X1 U1287 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1841), .Y(n1612) );
  MUX2X1 U1288 ( .B(n1611), .A(n1608), .S(n1804), .Y(n1615) );
  MUX2X1 U1289 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1841), .Y(n1619) );
  MUX2X1 U1290 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1841), .Y(n1618) );
  MUX2X1 U1291 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1841), .Y(n1622) );
  MUX2X1 U1292 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1841), .Y(n1621) );
  MUX2X1 U1293 ( .B(n1620), .A(n1617), .S(n1804), .Y(n1631) );
  MUX2X1 U1294 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1842), .Y(n1625) );
  MUX2X1 U1295 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1842), .Y(n1624) );
  MUX2X1 U1296 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1842), .Y(n1628) );
  MUX2X1 U1297 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1842), .Y(n1627) );
  MUX2X1 U1298 ( .B(n1626), .A(n1623), .S(n1804), .Y(n1630) );
  MUX2X1 U1299 ( .B(n1629), .A(n1614), .S(n1799), .Y(n1792) );
  MUX2X1 U1300 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1842), .Y(n1634) );
  MUX2X1 U1301 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1842), .Y(n1633) );
  MUX2X1 U1302 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1842), .Y(n1637) );
  MUX2X1 U1303 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1842), .Y(n1636) );
  MUX2X1 U1304 ( .B(n1635), .A(n1632), .S(n1804), .Y(n1646) );
  MUX2X1 U1305 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1842), .Y(n1640) );
  MUX2X1 U1306 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1842), .Y(n1639) );
  MUX2X1 U1307 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1842), .Y(n1643) );
  MUX2X1 U1308 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1842), .Y(n1642) );
  MUX2X1 U1309 ( .B(n1641), .A(n1638), .S(n1804), .Y(n1645) );
  MUX2X1 U1310 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1843), .Y(n1649) );
  MUX2X1 U1311 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1843), .Y(n1648) );
  MUX2X1 U1312 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1843), .Y(n1652) );
  MUX2X1 U1313 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1843), .Y(n1651) );
  MUX2X1 U1314 ( .B(n1650), .A(n1647), .S(n1804), .Y(n1661) );
  MUX2X1 U1315 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1843), .Y(n1655) );
  MUX2X1 U1316 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1843), .Y(n1654) );
  MUX2X1 U1317 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1843), .Y(n1658) );
  MUX2X1 U1318 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1843), .Y(n1657) );
  MUX2X1 U1319 ( .B(n1656), .A(n1653), .S(n1804), .Y(n1660) );
  MUX2X1 U1320 ( .B(n1659), .A(n1644), .S(n1799), .Y(n1793) );
  MUX2X1 U1321 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1843), .Y(n1664) );
  MUX2X1 U1322 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1843), .Y(n1663) );
  MUX2X1 U1323 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1843), .Y(n1667) );
  MUX2X1 U1324 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1843), .Y(n1666) );
  MUX2X1 U1325 ( .B(n1665), .A(n1662), .S(n1803), .Y(n1676) );
  MUX2X1 U1326 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1844), .Y(n1670) );
  MUX2X1 U1327 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1844), .Y(n1669) );
  MUX2X1 U1328 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1844), .Y(n1673) );
  MUX2X1 U1329 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1844), .Y(n1672) );
  MUX2X1 U1330 ( .B(n1671), .A(n1668), .S(n1803), .Y(n1675) );
  MUX2X1 U1331 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1844), .Y(n1679) );
  MUX2X1 U1332 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1844), .Y(n1678) );
  MUX2X1 U1333 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1844), .Y(n1682) );
  MUX2X1 U1334 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1844), .Y(n1681) );
  MUX2X1 U1335 ( .B(n1680), .A(n1677), .S(n1803), .Y(n1691) );
  MUX2X1 U1336 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1844), .Y(n1685) );
  MUX2X1 U1337 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1844), .Y(n1684) );
  MUX2X1 U1338 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1844), .Y(n1688) );
  MUX2X1 U1339 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1844), .Y(n1687) );
  MUX2X1 U1340 ( .B(n1686), .A(n1683), .S(n1803), .Y(n1690) );
  MUX2X1 U1341 ( .B(n1689), .A(n1674), .S(n1798), .Y(n1794) );
  MUX2X1 U1342 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1845), .Y(n1694) );
  MUX2X1 U1343 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1845), .Y(n1693) );
  MUX2X1 U1344 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1845), .Y(n1697) );
  MUX2X1 U1345 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1845), .Y(n1696) );
  MUX2X1 U1346 ( .B(n1695), .A(n1692), .S(n1803), .Y(n1706) );
  MUX2X1 U1347 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1845), .Y(n1700) );
  MUX2X1 U1348 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1845), .Y(n1699) );
  MUX2X1 U1349 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1845), .Y(n1703) );
  MUX2X1 U1350 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1845), .Y(n1702) );
  MUX2X1 U1351 ( .B(n1701), .A(n1698), .S(n1803), .Y(n1705) );
  MUX2X1 U1352 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1845), .Y(n1709) );
  MUX2X1 U1353 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1845), .Y(n1708) );
  MUX2X1 U1354 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1845), .Y(n1712) );
  MUX2X1 U1355 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1845), .Y(n1711) );
  MUX2X1 U1356 ( .B(n1710), .A(n1707), .S(n1803), .Y(n1721) );
  MUX2X1 U1357 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1846), .Y(n1715) );
  MUX2X1 U1358 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1846), .Y(n1714) );
  MUX2X1 U1359 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1846), .Y(n1718) );
  MUX2X1 U1360 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1846), .Y(n1717) );
  MUX2X1 U1361 ( .B(n1716), .A(n1713), .S(n1803), .Y(n1720) );
  MUX2X1 U1362 ( .B(n1719), .A(n1704), .S(n1798), .Y(n1795) );
  MUX2X1 U1363 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1846), .Y(n1724) );
  MUX2X1 U1364 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1846), .Y(n1723) );
  MUX2X1 U1365 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1846), .Y(n1727) );
  MUX2X1 U1366 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1846), .Y(n1726) );
  MUX2X1 U1367 ( .B(n1725), .A(n1722), .S(n1803), .Y(n1736) );
  MUX2X1 U1368 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1846), .Y(n1730) );
  MUX2X1 U1369 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1846), .Y(n1729) );
  MUX2X1 U1370 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1846), .Y(n1733) );
  MUX2X1 U1371 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1846), .Y(n1732) );
  MUX2X1 U1372 ( .B(n1731), .A(n1728), .S(n1803), .Y(n1735) );
  MUX2X1 U1373 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1847), .Y(n1739) );
  MUX2X1 U1374 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1847), .Y(n1738) );
  MUX2X1 U1375 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1847), .Y(n1742) );
  MUX2X1 U1376 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1847), .Y(n1741) );
  MUX2X1 U1377 ( .B(n1740), .A(n1737), .S(n1803), .Y(n1751) );
  MUX2X1 U1378 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1847), .Y(n1745) );
  MUX2X1 U1379 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1847), .Y(n1744) );
  MUX2X1 U1380 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1847), .Y(n1748) );
  MUX2X1 U1381 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1847), .Y(n1747) );
  MUX2X1 U1382 ( .B(n1746), .A(n1743), .S(n1803), .Y(n1750) );
  MUX2X1 U1383 ( .B(n1749), .A(n1734), .S(n1798), .Y(n1796) );
  MUX2X1 U1384 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1847), .Y(n1754) );
  MUX2X1 U1385 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1847), .Y(n1753) );
  MUX2X1 U1386 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1847), .Y(n1757) );
  MUX2X1 U1387 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1847), .Y(n1756) );
  MUX2X1 U1388 ( .B(n1755), .A(n1752), .S(n1803), .Y(n1766) );
  MUX2X1 U1389 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1848), .Y(n1760) );
  MUX2X1 U1390 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1848), .Y(n1759) );
  MUX2X1 U1391 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1848), .Y(n1763) );
  MUX2X1 U1392 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1848), .Y(n1762) );
  MUX2X1 U1393 ( .B(n1761), .A(n1758), .S(n1803), .Y(n1765) );
  MUX2X1 U1394 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1848), .Y(n1769) );
  MUX2X1 U1395 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1848), .Y(n1768) );
  MUX2X1 U1396 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1848), .Y(n1772) );
  MUX2X1 U1397 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1848), .Y(n1771) );
  MUX2X1 U1398 ( .B(n1770), .A(n1767), .S(n1803), .Y(n1781) );
  MUX2X1 U1399 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1848), .Y(n1775) );
  MUX2X1 U1400 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1848), .Y(n1774) );
  MUX2X1 U1401 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1848), .Y(n1778) );
  MUX2X1 U1402 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1848), .Y(n1777) );
  MUX2X1 U1403 ( .B(n1776), .A(n1773), .S(n1803), .Y(n1780) );
  MUX2X1 U1404 ( .B(n1779), .A(n1764), .S(n1798), .Y(n1797) );
  INVX8 U1405 ( .A(n1821), .Y(n1807) );
  INVX8 U1406 ( .A(n1821), .Y(n1808) );
  INVX8 U1407 ( .A(n1808), .Y(n1809) );
  INVX8 U1408 ( .A(n1808), .Y(n1810) );
  INVX8 U1409 ( .A(n1808), .Y(n1811) );
  INVX8 U1410 ( .A(n1807), .Y(n1812) );
  INVX8 U1411 ( .A(n1807), .Y(n1813) );
  INVX8 U1412 ( .A(n1807), .Y(n1814) );
  INVX8 U1413 ( .A(n1808), .Y(n1817) );
  INVX8 U1414 ( .A(n1808), .Y(n1818) );
  INVX8 U1415 ( .A(n1807), .Y(n1819) );
  INVX8 U1416 ( .A(n1850), .Y(n1822) );
  INVX8 U1417 ( .A(n1850), .Y(n1823) );
  INVX8 U1418 ( .A(n1850), .Y(n1824) );
  INVX8 U1419 ( .A(n1850), .Y(n1825) );
  INVX8 U1420 ( .A(n1850), .Y(n1827) );
  INVX8 U1421 ( .A(n1828), .Y(n1829) );
  INVX8 U1422 ( .A(n1828), .Y(n1830) );
  INVX8 U1423 ( .A(n1827), .Y(n1831) );
  INVX8 U1424 ( .A(n1827), .Y(n1832) );
  INVX8 U1425 ( .A(n1827), .Y(n1833) );
  INVX8 U1426 ( .A(n1826), .Y(n1834) );
  INVX8 U1427 ( .A(n1826), .Y(n1835) );
  INVX8 U1428 ( .A(n1825), .Y(n1836) );
  INVX8 U1429 ( .A(n1825), .Y(n1837) );
  INVX8 U1430 ( .A(n1825), .Y(n1838) );
  INVX8 U1431 ( .A(n1824), .Y(n1839) );
  INVX8 U1432 ( .A(n1824), .Y(n1840) );
  INVX8 U1433 ( .A(n1824), .Y(n1841) );
  INVX8 U1434 ( .A(n1823), .Y(n1842) );
  INVX8 U1435 ( .A(n1823), .Y(n1843) );
  INVX8 U1436 ( .A(n1823), .Y(n1844) );
  INVX8 U1437 ( .A(n1822), .Y(n1845) );
  INVX8 U1438 ( .A(n1822), .Y(n1846) );
  INVX8 U1439 ( .A(n1822), .Y(n1847) );
  INVX8 U1440 ( .A(n1822), .Y(n1848) );
  INVX8 U1441 ( .A(n1849), .Y(n1850) );
  INVX1 U1442 ( .A(N10), .Y(n1955) );
  INVX8 U1443 ( .A(n138), .Y(n1915) );
  INVX4 U1444 ( .A(n193), .Y(n1930) );
  INVX4 U1445 ( .A(n191), .Y(n1927) );
  INVX4 U1446 ( .A(n187), .Y(n1920) );
  INVX8 U1447 ( .A(n1915), .Y(n1914) );
  INVX8 U1448 ( .A(n185), .Y(n1917) );
  INVX8 U1449 ( .A(n1920), .Y(n1918) );
  INVX8 U1450 ( .A(n1920), .Y(n1919) );
  INVX8 U1451 ( .A(n188), .Y(n1921) );
  INVX8 U1452 ( .A(n188), .Y(n1922) );
  INVX8 U1453 ( .A(n189), .Y(n1923) );
  INVX8 U1454 ( .A(n189), .Y(n1924) );
  INVX8 U1455 ( .A(n1927), .Y(n1925) );
  INVX8 U1456 ( .A(n1927), .Y(n1926) );
  INVX8 U1457 ( .A(n1930), .Y(n1928) );
  INVX8 U1458 ( .A(n1930), .Y(n1929) );
  INVX8 U1459 ( .A(n194), .Y(n1931) );
  INVX8 U1460 ( .A(n194), .Y(n1932) );
  INVX8 U1461 ( .A(n1935), .Y(n1934) );
  INVX8 U1462 ( .A(n1938), .Y(n1936) );
  INVX8 U1463 ( .A(n1938), .Y(n1937) );
  INVX8 U1464 ( .A(n199), .Y(n1939) );
  INVX8 U1465 ( .A(n199), .Y(n1940) );
  INVX8 U1466 ( .A(n200), .Y(n1941) );
  INVX8 U1467 ( .A(n200), .Y(n1942) );
  INVX8 U1468 ( .A(n201), .Y(n1943) );
  INVX8 U1469 ( .A(n201), .Y(n1944) );
  INVX8 U1470 ( .A(n203), .Y(n1947) );
  INVX8 U1471 ( .A(n203), .Y(n1948) );
  INVX8 U1472 ( .A(n204), .Y(n1949) );
  INVX8 U1473 ( .A(n204), .Y(n1950) );
  INVX8 U1474 ( .A(n205), .Y(n1951) );
  INVX8 U1475 ( .A(n205), .Y(n1952) );
  NAND2X1 U1476 ( .A(\mem<31><0> ), .B(n117), .Y(n1964) );
  OAI21X1 U1477 ( .A(n1852), .B(n1916), .C(n1964), .Y(n2734) );
  OAI21X1 U1478 ( .A(n1918), .B(n1851), .C(n37), .Y(n2733) );
  OAI21X1 U1479 ( .A(n1922), .B(n1851), .C(n39), .Y(n2732) );
  OAI21X1 U1480 ( .A(n1924), .B(n1851), .C(n41), .Y(n2731) );
  OAI21X1 U1481 ( .A(n1925), .B(n1851), .C(n43), .Y(n2730) );
  OAI21X1 U1482 ( .A(n1928), .B(n1851), .C(n45), .Y(n2729) );
  OAI21X1 U1483 ( .A(n1932), .B(n1851), .C(n47), .Y(n2728) );
  OAI21X1 U1484 ( .A(n1934), .B(n1851), .C(n49), .Y(n2727) );
  NAND2X1 U1485 ( .A(\mem<31><8> ), .B(n117), .Y(n1965) );
  OAI21X1 U1486 ( .A(n1936), .B(n1851), .C(n1965), .Y(n2726) );
  NAND2X1 U1487 ( .A(\mem<31><9> ), .B(n117), .Y(n1966) );
  OAI21X1 U1488 ( .A(n1940), .B(n1852), .C(n1966), .Y(n2725) );
  NAND2X1 U1489 ( .A(\mem<31><10> ), .B(n117), .Y(n1967) );
  OAI21X1 U1490 ( .A(n1942), .B(n1852), .C(n1967), .Y(n2724) );
  NAND2X1 U1491 ( .A(\mem<31><11> ), .B(n117), .Y(n1968) );
  OAI21X1 U1492 ( .A(n1943), .B(n1852), .C(n1968), .Y(n2723) );
  NAND2X1 U1493 ( .A(\mem<31><12> ), .B(n117), .Y(n1969) );
  OAI21X1 U1494 ( .A(n1945), .B(n1852), .C(n1969), .Y(n2722) );
  NAND2X1 U1495 ( .A(\mem<31><13> ), .B(n117), .Y(n1970) );
  OAI21X1 U1496 ( .A(n1948), .B(n1852), .C(n1970), .Y(n2721) );
  NAND2X1 U1497 ( .A(\mem<31><14> ), .B(n117), .Y(n1971) );
  OAI21X1 U1498 ( .A(n1949), .B(n1852), .C(n1971), .Y(n2720) );
  NAND2X1 U1499 ( .A(\mem<31><15> ), .B(n117), .Y(n1972) );
  OAI21X1 U1500 ( .A(n1952), .B(n1852), .C(n1972), .Y(n2719) );
  NAND2X1 U1501 ( .A(\mem<30><0> ), .B(n183), .Y(n1973) );
  OAI21X1 U1502 ( .A(n1853), .B(n1916), .C(n1973), .Y(n2718) );
  NAND2X1 U1503 ( .A(\mem<30><1> ), .B(n490), .Y(n1974) );
  OAI21X1 U1504 ( .A(n1853), .B(n1918), .C(n1974), .Y(n2717) );
  NAND2X1 U1505 ( .A(\mem<30><2> ), .B(n1855), .Y(n1975) );
  OAI21X1 U1506 ( .A(n1853), .B(n1922), .C(n1975), .Y(n2716) );
  NAND2X1 U1507 ( .A(\mem<30><3> ), .B(n183), .Y(n1976) );
  OAI21X1 U1508 ( .A(n1853), .B(n1924), .C(n1976), .Y(n2715) );
  NAND2X1 U1509 ( .A(\mem<30><4> ), .B(n490), .Y(n1977) );
  OAI21X1 U1510 ( .A(n1853), .B(n1925), .C(n1977), .Y(n2714) );
  NAND2X1 U1511 ( .A(\mem<30><5> ), .B(n1855), .Y(n1978) );
  OAI21X1 U1512 ( .A(n1853), .B(n1928), .C(n1978), .Y(n2713) );
  NAND2X1 U1513 ( .A(\mem<30><6> ), .B(n183), .Y(n1979) );
  OAI21X1 U1514 ( .A(n1853), .B(n1932), .C(n1979), .Y(n2712) );
  NAND2X1 U1515 ( .A(\mem<30><7> ), .B(n490), .Y(n1980) );
  OAI21X1 U1516 ( .A(n1853), .B(n1934), .C(n1980), .Y(n2711) );
  NAND2X1 U1517 ( .A(\mem<30><8> ), .B(n183), .Y(n1981) );
  OAI21X1 U1518 ( .A(n1854), .B(n1937), .C(n1981), .Y(n2710) );
  NAND2X1 U1519 ( .A(\mem<30><9> ), .B(n1855), .Y(n1982) );
  OAI21X1 U1520 ( .A(n1854), .B(n1939), .C(n1982), .Y(n2709) );
  NAND2X1 U1521 ( .A(\mem<30><10> ), .B(n183), .Y(n1983) );
  OAI21X1 U1522 ( .A(n1854), .B(n1941), .C(n1983), .Y(n2708) );
  NAND2X1 U1523 ( .A(\mem<30><11> ), .B(n490), .Y(n1984) );
  OAI21X1 U1524 ( .A(n1854), .B(n1944), .C(n1984), .Y(n2707) );
  NAND2X1 U1525 ( .A(\mem<30><12> ), .B(n1855), .Y(n1985) );
  OAI21X1 U1526 ( .A(n1854), .B(n1946), .C(n1985), .Y(n2706) );
  NAND2X1 U1527 ( .A(\mem<30><13> ), .B(n183), .Y(n1986) );
  OAI21X1 U1528 ( .A(n1854), .B(n1947), .C(n1986), .Y(n2705) );
  NAND2X1 U1529 ( .A(\mem<30><14> ), .B(n490), .Y(n1987) );
  OAI21X1 U1530 ( .A(n1854), .B(n1950), .C(n1987), .Y(n2704) );
  NAND2X1 U1531 ( .A(\mem<30><15> ), .B(n1855), .Y(n1988) );
  OAI21X1 U1532 ( .A(n1854), .B(n1951), .C(n1988), .Y(n2703) );
  NAND3X1 U1533 ( .A(n1954), .B(n1958), .C(n1957), .Y(n1989) );
  NAND2X1 U1534 ( .A(\mem<29><0> ), .B(n24), .Y(n1990) );
  OAI21X1 U1535 ( .A(n1856), .B(n1917), .C(n1990), .Y(n2702) );
  NAND2X1 U1536 ( .A(\mem<29><1> ), .B(n24), .Y(n1991) );
  OAI21X1 U1537 ( .A(n1856), .B(n1918), .C(n1991), .Y(n2701) );
  NAND2X1 U1538 ( .A(\mem<29><2> ), .B(n24), .Y(n1992) );
  OAI21X1 U1539 ( .A(n1856), .B(n1921), .C(n1992), .Y(n2700) );
  NAND2X1 U1540 ( .A(\mem<29><3> ), .B(n24), .Y(n1993) );
  OAI21X1 U1541 ( .A(n1856), .B(n1923), .C(n1993), .Y(n2699) );
  NAND2X1 U1542 ( .A(\mem<29><4> ), .B(n24), .Y(n1994) );
  OAI21X1 U1543 ( .A(n1856), .B(n1925), .C(n1994), .Y(n2698) );
  NAND2X1 U1544 ( .A(\mem<29><5> ), .B(n141), .Y(n1995) );
  OAI21X1 U1545 ( .A(n1856), .B(n1928), .C(n1995), .Y(n2697) );
  NAND2X1 U1546 ( .A(\mem<29><6> ), .B(n141), .Y(n1996) );
  OAI21X1 U1547 ( .A(n1856), .B(n1931), .C(n1996), .Y(n2696) );
  NAND2X1 U1548 ( .A(\mem<29><7> ), .B(n141), .Y(n1997) );
  OAI21X1 U1549 ( .A(n1856), .B(n5), .C(n1997), .Y(n2695) );
  NAND2X1 U1550 ( .A(\mem<29><8> ), .B(n24), .Y(n1998) );
  OAI21X1 U1551 ( .A(n1857), .B(n16), .C(n1998), .Y(n2694) );
  NAND2X1 U1552 ( .A(\mem<29><9> ), .B(n140), .Y(n1999) );
  OAI21X1 U1553 ( .A(n1857), .B(n1940), .C(n1999), .Y(n2693) );
  NAND2X1 U1554 ( .A(\mem<29><10> ), .B(n24), .Y(n2000) );
  OAI21X1 U1555 ( .A(n1857), .B(n1942), .C(n2000), .Y(n2692) );
  NAND2X1 U1556 ( .A(\mem<29><11> ), .B(n140), .Y(n2001) );
  OAI21X1 U1557 ( .A(n1857), .B(n1943), .C(n2001), .Y(n2691) );
  NAND2X1 U1558 ( .A(\mem<29><12> ), .B(n24), .Y(n2002) );
  OAI21X1 U1559 ( .A(n1857), .B(n1945), .C(n2002), .Y(n2690) );
  NAND2X1 U1560 ( .A(\mem<29><13> ), .B(n140), .Y(n2003) );
  OAI21X1 U1561 ( .A(n1857), .B(n1948), .C(n2003), .Y(n2689) );
  NAND2X1 U1562 ( .A(\mem<29><14> ), .B(n141), .Y(n2004) );
  OAI21X1 U1563 ( .A(n1857), .B(n1949), .C(n2004), .Y(n2688) );
  NAND2X1 U1564 ( .A(\mem<29><15> ), .B(n140), .Y(n2005) );
  OAI21X1 U1565 ( .A(n1857), .B(n1952), .C(n2005), .Y(n2687) );
  NAND3X1 U1566 ( .A(n1958), .B(n1957), .C(n1955), .Y(n2006) );
  NAND2X1 U1567 ( .A(\mem<28><0> ), .B(n23), .Y(n2007) );
  OAI21X1 U1568 ( .A(n1858), .B(n1916), .C(n2007), .Y(n2686) );
  NAND2X1 U1569 ( .A(\mem<28><1> ), .B(n23), .Y(n2008) );
  OAI21X1 U1570 ( .A(n1858), .B(n13), .C(n2008), .Y(n2685) );
  NAND2X1 U1571 ( .A(\mem<28><2> ), .B(n23), .Y(n2009) );
  OAI21X1 U1572 ( .A(n1858), .B(n1922), .C(n2009), .Y(n2684) );
  NAND2X1 U1573 ( .A(\mem<28><3> ), .B(n23), .Y(n2010) );
  OAI21X1 U1574 ( .A(n1858), .B(n1924), .C(n2010), .Y(n2683) );
  NAND2X1 U1575 ( .A(\mem<28><4> ), .B(n23), .Y(n2011) );
  OAI21X1 U1576 ( .A(n1858), .B(n14), .C(n2011), .Y(n2682) );
  NAND2X1 U1577 ( .A(\mem<28><5> ), .B(n144), .Y(n2012) );
  OAI21X1 U1578 ( .A(n1858), .B(n15), .C(n2012), .Y(n2681) );
  NAND2X1 U1579 ( .A(\mem<28><6> ), .B(n144), .Y(n2013) );
  OAI21X1 U1580 ( .A(n1858), .B(n1932), .C(n2013), .Y(n2680) );
  NAND2X1 U1581 ( .A(\mem<28><7> ), .B(n144), .Y(n2014) );
  OAI21X1 U1582 ( .A(n1858), .B(n17), .C(n2014), .Y(n2679) );
  NAND2X1 U1583 ( .A(\mem<28><8> ), .B(n23), .Y(n2015) );
  OAI21X1 U1584 ( .A(n1859), .B(n1937), .C(n2015), .Y(n2678) );
  NAND2X1 U1585 ( .A(\mem<28><9> ), .B(n143), .Y(n2016) );
  OAI21X1 U1586 ( .A(n1859), .B(n1939), .C(n2016), .Y(n2677) );
  NAND2X1 U1587 ( .A(\mem<28><10> ), .B(n23), .Y(n2017) );
  OAI21X1 U1588 ( .A(n1859), .B(n1942), .C(n2017), .Y(n2676) );
  NAND2X1 U1589 ( .A(\mem<28><11> ), .B(n143), .Y(n2018) );
  OAI21X1 U1590 ( .A(n1859), .B(n1944), .C(n2018), .Y(n2675) );
  NAND2X1 U1591 ( .A(\mem<28><12> ), .B(n23), .Y(n2019) );
  OAI21X1 U1592 ( .A(n1859), .B(n1946), .C(n2019), .Y(n2674) );
  NAND2X1 U1593 ( .A(\mem<28><13> ), .B(n143), .Y(n2020) );
  OAI21X1 U1594 ( .A(n1859), .B(n1947), .C(n2020), .Y(n2673) );
  NAND2X1 U1595 ( .A(\mem<28><14> ), .B(n144), .Y(n2021) );
  OAI21X1 U1596 ( .A(n1859), .B(n1950), .C(n2021), .Y(n2672) );
  NAND2X1 U1597 ( .A(\mem<28><15> ), .B(n143), .Y(n2022) );
  OAI21X1 U1598 ( .A(n1859), .B(n1951), .C(n2022), .Y(n2671) );
  NAND3X1 U1599 ( .A(n1954), .B(n1956), .C(n1959), .Y(n2023) );
  NAND2X1 U1600 ( .A(\mem<27><0> ), .B(n22), .Y(n2024) );
  OAI21X1 U1601 ( .A(n1860), .B(n1917), .C(n2024), .Y(n2670) );
  NAND2X1 U1602 ( .A(\mem<27><1> ), .B(n22), .Y(n2025) );
  OAI21X1 U1603 ( .A(n1860), .B(n1919), .C(n2025), .Y(n2669) );
  NAND2X1 U1604 ( .A(\mem<27><2> ), .B(n22), .Y(n2026) );
  OAI21X1 U1605 ( .A(n1860), .B(n1921), .C(n2026), .Y(n2668) );
  NAND2X1 U1606 ( .A(\mem<27><3> ), .B(n22), .Y(n2027) );
  OAI21X1 U1607 ( .A(n1860), .B(n1923), .C(n2027), .Y(n2667) );
  NAND2X1 U1608 ( .A(\mem<27><4> ), .B(n22), .Y(n2028) );
  OAI21X1 U1609 ( .A(n1860), .B(n1926), .C(n2028), .Y(n2666) );
  NAND2X1 U1610 ( .A(\mem<27><5> ), .B(n147), .Y(n2029) );
  OAI21X1 U1611 ( .A(n1860), .B(n1929), .C(n2029), .Y(n2665) );
  NAND2X1 U1612 ( .A(\mem<27><6> ), .B(n147), .Y(n2030) );
  OAI21X1 U1613 ( .A(n1860), .B(n1931), .C(n2030), .Y(n2664) );
  NAND2X1 U1614 ( .A(\mem<27><7> ), .B(n147), .Y(n2031) );
  OAI21X1 U1615 ( .A(n1860), .B(n5), .C(n2031), .Y(n2663) );
  NAND2X1 U1616 ( .A(\mem<27><8> ), .B(n22), .Y(n2032) );
  OAI21X1 U1617 ( .A(n1861), .B(n1936), .C(n2032), .Y(n2662) );
  NAND2X1 U1618 ( .A(\mem<27><9> ), .B(n146), .Y(n2033) );
  OAI21X1 U1619 ( .A(n1861), .B(n1940), .C(n2033), .Y(n2661) );
  NAND2X1 U1620 ( .A(\mem<27><10> ), .B(n22), .Y(n2034) );
  OAI21X1 U1621 ( .A(n1861), .B(n1941), .C(n2034), .Y(n2660) );
  NAND2X1 U1622 ( .A(\mem<27><11> ), .B(n146), .Y(n2035) );
  OAI21X1 U1623 ( .A(n1861), .B(n1943), .C(n2035), .Y(n2659) );
  NAND2X1 U1624 ( .A(\mem<27><12> ), .B(n22), .Y(n2036) );
  OAI21X1 U1625 ( .A(n1861), .B(n12), .C(n2036), .Y(n2658) );
  NAND2X1 U1626 ( .A(\mem<27><13> ), .B(n146), .Y(n2037) );
  OAI21X1 U1627 ( .A(n1861), .B(n1948), .C(n2037), .Y(n2657) );
  NAND2X1 U1628 ( .A(\mem<27><14> ), .B(n147), .Y(n2038) );
  OAI21X1 U1629 ( .A(n1861), .B(n1950), .C(n2038), .Y(n2656) );
  NAND2X1 U1630 ( .A(\mem<27><15> ), .B(n146), .Y(n2039) );
  OAI21X1 U1631 ( .A(n1861), .B(n1951), .C(n2039), .Y(n2655) );
  NAND3X1 U1632 ( .A(n1959), .B(n1956), .C(n1955), .Y(n2040) );
  NAND2X1 U1633 ( .A(\mem<26><0> ), .B(n21), .Y(n2041) );
  OAI21X1 U1634 ( .A(n1862), .B(n1916), .C(n2041), .Y(n2654) );
  NAND2X1 U1635 ( .A(\mem<26><1> ), .B(n21), .Y(n2042) );
  OAI21X1 U1636 ( .A(n1862), .B(n1918), .C(n2042), .Y(n2653) );
  NAND2X1 U1637 ( .A(\mem<26><2> ), .B(n21), .Y(n2043) );
  OAI21X1 U1638 ( .A(n1862), .B(n1922), .C(n2043), .Y(n2652) );
  NAND2X1 U1639 ( .A(\mem<26><3> ), .B(n21), .Y(n2044) );
  OAI21X1 U1640 ( .A(n1862), .B(n1924), .C(n2044), .Y(n2651) );
  NAND2X1 U1641 ( .A(\mem<26><4> ), .B(n21), .Y(n2045) );
  OAI21X1 U1642 ( .A(n1862), .B(n1925), .C(n2045), .Y(n2650) );
  NAND2X1 U1643 ( .A(\mem<26><5> ), .B(n150), .Y(n2046) );
  OAI21X1 U1644 ( .A(n1862), .B(n1928), .C(n2046), .Y(n2649) );
  NAND2X1 U1645 ( .A(\mem<26><6> ), .B(n150), .Y(n2047) );
  OAI21X1 U1646 ( .A(n1862), .B(n1932), .C(n2047), .Y(n2648) );
  NAND2X1 U1647 ( .A(\mem<26><7> ), .B(n150), .Y(n2048) );
  OAI21X1 U1648 ( .A(n1862), .B(n1934), .C(n2048), .Y(n2647) );
  NAND2X1 U1649 ( .A(\mem<26><8> ), .B(n21), .Y(n2049) );
  OAI21X1 U1650 ( .A(n1863), .B(n1937), .C(n2049), .Y(n2646) );
  NAND2X1 U1651 ( .A(\mem<26><9> ), .B(n149), .Y(n2050) );
  OAI21X1 U1652 ( .A(n1863), .B(n1939), .C(n2050), .Y(n2645) );
  NAND2X1 U1653 ( .A(\mem<26><10> ), .B(n21), .Y(n2051) );
  OAI21X1 U1654 ( .A(n1863), .B(n1941), .C(n2051), .Y(n2644) );
  NAND2X1 U1655 ( .A(\mem<26><11> ), .B(n149), .Y(n2052) );
  OAI21X1 U1656 ( .A(n1863), .B(n1944), .C(n2052), .Y(n2643) );
  NAND2X1 U1657 ( .A(\mem<26><12> ), .B(n21), .Y(n2053) );
  OAI21X1 U1658 ( .A(n1863), .B(n1946), .C(n2053), .Y(n2642) );
  NAND2X1 U1659 ( .A(\mem<26><13> ), .B(n149), .Y(n2054) );
  OAI21X1 U1660 ( .A(n1863), .B(n1947), .C(n2054), .Y(n2641) );
  NAND2X1 U1661 ( .A(\mem<26><14> ), .B(n150), .Y(n2055) );
  OAI21X1 U1662 ( .A(n1863), .B(n1950), .C(n2055), .Y(n2640) );
  NAND2X1 U1663 ( .A(\mem<26><15> ), .B(n149), .Y(n2056) );
  OAI21X1 U1664 ( .A(n1863), .B(n1952), .C(n2056), .Y(n2639) );
  NAND3X1 U1665 ( .A(n1954), .B(n1959), .C(n1957), .Y(n2057) );
  NAND2X1 U1666 ( .A(\mem<25><0> ), .B(n20), .Y(n2058) );
  OAI21X1 U1667 ( .A(n1864), .B(n1917), .C(n2058), .Y(n2638) );
  NAND2X1 U1668 ( .A(\mem<25><1> ), .B(n20), .Y(n2059) );
  OAI21X1 U1669 ( .A(n1864), .B(n1919), .C(n2059), .Y(n2637) );
  NAND2X1 U1670 ( .A(\mem<25><2> ), .B(n20), .Y(n2060) );
  OAI21X1 U1671 ( .A(n1864), .B(n1921), .C(n2060), .Y(n2636) );
  NAND2X1 U1672 ( .A(\mem<25><3> ), .B(n20), .Y(n2061) );
  OAI21X1 U1673 ( .A(n1864), .B(n1923), .C(n2061), .Y(n2635) );
  NAND2X1 U1674 ( .A(\mem<25><4> ), .B(n20), .Y(n2062) );
  OAI21X1 U1675 ( .A(n1864), .B(n1926), .C(n2062), .Y(n2634) );
  NAND2X1 U1676 ( .A(\mem<25><5> ), .B(n153), .Y(n2063) );
  OAI21X1 U1677 ( .A(n1864), .B(n1929), .C(n2063), .Y(n2633) );
  NAND2X1 U1678 ( .A(\mem<25><6> ), .B(n153), .Y(n2064) );
  OAI21X1 U1679 ( .A(n1864), .B(n1931), .C(n2064), .Y(n2632) );
  NAND2X1 U1680 ( .A(\mem<25><7> ), .B(n153), .Y(n2065) );
  OAI21X1 U1681 ( .A(n1864), .B(n5), .C(n2065), .Y(n2631) );
  NAND2X1 U1682 ( .A(\mem<25><8> ), .B(n20), .Y(n2066) );
  OAI21X1 U1683 ( .A(n1865), .B(n6), .C(n2066), .Y(n2630) );
  NAND2X1 U1684 ( .A(\mem<25><9> ), .B(n152), .Y(n2067) );
  OAI21X1 U1685 ( .A(n1865), .B(n1940), .C(n2067), .Y(n2629) );
  NAND2X1 U1686 ( .A(\mem<25><10> ), .B(n20), .Y(n2068) );
  OAI21X1 U1687 ( .A(n1865), .B(n1941), .C(n2068), .Y(n2628) );
  NAND2X1 U1688 ( .A(\mem<25><11> ), .B(n152), .Y(n2069) );
  OAI21X1 U1689 ( .A(n1865), .B(n1943), .C(n2069), .Y(n2627) );
  NAND2X1 U1690 ( .A(\mem<25><12> ), .B(n20), .Y(n2070) );
  OAI21X1 U1691 ( .A(n1865), .B(n12), .C(n2070), .Y(n2626) );
  NAND2X1 U1692 ( .A(\mem<25><13> ), .B(n152), .Y(n2071) );
  OAI21X1 U1693 ( .A(n1865), .B(n1948), .C(n2071), .Y(n2625) );
  NAND2X1 U1694 ( .A(\mem<25><14> ), .B(n153), .Y(n2072) );
  OAI21X1 U1695 ( .A(n1865), .B(n1950), .C(n2072), .Y(n2624) );
  NAND2X1 U1696 ( .A(\mem<25><15> ), .B(n152), .Y(n2073) );
  OAI21X1 U1697 ( .A(n1865), .B(n1952), .C(n2073), .Y(n2623) );
  NOR3X1 U1698 ( .A(n1954), .B(n1956), .C(n1958), .Y(n2206) );
  NAND2X1 U1699 ( .A(\mem<24><0> ), .B(n25), .Y(n2074) );
  OAI21X1 U1700 ( .A(n1866), .B(n1916), .C(n2074), .Y(n2622) );
  NAND2X1 U1701 ( .A(\mem<24><1> ), .B(n25), .Y(n2075) );
  OAI21X1 U1702 ( .A(n1866), .B(n10), .C(n2075), .Y(n2621) );
  NAND2X1 U1703 ( .A(\mem<24><2> ), .B(n156), .Y(n2076) );
  OAI21X1 U1704 ( .A(n1866), .B(n1921), .C(n2076), .Y(n2620) );
  NAND2X1 U1705 ( .A(\mem<24><3> ), .B(n156), .Y(n2077) );
  OAI21X1 U1706 ( .A(n1866), .B(n1923), .C(n2077), .Y(n2619) );
  NAND2X1 U1707 ( .A(\mem<24><4> ), .B(n25), .Y(n2078) );
  OAI21X1 U1708 ( .A(n1866), .B(n8), .C(n2078), .Y(n2618) );
  NAND2X1 U1709 ( .A(\mem<24><5> ), .B(n25), .Y(n2079) );
  OAI21X1 U1710 ( .A(n1866), .B(n9), .C(n2079), .Y(n2617) );
  NAND2X1 U1711 ( .A(\mem<24><6> ), .B(n156), .Y(n2080) );
  OAI21X1 U1712 ( .A(n1866), .B(n1931), .C(n2080), .Y(n2616) );
  NAND2X1 U1713 ( .A(\mem<24><7> ), .B(n156), .Y(n2081) );
  OAI21X1 U1714 ( .A(n1866), .B(n1933), .C(n2081), .Y(n2615) );
  NAND2X1 U1715 ( .A(\mem<24><8> ), .B(n155), .Y(n2082) );
  OAI21X1 U1716 ( .A(n1866), .B(n1936), .C(n2082), .Y(n2614) );
  NAND2X1 U1717 ( .A(\mem<24><9> ), .B(n25), .Y(n2083) );
  OAI21X1 U1718 ( .A(n1866), .B(n1939), .C(n2083), .Y(n2613) );
  NAND2X1 U1719 ( .A(\mem<24><10> ), .B(n155), .Y(n2084) );
  OAI21X1 U1720 ( .A(n1866), .B(n1942), .C(n2084), .Y(n2612) );
  NAND2X1 U1721 ( .A(\mem<24><11> ), .B(n25), .Y(n2085) );
  OAI21X1 U1722 ( .A(n1866), .B(n1944), .C(n2085), .Y(n2611) );
  NAND2X1 U1723 ( .A(\mem<24><12> ), .B(n155), .Y(n2086) );
  OAI21X1 U1724 ( .A(n1866), .B(n1945), .C(n2086), .Y(n2610) );
  NAND2X1 U1725 ( .A(\mem<24><13> ), .B(n25), .Y(n2087) );
  OAI21X1 U1726 ( .A(n1866), .B(n1947), .C(n2087), .Y(n2609) );
  NAND2X1 U1727 ( .A(\mem<24><14> ), .B(n155), .Y(n2088) );
  OAI21X1 U1728 ( .A(n1866), .B(n1950), .C(n2088), .Y(n2608) );
  NAND2X1 U1729 ( .A(\mem<24><15> ), .B(n25), .Y(n2089) );
  OAI21X1 U1730 ( .A(n1866), .B(n1951), .C(n2089), .Y(n2607) );
  NAND2X1 U1731 ( .A(\mem<23><0> ), .B(n19), .Y(n2090) );
  OAI21X1 U1732 ( .A(n1867), .B(n1917), .C(n2090), .Y(n2606) );
  NAND2X1 U1733 ( .A(\mem<23><1> ), .B(n19), .Y(n2091) );
  OAI21X1 U1734 ( .A(n1867), .B(n13), .C(n2091), .Y(n2605) );
  NAND2X1 U1735 ( .A(\mem<23><2> ), .B(n19), .Y(n2092) );
  OAI21X1 U1736 ( .A(n1867), .B(n1922), .C(n2092), .Y(n2604) );
  NAND2X1 U1737 ( .A(\mem<23><3> ), .B(n19), .Y(n2093) );
  OAI21X1 U1738 ( .A(n1867), .B(n1924), .C(n2093), .Y(n2603) );
  NAND2X1 U1739 ( .A(\mem<23><4> ), .B(n19), .Y(n2094) );
  OAI21X1 U1740 ( .A(n1867), .B(n14), .C(n2094), .Y(n2602) );
  NAND2X1 U1741 ( .A(\mem<23><5> ), .B(n159), .Y(n2095) );
  OAI21X1 U1742 ( .A(n1867), .B(n15), .C(n2095), .Y(n2601) );
  NAND2X1 U1743 ( .A(\mem<23><6> ), .B(n159), .Y(n2096) );
  OAI21X1 U1744 ( .A(n1867), .B(n1932), .C(n2096), .Y(n2600) );
  NAND2X1 U1745 ( .A(\mem<23><7> ), .B(n159), .Y(n2097) );
  OAI21X1 U1746 ( .A(n1867), .B(n17), .C(n2097), .Y(n2599) );
  NAND2X1 U1747 ( .A(\mem<23><8> ), .B(n19), .Y(n2098) );
  OAI21X1 U1748 ( .A(n1868), .B(n1936), .C(n2098), .Y(n2598) );
  NAND2X1 U1749 ( .A(\mem<23><9> ), .B(n158), .Y(n2099) );
  OAI21X1 U1750 ( .A(n1868), .B(n1940), .C(n2099), .Y(n2597) );
  NAND2X1 U1751 ( .A(\mem<23><10> ), .B(n19), .Y(n2100) );
  OAI21X1 U1752 ( .A(n1868), .B(n1942), .C(n2100), .Y(n2596) );
  NAND2X1 U1753 ( .A(\mem<23><11> ), .B(n158), .Y(n2101) );
  OAI21X1 U1754 ( .A(n1868), .B(n1943), .C(n2101), .Y(n2595) );
  NAND2X1 U1755 ( .A(\mem<23><12> ), .B(n19), .Y(n2102) );
  OAI21X1 U1756 ( .A(n1868), .B(n1945), .C(n2102), .Y(n2594) );
  NAND2X1 U1757 ( .A(\mem<23><13> ), .B(n158), .Y(n2103) );
  OAI21X1 U1758 ( .A(n1868), .B(n1948), .C(n2103), .Y(n2593) );
  NAND2X1 U1759 ( .A(\mem<23><14> ), .B(n159), .Y(n2104) );
  OAI21X1 U1760 ( .A(n1868), .B(n1949), .C(n2104), .Y(n2592) );
  NAND2X1 U1761 ( .A(\mem<23><15> ), .B(n158), .Y(n2105) );
  OAI21X1 U1762 ( .A(n1868), .B(n1951), .C(n2105), .Y(n2591) );
  NAND2X1 U1763 ( .A(\mem<22><0> ), .B(n119), .Y(n2106) );
  OAI21X1 U1764 ( .A(n1869), .B(n1917), .C(n2106), .Y(n2590) );
  NAND2X1 U1765 ( .A(\mem<22><1> ), .B(n119), .Y(n2107) );
  OAI21X1 U1766 ( .A(n1869), .B(n1918), .C(n2107), .Y(n2589) );
  NAND2X1 U1767 ( .A(\mem<22><2> ), .B(n119), .Y(n2108) );
  OAI21X1 U1768 ( .A(n1869), .B(n1922), .C(n2108), .Y(n2588) );
  NAND2X1 U1769 ( .A(\mem<22><3> ), .B(n119), .Y(n2109) );
  OAI21X1 U1770 ( .A(n1869), .B(n1924), .C(n2109), .Y(n2587) );
  NAND2X1 U1771 ( .A(\mem<22><4> ), .B(n119), .Y(n2110) );
  OAI21X1 U1772 ( .A(n1869), .B(n1925), .C(n2110), .Y(n2586) );
  NAND2X1 U1773 ( .A(\mem<22><5> ), .B(n119), .Y(n2111) );
  OAI21X1 U1774 ( .A(n1869), .B(n1928), .C(n2111), .Y(n2585) );
  NAND2X1 U1775 ( .A(\mem<22><6> ), .B(n119), .Y(n2112) );
  OAI21X1 U1776 ( .A(n1869), .B(n1932), .C(n2112), .Y(n2584) );
  NAND2X1 U1777 ( .A(\mem<22><7> ), .B(n119), .Y(n2113) );
  OAI21X1 U1778 ( .A(n1869), .B(n1934), .C(n2113), .Y(n2583) );
  OAI21X1 U1779 ( .A(n1870), .B(n6), .C(n51), .Y(n2582) );
  OAI21X1 U1780 ( .A(n1870), .B(n1940), .C(n53), .Y(n2581) );
  OAI21X1 U1781 ( .A(n1870), .B(n1942), .C(n55), .Y(n2580) );
  OAI21X1 U1782 ( .A(n1870), .B(n1943), .C(n57), .Y(n2579) );
  OAI21X1 U1783 ( .A(n1870), .B(n1945), .C(n59), .Y(n2578) );
  OAI21X1 U1784 ( .A(n1870), .B(n1948), .C(n61), .Y(n2577) );
  OAI21X1 U1785 ( .A(n1870), .B(n1949), .C(n63), .Y(n2576) );
  NAND2X1 U1786 ( .A(\mem<22><15> ), .B(n119), .Y(n2114) );
  OAI21X1 U1787 ( .A(n1870), .B(n1952), .C(n2114), .Y(n2575) );
  NAND2X1 U1788 ( .A(\mem<21><0> ), .B(n121), .Y(n2115) );
  OAI21X1 U1789 ( .A(n1871), .B(n1917), .C(n2115), .Y(n2574) );
  NAND2X1 U1790 ( .A(\mem<21><1> ), .B(n121), .Y(n2116) );
  OAI21X1 U1791 ( .A(n1871), .B(n1919), .C(n2116), .Y(n2573) );
  NAND2X1 U1792 ( .A(\mem<21><2> ), .B(n121), .Y(n2117) );
  OAI21X1 U1793 ( .A(n1871), .B(n1922), .C(n2117), .Y(n2572) );
  NAND2X1 U1794 ( .A(\mem<21><3> ), .B(n121), .Y(n2118) );
  OAI21X1 U1795 ( .A(n1871), .B(n1924), .C(n2118), .Y(n2571) );
  NAND2X1 U1796 ( .A(\mem<21><4> ), .B(n121), .Y(n2119) );
  OAI21X1 U1797 ( .A(n1871), .B(n1926), .C(n2119), .Y(n2570) );
  NAND2X1 U1798 ( .A(\mem<21><5> ), .B(n121), .Y(n2120) );
  OAI21X1 U1799 ( .A(n1871), .B(n1929), .C(n2120), .Y(n2569) );
  NAND2X1 U1800 ( .A(\mem<21><6> ), .B(n121), .Y(n2121) );
  OAI21X1 U1801 ( .A(n1871), .B(n1932), .C(n2121), .Y(n2568) );
  NAND2X1 U1802 ( .A(\mem<21><7> ), .B(n121), .Y(n2122) );
  OAI21X1 U1803 ( .A(n1871), .B(n17), .C(n2122), .Y(n2567) );
  OAI21X1 U1804 ( .A(n1872), .B(n1936), .C(n65), .Y(n2566) );
  OAI21X1 U1805 ( .A(n1872), .B(n1940), .C(n67), .Y(n2565) );
  OAI21X1 U1806 ( .A(n1872), .B(n1941), .C(n69), .Y(n2564) );
  OAI21X1 U1807 ( .A(n1872), .B(n1943), .C(n71), .Y(n2563) );
  OAI21X1 U1808 ( .A(n1872), .B(n12), .C(n73), .Y(n2562) );
  OAI21X1 U1809 ( .A(n1872), .B(n1948), .C(n75), .Y(n2561) );
  OAI21X1 U1810 ( .A(n1872), .B(n1949), .C(n77), .Y(n2560) );
  NAND2X1 U1811 ( .A(\mem<21><15> ), .B(n121), .Y(n2123) );
  OAI21X1 U1812 ( .A(n1872), .B(n1951), .C(n2123), .Y(n2559) );
  NAND2X1 U1813 ( .A(\mem<20><0> ), .B(n123), .Y(n2124) );
  OAI21X1 U1814 ( .A(n1873), .B(n1916), .C(n2124), .Y(n2558) );
  NAND2X1 U1815 ( .A(\mem<20><1> ), .B(n123), .Y(n2125) );
  OAI21X1 U1816 ( .A(n1873), .B(n13), .C(n2125), .Y(n2557) );
  NAND2X1 U1817 ( .A(\mem<20><2> ), .B(n123), .Y(n2126) );
  OAI21X1 U1818 ( .A(n1873), .B(n1922), .C(n2126), .Y(n2556) );
  NAND2X1 U1819 ( .A(\mem<20><3> ), .B(n123), .Y(n2127) );
  OAI21X1 U1820 ( .A(n1873), .B(n1924), .C(n2127), .Y(n2555) );
  NAND2X1 U1821 ( .A(\mem<20><4> ), .B(n123), .Y(n2128) );
  OAI21X1 U1822 ( .A(n1873), .B(n14), .C(n2128), .Y(n2554) );
  NAND2X1 U1823 ( .A(\mem<20><5> ), .B(n123), .Y(n2129) );
  OAI21X1 U1824 ( .A(n1873), .B(n15), .C(n2129), .Y(n2553) );
  NAND2X1 U1825 ( .A(\mem<20><6> ), .B(n123), .Y(n2130) );
  OAI21X1 U1826 ( .A(n1873), .B(n1932), .C(n2130), .Y(n2552) );
  NAND2X1 U1827 ( .A(\mem<20><7> ), .B(n123), .Y(n2131) );
  OAI21X1 U1828 ( .A(n1873), .B(n1934), .C(n2131), .Y(n2551) );
  OAI21X1 U1829 ( .A(n1874), .B(n6), .C(n79), .Y(n2550) );
  OAI21X1 U1830 ( .A(n1874), .B(n1940), .C(n81), .Y(n2549) );
  OAI21X1 U1831 ( .A(n1874), .B(n1942), .C(n83), .Y(n2548) );
  OAI21X1 U1832 ( .A(n1874), .B(n1943), .C(n85), .Y(n2547) );
  OAI21X1 U1833 ( .A(n1874), .B(n12), .C(n87), .Y(n2546) );
  OAI21X1 U1834 ( .A(n1874), .B(n1948), .C(n89), .Y(n2545) );
  OAI21X1 U1835 ( .A(n1874), .B(n1950), .C(n91), .Y(n2544) );
  NAND2X1 U1836 ( .A(\mem<20><15> ), .B(n123), .Y(n2132) );
  OAI21X1 U1837 ( .A(n1874), .B(n1952), .C(n2132), .Y(n2543) );
  OAI21X1 U1838 ( .A(n1875), .B(n1916), .C(n494), .Y(n2542) );
  OAI21X1 U1839 ( .A(n1875), .B(n13), .C(n208), .Y(n2541) );
  OAI21X1 U1840 ( .A(n1875), .B(n1922), .C(n210), .Y(n2540) );
  OAI21X1 U1841 ( .A(n1875), .B(n1924), .C(n212), .Y(n2539) );
  OAI21X1 U1842 ( .A(n1875), .B(n14), .C(n215), .Y(n2538) );
  OAI21X1 U1843 ( .A(n1875), .B(n15), .C(n217), .Y(n2537) );
  OAI21X1 U1844 ( .A(n1875), .B(n1932), .C(n219), .Y(n2536) );
  OAI21X1 U1845 ( .A(n1875), .B(n17), .C(n221), .Y(n2535) );
  OAI21X1 U1846 ( .A(n1876), .B(n1936), .C(n496), .Y(n2534) );
  OAI21X1 U1847 ( .A(n1876), .B(n1940), .C(n498), .Y(n2533) );
  OAI21X1 U1848 ( .A(n1876), .B(n1941), .C(n500), .Y(n2532) );
  OAI21X1 U1849 ( .A(n1876), .B(n1943), .C(n502), .Y(n2531) );
  OAI21X1 U1850 ( .A(n1876), .B(n1945), .C(n504), .Y(n2530) );
  OAI21X1 U1851 ( .A(n1876), .B(n1948), .C(n506), .Y(n2529) );
  OAI21X1 U1852 ( .A(n1876), .B(n1949), .C(n508), .Y(n2528) );
  OAI21X1 U1853 ( .A(n1876), .B(n1951), .C(n510), .Y(n2527) );
  OAI21X1 U1854 ( .A(n1877), .B(n1917), .C(n512), .Y(n2526) );
  OAI21X1 U1855 ( .A(n1877), .B(n1919), .C(n223), .Y(n2525) );
  OAI21X1 U1856 ( .A(n1877), .B(n1922), .C(n225), .Y(n2524) );
  OAI21X1 U1857 ( .A(n1877), .B(n1924), .C(n227), .Y(n2523) );
  OAI21X1 U1858 ( .A(n1877), .B(n1926), .C(n229), .Y(n2522) );
  OAI21X1 U1859 ( .A(n1877), .B(n1929), .C(n231), .Y(n2521) );
  OAI21X1 U1860 ( .A(n1877), .B(n1932), .C(n233), .Y(n2520) );
  OAI21X1 U1861 ( .A(n1877), .B(n1934), .C(n235), .Y(n2519) );
  OAI21X1 U1862 ( .A(n1878), .B(n16), .C(n514), .Y(n2518) );
  OAI21X1 U1863 ( .A(n1878), .B(n1940), .C(n516), .Y(n2517) );
  OAI21X1 U1864 ( .A(n1878), .B(n1941), .C(n518), .Y(n2516) );
  OAI21X1 U1865 ( .A(n1878), .B(n1943), .C(n520), .Y(n2515) );
  OAI21X1 U1866 ( .A(n1878), .B(n1945), .C(n522), .Y(n2514) );
  OAI21X1 U1867 ( .A(n1878), .B(n1948), .C(n524), .Y(n2513) );
  OAI21X1 U1868 ( .A(n1878), .B(n1949), .C(n526), .Y(n2512) );
  OAI21X1 U1869 ( .A(n1878), .B(n1952), .C(n528), .Y(n2511) );
  OAI21X1 U1870 ( .A(n1879), .B(n1916), .C(n530), .Y(n2510) );
  OAI21X1 U1871 ( .A(n1879), .B(n1918), .C(n237), .Y(n2509) );
  OAI21X1 U1872 ( .A(n1879), .B(n1922), .C(n239), .Y(n2508) );
  OAI21X1 U1873 ( .A(n1879), .B(n1924), .C(n241), .Y(n2507) );
  OAI21X1 U1874 ( .A(n1879), .B(n1925), .C(n243), .Y(n2506) );
  OAI21X1 U1875 ( .A(n1879), .B(n1928), .C(n245), .Y(n2505) );
  OAI21X1 U1876 ( .A(n1879), .B(n1932), .C(n247), .Y(n2504) );
  OAI21X1 U1877 ( .A(n1879), .B(n17), .C(n249), .Y(n2503) );
  OAI21X1 U1878 ( .A(n1880), .B(n1936), .C(n532), .Y(n2502) );
  OAI21X1 U1879 ( .A(n1880), .B(n1940), .C(n534), .Y(n2501) );
  OAI21X1 U1880 ( .A(n1880), .B(n1942), .C(n536), .Y(n2500) );
  OAI21X1 U1881 ( .A(n1880), .B(n1944), .C(n538), .Y(n2499) );
  OAI21X1 U1882 ( .A(n1880), .B(n1945), .C(n540), .Y(n2498) );
  OAI21X1 U1883 ( .A(n1880), .B(n1948), .C(n542), .Y(n2497) );
  OAI21X1 U1884 ( .A(n1880), .B(n1949), .C(n544), .Y(n2496) );
  OAI21X1 U1885 ( .A(n1880), .B(n1951), .C(n546), .Y(n2495) );
  OAI21X1 U1886 ( .A(n1881), .B(n1916), .C(n548), .Y(n2494) );
  OAI21X1 U1887 ( .A(n1881), .B(n10), .C(n251), .Y(n2493) );
  OAI21X1 U1888 ( .A(n1881), .B(n1922), .C(n253), .Y(n2492) );
  OAI21X1 U1889 ( .A(n1881), .B(n1924), .C(n255), .Y(n2491) );
  OAI21X1 U1890 ( .A(n1881), .B(n8), .C(n257), .Y(n2490) );
  OAI21X1 U1891 ( .A(n1881), .B(n9), .C(n259), .Y(n2489) );
  OAI21X1 U1892 ( .A(n1881), .B(n1932), .C(n261), .Y(n2488) );
  OAI21X1 U1893 ( .A(n1881), .B(n1933), .C(n263), .Y(n2487) );
  OAI21X1 U1894 ( .A(n1881), .B(n11), .C(n550), .Y(n2486) );
  OAI21X1 U1895 ( .A(n1881), .B(n1940), .C(n552), .Y(n2485) );
  OAI21X1 U1896 ( .A(n1881), .B(n1941), .C(n554), .Y(n2484) );
  OAI21X1 U1897 ( .A(n1881), .B(n1943), .C(n556), .Y(n2483) );
  OAI21X1 U1898 ( .A(n1881), .B(n1946), .C(n558), .Y(n2482) );
  OAI21X1 U1899 ( .A(n1881), .B(n1948), .C(n560), .Y(n2481) );
  OAI21X1 U1900 ( .A(n1881), .B(n1949), .C(n562), .Y(n2480) );
  OAI21X1 U1901 ( .A(n1881), .B(n1952), .C(n564), .Y(n2479) );
  NAND3X1 U1902 ( .A(n1960), .B(n2735), .C(n1963), .Y(n2133) );
  OAI21X1 U1903 ( .A(n1882), .B(n1917), .C(n566), .Y(n2478) );
  OAI21X1 U1904 ( .A(n1882), .B(n1919), .C(n265), .Y(n2477) );
  OAI21X1 U1905 ( .A(n1882), .B(n1922), .C(n267), .Y(n2476) );
  OAI21X1 U1906 ( .A(n1882), .B(n1924), .C(n269), .Y(n2475) );
  OAI21X1 U1907 ( .A(n1882), .B(n1926), .C(n271), .Y(n2474) );
  OAI21X1 U1908 ( .A(n1882), .B(n1929), .C(n273), .Y(n2473) );
  OAI21X1 U1909 ( .A(n1882), .B(n1932), .C(n275), .Y(n2472) );
  OAI21X1 U1910 ( .A(n1882), .B(n1934), .C(n277), .Y(n2471) );
  OAI21X1 U1911 ( .A(n1883), .B(n6), .C(n568), .Y(n2470) );
  OAI21X1 U1912 ( .A(n1883), .B(n1940), .C(n570), .Y(n2469) );
  OAI21X1 U1913 ( .A(n1883), .B(n1942), .C(n572), .Y(n2468) );
  OAI21X1 U1914 ( .A(n1883), .B(n1944), .C(n574), .Y(n2467) );
  OAI21X1 U1915 ( .A(n1883), .B(n12), .C(n576), .Y(n2466) );
  OAI21X1 U1916 ( .A(n1883), .B(n1948), .C(n578), .Y(n2465) );
  OAI21X1 U1917 ( .A(n1883), .B(n1950), .C(n580), .Y(n2464) );
  OAI21X1 U1918 ( .A(n1883), .B(n1952), .C(n582), .Y(n2463) );
  OAI21X1 U1919 ( .A(n1884), .B(n1916), .C(n584), .Y(n2462) );
  OAI21X1 U1920 ( .A(n1884), .B(n1919), .C(n279), .Y(n2461) );
  OAI21X1 U1921 ( .A(n1884), .B(n1922), .C(n281), .Y(n2460) );
  OAI21X1 U1922 ( .A(n1884), .B(n1924), .C(n283), .Y(n2459) );
  OAI21X1 U1923 ( .A(n1884), .B(n1926), .C(n285), .Y(n2458) );
  OAI21X1 U1924 ( .A(n1884), .B(n1929), .C(n287), .Y(n2457) );
  OAI21X1 U1925 ( .A(n1884), .B(n1932), .C(n289), .Y(n2456) );
  OAI21X1 U1926 ( .A(n1884), .B(n17), .C(n291), .Y(n2455) );
  OAI21X1 U1927 ( .A(n1885), .B(n1936), .C(n586), .Y(n2454) );
  OAI21X1 U1928 ( .A(n1885), .B(n1940), .C(n588), .Y(n2453) );
  OAI21X1 U1929 ( .A(n1885), .B(n1941), .C(n590), .Y(n2452) );
  OAI21X1 U1930 ( .A(n1885), .B(n1943), .C(n592), .Y(n2451) );
  OAI21X1 U1931 ( .A(n1885), .B(n1945), .C(n594), .Y(n2450) );
  OAI21X1 U1932 ( .A(n1885), .B(n1948), .C(n596), .Y(n2449) );
  OAI21X1 U1933 ( .A(n1885), .B(n1949), .C(n598), .Y(n2448) );
  OAI21X1 U1934 ( .A(n1885), .B(n1951), .C(n600), .Y(n2447) );
  OAI21X1 U1935 ( .A(n1886), .B(n1917), .C(n602), .Y(n2446) );
  OAI21X1 U1936 ( .A(n1886), .B(n1918), .C(n293), .Y(n2445) );
  OAI21X1 U1937 ( .A(n1886), .B(n1922), .C(n295), .Y(n2444) );
  OAI21X1 U1938 ( .A(n1886), .B(n1924), .C(n297), .Y(n2443) );
  OAI21X1 U1939 ( .A(n1886), .B(n1925), .C(n299), .Y(n2442) );
  OAI21X1 U1940 ( .A(n1886), .B(n1928), .C(n301), .Y(n2441) );
  OAI21X1 U1941 ( .A(n1886), .B(n1932), .C(n303), .Y(n2440) );
  OAI21X1 U1942 ( .A(n1886), .B(n1934), .C(n305), .Y(n2439) );
  OAI21X1 U1943 ( .A(n1887), .B(n6), .C(n604), .Y(n2438) );
  OAI21X1 U1944 ( .A(n1887), .B(n1940), .C(n606), .Y(n2437) );
  OAI21X1 U1945 ( .A(n1887), .B(n1942), .C(n608), .Y(n2436) );
  OAI21X1 U1946 ( .A(n1887), .B(n1943), .C(n610), .Y(n2435) );
  OAI21X1 U1947 ( .A(n1887), .B(n1945), .C(n612), .Y(n2434) );
  OAI21X1 U1948 ( .A(n1887), .B(n1948), .C(n614), .Y(n2433) );
  OAI21X1 U1949 ( .A(n1887), .B(n1949), .C(n616), .Y(n2432) );
  OAI21X1 U1950 ( .A(n1887), .B(n1952), .C(n618), .Y(n2431) );
  OAI21X1 U1951 ( .A(n1888), .B(n1916), .C(n620), .Y(n2430) );
  OAI21X1 U1952 ( .A(n1888), .B(n1919), .C(n307), .Y(n2429) );
  OAI21X1 U1953 ( .A(n1888), .B(n1922), .C(n309), .Y(n2428) );
  OAI21X1 U1954 ( .A(n1888), .B(n1924), .C(n311), .Y(n2427) );
  OAI21X1 U1955 ( .A(n1888), .B(n1926), .C(n313), .Y(n2426) );
  OAI21X1 U1956 ( .A(n1888), .B(n1929), .C(n315), .Y(n2425) );
  OAI21X1 U1957 ( .A(n1888), .B(n1932), .C(n317), .Y(n2424) );
  OAI21X1 U1958 ( .A(n1888), .B(n17), .C(n319), .Y(n2423) );
  OAI21X1 U1959 ( .A(n1889), .B(n1936), .C(n622), .Y(n2422) );
  OAI21X1 U1960 ( .A(n1889), .B(n1940), .C(n624), .Y(n2421) );
  OAI21X1 U1961 ( .A(n1889), .B(n1941), .C(n626), .Y(n2420) );
  OAI21X1 U1962 ( .A(n1889), .B(n1944), .C(n628), .Y(n2419) );
  OAI21X1 U1963 ( .A(n1889), .B(n12), .C(n630), .Y(n2418) );
  OAI21X1 U1964 ( .A(n1889), .B(n1948), .C(n632), .Y(n2417) );
  OAI21X1 U1965 ( .A(n1889), .B(n1949), .C(n634), .Y(n2416) );
  OAI21X1 U1966 ( .A(n1889), .B(n1951), .C(n636), .Y(n2415) );
  OAI21X1 U1967 ( .A(n1890), .B(n1917), .C(n638), .Y(n2414) );
  OAI21X1 U1968 ( .A(n1890), .B(n13), .C(n321), .Y(n2413) );
  OAI21X1 U1969 ( .A(n1890), .B(n1921), .C(n323), .Y(n2412) );
  OAI21X1 U1970 ( .A(n1890), .B(n1923), .C(n325), .Y(n2411) );
  OAI21X1 U1971 ( .A(n1890), .B(n14), .C(n327), .Y(n2410) );
  OAI21X1 U1972 ( .A(n1890), .B(n15), .C(n329), .Y(n2409) );
  OAI21X1 U1973 ( .A(n1890), .B(n1931), .C(n331), .Y(n2408) );
  OAI21X1 U1974 ( .A(n1890), .B(n5), .C(n333), .Y(n2407) );
  OAI21X1 U1975 ( .A(n1891), .B(n1937), .C(n640), .Y(n2406) );
  OAI21X1 U1976 ( .A(n1891), .B(n1939), .C(n642), .Y(n2405) );
  OAI21X1 U1977 ( .A(n1891), .B(n1941), .C(n644), .Y(n2404) );
  OAI21X1 U1978 ( .A(n1891), .B(n1944), .C(n646), .Y(n2403) );
  OAI21X1 U1979 ( .A(n1891), .B(n1946), .C(n648), .Y(n2402) );
  OAI21X1 U1980 ( .A(n1891), .B(n1947), .C(n650), .Y(n2401) );
  OAI21X1 U1981 ( .A(n1891), .B(n1950), .C(n1164), .Y(n2400) );
  OAI21X1 U1982 ( .A(n1891), .B(n1951), .C(n1166), .Y(n2399) );
  OAI21X1 U1983 ( .A(n1892), .B(n1916), .C(n1168), .Y(n2398) );
  OAI21X1 U1984 ( .A(n1892), .B(n1919), .C(n335), .Y(n2397) );
  OAI21X1 U1985 ( .A(n1892), .B(n1921), .C(n337), .Y(n2396) );
  OAI21X1 U1986 ( .A(n1892), .B(n1923), .C(n339), .Y(n2395) );
  OAI21X1 U1987 ( .A(n1892), .B(n1926), .C(n341), .Y(n2394) );
  OAI21X1 U1988 ( .A(n1892), .B(n1929), .C(n343), .Y(n2393) );
  OAI21X1 U1989 ( .A(n1892), .B(n1931), .C(n345), .Y(n2392) );
  OAI21X1 U1990 ( .A(n1892), .B(n7), .C(n347), .Y(n2391) );
  OAI21X1 U1991 ( .A(n1893), .B(n1937), .C(n1170), .Y(n2390) );
  OAI21X1 U1992 ( .A(n1893), .B(n1939), .C(n1172), .Y(n2389) );
  OAI21X1 U1993 ( .A(n1893), .B(n1942), .C(n1174), .Y(n2388) );
  OAI21X1 U1994 ( .A(n1893), .B(n1944), .C(n1176), .Y(n2387) );
  OAI21X1 U1995 ( .A(n1893), .B(n1946), .C(n1178), .Y(n2386) );
  OAI21X1 U1996 ( .A(n1893), .B(n1947), .C(n1180), .Y(n2385) );
  OAI21X1 U1997 ( .A(n1893), .B(n1950), .C(n1182), .Y(n2384) );
  OAI21X1 U1998 ( .A(n1893), .B(n1952), .C(n1184), .Y(n2383) );
  OAI21X1 U1999 ( .A(n1894), .B(n1917), .C(n1186), .Y(n2382) );
  OAI21X1 U2000 ( .A(n1894), .B(n13), .C(n349), .Y(n2381) );
  OAI21X1 U2001 ( .A(n1894), .B(n1921), .C(n351), .Y(n2380) );
  OAI21X1 U2002 ( .A(n1894), .B(n1923), .C(n353), .Y(n2379) );
  OAI21X1 U2003 ( .A(n1894), .B(n14), .C(n355), .Y(n2378) );
  OAI21X1 U2004 ( .A(n1894), .B(n15), .C(n357), .Y(n2377) );
  OAI21X1 U2005 ( .A(n1894), .B(n1931), .C(n359), .Y(n2376) );
  OAI21X1 U2006 ( .A(n1894), .B(n7), .C(n361), .Y(n2375) );
  OAI21X1 U2007 ( .A(n1895), .B(n1937), .C(n1188), .Y(n2374) );
  OAI21X1 U2008 ( .A(n1895), .B(n1939), .C(n1190), .Y(n2373) );
  OAI21X1 U2009 ( .A(n1895), .B(n1942), .C(n1192), .Y(n2372) );
  OAI21X1 U2010 ( .A(n1895), .B(n1944), .C(n1194), .Y(n2371) );
  OAI21X1 U2011 ( .A(n1895), .B(n1946), .C(n1196), .Y(n2370) );
  OAI21X1 U2012 ( .A(n1895), .B(n1947), .C(n1198), .Y(n2369) );
  OAI21X1 U2013 ( .A(n1895), .B(n1950), .C(n1200), .Y(n2368) );
  OAI21X1 U2014 ( .A(n1895), .B(n1951), .C(n1202), .Y(n2367) );
  NAND2X1 U2015 ( .A(\mem<8><0> ), .B(n93), .Y(n2135) );
  OAI21X1 U2016 ( .A(n1896), .B(n1916), .C(n2135), .Y(n2366) );
  NAND2X1 U2017 ( .A(\mem<8><1> ), .B(n93), .Y(n2136) );
  OAI21X1 U2018 ( .A(n1896), .B(n13), .C(n2136), .Y(n2365) );
  NAND2X1 U2019 ( .A(\mem<8><2> ), .B(n93), .Y(n2137) );
  OAI21X1 U2020 ( .A(n1896), .B(n1921), .C(n2137), .Y(n2364) );
  NAND2X1 U2021 ( .A(\mem<8><3> ), .B(n93), .Y(n2138) );
  OAI21X1 U2022 ( .A(n1896), .B(n1923), .C(n2138), .Y(n2363) );
  NAND2X1 U2023 ( .A(\mem<8><4> ), .B(n93), .Y(n2139) );
  OAI21X1 U2024 ( .A(n1896), .B(n14), .C(n2139), .Y(n2362) );
  NAND2X1 U2025 ( .A(\mem<8><5> ), .B(n93), .Y(n2140) );
  OAI21X1 U2026 ( .A(n1896), .B(n15), .C(n2140), .Y(n2361) );
  NAND2X1 U2027 ( .A(\mem<8><6> ), .B(n93), .Y(n2141) );
  OAI21X1 U2028 ( .A(n1896), .B(n1931), .C(n2141), .Y(n2360) );
  NAND2X1 U2029 ( .A(\mem<8><7> ), .B(n93), .Y(n2142) );
  OAI21X1 U2030 ( .A(n1896), .B(n5), .C(n2142), .Y(n2359) );
  OAI21X1 U2031 ( .A(n1896), .B(n11), .C(n363), .Y(n2358) );
  OAI21X1 U2032 ( .A(n1896), .B(n1939), .C(n365), .Y(n2357) );
  OAI21X1 U2033 ( .A(n1896), .B(n1942), .C(n367), .Y(n2356) );
  OAI21X1 U2034 ( .A(n1896), .B(n1943), .C(n369), .Y(n2355) );
  OAI21X1 U2035 ( .A(n1896), .B(n1945), .C(n371), .Y(n2354) );
  OAI21X1 U2036 ( .A(n1896), .B(n1947), .C(n373), .Y(n2353) );
  OAI21X1 U2037 ( .A(n1896), .B(n1949), .C(n375), .Y(n2352) );
  OAI21X1 U2038 ( .A(n1896), .B(n1952), .C(n377), .Y(n2351) );
  NAND3X1 U2039 ( .A(n1961), .B(n2735), .C(n1963), .Y(n2143) );
  NAND2X1 U2040 ( .A(\mem<7><0> ), .B(n95), .Y(n2144) );
  OAI21X1 U2041 ( .A(n1897), .B(n1917), .C(n2144), .Y(n2350) );
  NAND2X1 U2042 ( .A(\mem<7><1> ), .B(n95), .Y(n2145) );
  OAI21X1 U2043 ( .A(n1897), .B(n1918), .C(n2145), .Y(n2349) );
  NAND2X1 U2044 ( .A(\mem<7><2> ), .B(n95), .Y(n2146) );
  OAI21X1 U2045 ( .A(n1897), .B(n1921), .C(n2146), .Y(n2348) );
  NAND2X1 U2046 ( .A(\mem<7><3> ), .B(n95), .Y(n2147) );
  OAI21X1 U2047 ( .A(n1897), .B(n1923), .C(n2147), .Y(n2347) );
  NAND2X1 U2048 ( .A(\mem<7><4> ), .B(n95), .Y(n2148) );
  OAI21X1 U2049 ( .A(n1897), .B(n1925), .C(n2148), .Y(n2346) );
  NAND2X1 U2050 ( .A(\mem<7><5> ), .B(n95), .Y(n2149) );
  OAI21X1 U2051 ( .A(n1897), .B(n1928), .C(n2149), .Y(n2345) );
  NAND2X1 U2052 ( .A(\mem<7><6> ), .B(n95), .Y(n2150) );
  OAI21X1 U2053 ( .A(n1897), .B(n1931), .C(n2150), .Y(n2344) );
  NAND2X1 U2054 ( .A(\mem<7><7> ), .B(n95), .Y(n2151) );
  OAI21X1 U2055 ( .A(n1897), .B(n17), .C(n2151), .Y(n2343) );
  OAI21X1 U2056 ( .A(n1898), .B(n1937), .C(n379), .Y(n2342) );
  OAI21X1 U2057 ( .A(n1898), .B(n1939), .C(n381), .Y(n2341) );
  OAI21X1 U2058 ( .A(n1898), .B(n1941), .C(n383), .Y(n2340) );
  OAI21X1 U2059 ( .A(n1898), .B(n1944), .C(n385), .Y(n2339) );
  OAI21X1 U2060 ( .A(n1898), .B(n1946), .C(n387), .Y(n2338) );
  OAI21X1 U2061 ( .A(n1898), .B(n1947), .C(n389), .Y(n2337) );
  OAI21X1 U2062 ( .A(n1898), .B(n1950), .C(n391), .Y(n2336) );
  OAI21X1 U2063 ( .A(n1898), .B(n1952), .C(n393), .Y(n2335) );
  NAND2X1 U2064 ( .A(\mem<6><0> ), .B(n97), .Y(n2152) );
  OAI21X1 U2065 ( .A(n1899), .B(n1917), .C(n2152), .Y(n2334) );
  NAND2X1 U2066 ( .A(\mem<6><1> ), .B(n97), .Y(n2153) );
  OAI21X1 U2067 ( .A(n1899), .B(n1919), .C(n2153), .Y(n2333) );
  NAND2X1 U2068 ( .A(\mem<6><2> ), .B(n97), .Y(n2154) );
  OAI21X1 U2069 ( .A(n1899), .B(n1921), .C(n2154), .Y(n2332) );
  NAND2X1 U2070 ( .A(\mem<6><3> ), .B(n97), .Y(n2155) );
  OAI21X1 U2071 ( .A(n1899), .B(n1923), .C(n2155), .Y(n2331) );
  NAND2X1 U2072 ( .A(\mem<6><4> ), .B(n97), .Y(n2156) );
  OAI21X1 U2073 ( .A(n1899), .B(n1926), .C(n2156), .Y(n2330) );
  NAND2X1 U2074 ( .A(\mem<6><5> ), .B(n97), .Y(n2157) );
  OAI21X1 U2075 ( .A(n1899), .B(n1929), .C(n2157), .Y(n2329) );
  NAND2X1 U2076 ( .A(\mem<6><6> ), .B(n97), .Y(n2158) );
  OAI21X1 U2077 ( .A(n1899), .B(n1931), .C(n2158), .Y(n2328) );
  NAND2X1 U2078 ( .A(\mem<6><7> ), .B(n97), .Y(n2159) );
  OAI21X1 U2079 ( .A(n1899), .B(n1934), .C(n2159), .Y(n2327) );
  OAI21X1 U2080 ( .A(n1900), .B(n1937), .C(n395), .Y(n2326) );
  OAI21X1 U2081 ( .A(n1900), .B(n1939), .C(n397), .Y(n2325) );
  OAI21X1 U2082 ( .A(n1900), .B(n1942), .C(n399), .Y(n2324) );
  OAI21X1 U2083 ( .A(n1900), .B(n1944), .C(n401), .Y(n2323) );
  OAI21X1 U2084 ( .A(n1900), .B(n1946), .C(n403), .Y(n2322) );
  OAI21X1 U2085 ( .A(n1900), .B(n1947), .C(n405), .Y(n2321) );
  OAI21X1 U2086 ( .A(n1900), .B(n1950), .C(n407), .Y(n2320) );
  OAI21X1 U2087 ( .A(n1900), .B(n1951), .C(n409), .Y(n2319) );
  NAND2X1 U2088 ( .A(\mem<5><0> ), .B(n99), .Y(n2161) );
  OAI21X1 U2089 ( .A(n1901), .B(n1917), .C(n2161), .Y(n2318) );
  NAND2X1 U2090 ( .A(\mem<5><1> ), .B(n99), .Y(n2162) );
  OAI21X1 U2091 ( .A(n1901), .B(n1918), .C(n2162), .Y(n2317) );
  NAND2X1 U2092 ( .A(\mem<5><2> ), .B(n99), .Y(n2163) );
  OAI21X1 U2093 ( .A(n1901), .B(n1921), .C(n2163), .Y(n2316) );
  NAND2X1 U2094 ( .A(\mem<5><3> ), .B(n99), .Y(n2164) );
  OAI21X1 U2095 ( .A(n1901), .B(n1923), .C(n2164), .Y(n2315) );
  NAND2X1 U2096 ( .A(\mem<5><4> ), .B(n99), .Y(n2165) );
  OAI21X1 U2097 ( .A(n1901), .B(n1925), .C(n2165), .Y(n2314) );
  NAND2X1 U2098 ( .A(\mem<5><5> ), .B(n99), .Y(n2166) );
  OAI21X1 U2099 ( .A(n1901), .B(n1928), .C(n2166), .Y(n2313) );
  NAND2X1 U2100 ( .A(\mem<5><6> ), .B(n99), .Y(n2167) );
  OAI21X1 U2101 ( .A(n1901), .B(n1931), .C(n2167), .Y(n2312) );
  NAND2X1 U2102 ( .A(\mem<5><7> ), .B(n99), .Y(n2168) );
  OAI21X1 U2103 ( .A(n1901), .B(n17), .C(n2168), .Y(n2311) );
  OAI21X1 U2104 ( .A(n1902), .B(n1937), .C(n411), .Y(n2310) );
  OAI21X1 U2105 ( .A(n1902), .B(n1939), .C(n413), .Y(n2309) );
  OAI21X1 U2106 ( .A(n1902), .B(n1942), .C(n415), .Y(n2308) );
  OAI21X1 U2107 ( .A(n1902), .B(n1944), .C(n417), .Y(n2307) );
  OAI21X1 U2108 ( .A(n1902), .B(n1946), .C(n419), .Y(n2306) );
  OAI21X1 U2109 ( .A(n1902), .B(n1947), .C(n421), .Y(n2305) );
  OAI21X1 U2110 ( .A(n1902), .B(n1950), .C(n423), .Y(n2304) );
  OAI21X1 U2111 ( .A(n1902), .B(n1952), .C(n425), .Y(n2303) );
  NAND2X1 U2112 ( .A(\mem<4><0> ), .B(n101), .Y(n2170) );
  OAI21X1 U2113 ( .A(n1903), .B(n1916), .C(n2170), .Y(n2302) );
  NAND2X1 U2114 ( .A(\mem<4><1> ), .B(n101), .Y(n2171) );
  OAI21X1 U2115 ( .A(n1903), .B(n13), .C(n2171), .Y(n2301) );
  NAND2X1 U2116 ( .A(\mem<4><2> ), .B(n101), .Y(n2172) );
  OAI21X1 U2117 ( .A(n1903), .B(n1921), .C(n2172), .Y(n2300) );
  NAND2X1 U2118 ( .A(\mem<4><3> ), .B(n101), .Y(n2173) );
  OAI21X1 U2119 ( .A(n1903), .B(n1923), .C(n2173), .Y(n2299) );
  NAND2X1 U2120 ( .A(\mem<4><4> ), .B(n101), .Y(n2174) );
  OAI21X1 U2121 ( .A(n1903), .B(n14), .C(n2174), .Y(n2298) );
  NAND2X1 U2122 ( .A(\mem<4><5> ), .B(n101), .Y(n2175) );
  OAI21X1 U2123 ( .A(n1903), .B(n15), .C(n2175), .Y(n2297) );
  NAND2X1 U2124 ( .A(\mem<4><6> ), .B(n101), .Y(n2176) );
  OAI21X1 U2125 ( .A(n1903), .B(n1931), .C(n2176), .Y(n2296) );
  NAND2X1 U2126 ( .A(\mem<4><7> ), .B(n101), .Y(n2177) );
  OAI21X1 U2127 ( .A(n1903), .B(n1934), .C(n2177), .Y(n2295) );
  OAI21X1 U2128 ( .A(n1904), .B(n1937), .C(n427), .Y(n2294) );
  OAI21X1 U2129 ( .A(n1904), .B(n1939), .C(n429), .Y(n2293) );
  OAI21X1 U2130 ( .A(n1904), .B(n1941), .C(n431), .Y(n2292) );
  OAI21X1 U2131 ( .A(n1904), .B(n1943), .C(n433), .Y(n2291) );
  OAI21X1 U2132 ( .A(n1904), .B(n1945), .C(n435), .Y(n2290) );
  OAI21X1 U2133 ( .A(n1904), .B(n1947), .C(n437), .Y(n2289) );
  OAI21X1 U2134 ( .A(n1904), .B(n1949), .C(n439), .Y(n2288) );
  OAI21X1 U2135 ( .A(n1904), .B(n1951), .C(n441), .Y(n2287) );
  NAND2X1 U2136 ( .A(\mem<3><0> ), .B(n103), .Y(n2179) );
  OAI21X1 U2137 ( .A(n1905), .B(n1917), .C(n2179), .Y(n2286) );
  NAND2X1 U2138 ( .A(\mem<3><1> ), .B(n103), .Y(n2180) );
  OAI21X1 U2139 ( .A(n1905), .B(n13), .C(n2180), .Y(n2285) );
  NAND2X1 U2140 ( .A(\mem<3><2> ), .B(n103), .Y(n2181) );
  OAI21X1 U2141 ( .A(n1905), .B(n1921), .C(n2181), .Y(n2284) );
  NAND2X1 U2142 ( .A(\mem<3><3> ), .B(n103), .Y(n2182) );
  OAI21X1 U2143 ( .A(n1905), .B(n1923), .C(n2182), .Y(n2283) );
  NAND2X1 U2144 ( .A(\mem<3><4> ), .B(n103), .Y(n2183) );
  OAI21X1 U2145 ( .A(n1905), .B(n14), .C(n2183), .Y(n2282) );
  NAND2X1 U2146 ( .A(\mem<3><5> ), .B(n103), .Y(n2184) );
  OAI21X1 U2147 ( .A(n1905), .B(n15), .C(n2184), .Y(n2281) );
  NAND2X1 U2148 ( .A(\mem<3><6> ), .B(n103), .Y(n2185) );
  OAI21X1 U2149 ( .A(n1905), .B(n1931), .C(n2185), .Y(n2280) );
  NAND2X1 U2150 ( .A(\mem<3><7> ), .B(n103), .Y(n2186) );
  OAI21X1 U2151 ( .A(n1905), .B(n17), .C(n2186), .Y(n2279) );
  OAI21X1 U2152 ( .A(n1906), .B(n1937), .C(n443), .Y(n2278) );
  OAI21X1 U2153 ( .A(n1906), .B(n1939), .C(n445), .Y(n2277) );
  OAI21X1 U2154 ( .A(n1906), .B(n1942), .C(n447), .Y(n2276) );
  OAI21X1 U2155 ( .A(n1906), .B(n1944), .C(n449), .Y(n2275) );
  OAI21X1 U2156 ( .A(n1906), .B(n1946), .C(n451), .Y(n2274) );
  OAI21X1 U2157 ( .A(n1906), .B(n1947), .C(n453), .Y(n2273) );
  OAI21X1 U2158 ( .A(n1906), .B(n1950), .C(n455), .Y(n2272) );
  OAI21X1 U2159 ( .A(n1906), .B(n1952), .C(n457), .Y(n2271) );
  NAND2X1 U2160 ( .A(\mem<2><0> ), .B(n105), .Y(n2188) );
  OAI21X1 U2161 ( .A(n1907), .B(n1917), .C(n2188), .Y(n2270) );
  NAND2X1 U2162 ( .A(\mem<2><1> ), .B(n105), .Y(n2189) );
  OAI21X1 U2163 ( .A(n1907), .B(n1918), .C(n2189), .Y(n2269) );
  NAND2X1 U2164 ( .A(\mem<2><2> ), .B(n105), .Y(n2190) );
  OAI21X1 U2165 ( .A(n1907), .B(n1921), .C(n2190), .Y(n2268) );
  NAND2X1 U2166 ( .A(\mem<2><3> ), .B(n105), .Y(n2191) );
  OAI21X1 U2167 ( .A(n1907), .B(n1923), .C(n2191), .Y(n2267) );
  NAND2X1 U2168 ( .A(\mem<2><4> ), .B(n105), .Y(n2192) );
  OAI21X1 U2169 ( .A(n1907), .B(n1925), .C(n2192), .Y(n2266) );
  NAND2X1 U2170 ( .A(\mem<2><5> ), .B(n105), .Y(n2193) );
  OAI21X1 U2171 ( .A(n1907), .B(n1928), .C(n2193), .Y(n2265) );
  NAND2X1 U2172 ( .A(\mem<2><6> ), .B(n105), .Y(n2194) );
  OAI21X1 U2173 ( .A(n1907), .B(n1931), .C(n2194), .Y(n2264) );
  NAND2X1 U2174 ( .A(\mem<2><7> ), .B(n105), .Y(n2195) );
  OAI21X1 U2175 ( .A(n1907), .B(n1934), .C(n2195), .Y(n2263) );
  OAI21X1 U2176 ( .A(n1908), .B(n1936), .C(n459), .Y(n2262) );
  OAI21X1 U2177 ( .A(n1908), .B(n1939), .C(n461), .Y(n2261) );
  OAI21X1 U2178 ( .A(n1908), .B(n1941), .C(n463), .Y(n2260) );
  OAI21X1 U2179 ( .A(n1908), .B(n1944), .C(n465), .Y(n2259) );
  OAI21X1 U2180 ( .A(n1908), .B(n12), .C(n467), .Y(n2258) );
  OAI21X1 U2181 ( .A(n1908), .B(n1947), .C(n469), .Y(n2257) );
  OAI21X1 U2182 ( .A(n1908), .B(n1949), .C(n471), .Y(n2256) );
  OAI21X1 U2183 ( .A(n1908), .B(n1951), .C(n473), .Y(n2255) );
  NAND2X1 U2184 ( .A(\mem<1><0> ), .B(n107), .Y(n2197) );
  OAI21X1 U2185 ( .A(n1909), .B(n1917), .C(n2197), .Y(n2254) );
  NAND2X1 U2186 ( .A(\mem<1><1> ), .B(n107), .Y(n2198) );
  OAI21X1 U2187 ( .A(n1909), .B(n13), .C(n2198), .Y(n2253) );
  NAND2X1 U2188 ( .A(\mem<1><2> ), .B(n107), .Y(n2199) );
  OAI21X1 U2189 ( .A(n1909), .B(n1921), .C(n2199), .Y(n2252) );
  NAND2X1 U2190 ( .A(\mem<1><3> ), .B(n107), .Y(n2200) );
  OAI21X1 U2191 ( .A(n1909), .B(n1923), .C(n2200), .Y(n2251) );
  NAND2X1 U2192 ( .A(\mem<1><4> ), .B(n107), .Y(n2201) );
  OAI21X1 U2193 ( .A(n1909), .B(n14), .C(n2201), .Y(n2250) );
  NAND2X1 U2194 ( .A(\mem<1><5> ), .B(n107), .Y(n2202) );
  OAI21X1 U2195 ( .A(n1909), .B(n15), .C(n2202), .Y(n2249) );
  NAND2X1 U2196 ( .A(\mem<1><6> ), .B(n107), .Y(n2203) );
  OAI21X1 U2197 ( .A(n1909), .B(n1931), .C(n2203), .Y(n2248) );
  NAND2X1 U2198 ( .A(\mem<1><7> ), .B(n107), .Y(n2204) );
  OAI21X1 U2199 ( .A(n1909), .B(n17), .C(n2204), .Y(n2247) );
  OAI21X1 U2200 ( .A(n1910), .B(n6), .C(n475), .Y(n2246) );
  OAI21X1 U2201 ( .A(n1910), .B(n1939), .C(n477), .Y(n2245) );
  OAI21X1 U2202 ( .A(n1910), .B(n1941), .C(n479), .Y(n2244) );
  OAI21X1 U2203 ( .A(n1910), .B(n1944), .C(n481), .Y(n2243) );
  OAI21X1 U2204 ( .A(n1910), .B(n1946), .C(n483), .Y(n2242) );
  OAI21X1 U2205 ( .A(n1910), .B(n1947), .C(n485), .Y(n2241) );
  OAI21X1 U2206 ( .A(n1910), .B(n1950), .C(n487), .Y(n2240) );
  OAI21X1 U2207 ( .A(n1910), .B(n1952), .C(n489), .Y(n2239) );
  NAND2X1 U2208 ( .A(\mem<0><0> ), .B(n109), .Y(n2207) );
  OAI21X1 U2209 ( .A(n1911), .B(n1916), .C(n2207), .Y(n2238) );
  NAND2X1 U2210 ( .A(\mem<0><1> ), .B(n109), .Y(n2208) );
  OAI21X1 U2211 ( .A(n1911), .B(n1919), .C(n2208), .Y(n2237) );
  NAND2X1 U2212 ( .A(\mem<0><2> ), .B(n109), .Y(n2209) );
  OAI21X1 U2213 ( .A(n1911), .B(n1921), .C(n2209), .Y(n2236) );
  NAND2X1 U2214 ( .A(\mem<0><3> ), .B(n109), .Y(n2210) );
  OAI21X1 U2215 ( .A(n1911), .B(n1923), .C(n2210), .Y(n2235) );
  NAND2X1 U2216 ( .A(\mem<0><4> ), .B(n109), .Y(n2211) );
  OAI21X1 U2217 ( .A(n1911), .B(n1926), .C(n2211), .Y(n2234) );
  NAND2X1 U2218 ( .A(\mem<0><5> ), .B(n109), .Y(n2212) );
  OAI21X1 U2219 ( .A(n1911), .B(n1929), .C(n2212), .Y(n2233) );
  NAND2X1 U2220 ( .A(\mem<0><6> ), .B(n109), .Y(n2213) );
  OAI21X1 U2221 ( .A(n1911), .B(n1931), .C(n2213), .Y(n2232) );
  NAND2X1 U2222 ( .A(\mem<0><7> ), .B(n109), .Y(n2214) );
  OAI21X1 U2223 ( .A(n1911), .B(n1933), .C(n2214), .Y(n2231) );
  NAND2X1 U2224 ( .A(\mem<0><8> ), .B(n109), .Y(n2215) );
  OAI21X1 U2225 ( .A(n1911), .B(n1936), .C(n2215), .Y(n2230) );
  NAND2X1 U2226 ( .A(\mem<0><9> ), .B(n109), .Y(n2216) );
  OAI21X1 U2227 ( .A(n1911), .B(n1939), .C(n2216), .Y(n2229) );
  NAND2X1 U2228 ( .A(\mem<0><10> ), .B(n109), .Y(n2217) );
  OAI21X1 U2229 ( .A(n1911), .B(n1941), .C(n2217), .Y(n2228) );
  NAND2X1 U2230 ( .A(\mem<0><11> ), .B(n109), .Y(n2218) );
  OAI21X1 U2231 ( .A(n1911), .B(n1943), .C(n2218), .Y(n2227) );
  NAND2X1 U2232 ( .A(\mem<0><12> ), .B(n109), .Y(n2219) );
  OAI21X1 U2233 ( .A(n1911), .B(n1945), .C(n2219), .Y(n2226) );
  NAND2X1 U2234 ( .A(\mem<0><13> ), .B(n109), .Y(n2220) );
  OAI21X1 U2235 ( .A(n1911), .B(n1947), .C(n2220), .Y(n2225) );
  NAND2X1 U2236 ( .A(\mem<0><14> ), .B(n109), .Y(n2221) );
  OAI21X1 U2237 ( .A(n1911), .B(n1949), .C(n2221), .Y(n2224) );
  NAND2X1 U2238 ( .A(\mem<0><15> ), .B(n109), .Y(n2222) );
  OAI21X1 U2239 ( .A(n1911), .B(n1951), .C(n2222), .Y(n2223) );
endmodule


module memc_Size5_1 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , n56, n57, n65, n73, n81, n89, n97, n105,
         n113, n114, n115, n172, n229, n286, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, net85891, net85954, net86080, net89225, net89223, net89361,
         net89359, net89515, net89513, net89511, net89783, net89781, net89779,
         net89777, net89775, net90255, net90251, net90249, net90247, net90245,
         net90243, net90241, net90239, net90935, net96102, net102546,
         net102545, net102667, net102825, net102831, net102837, net102839,
         net102846, net103275, net117952, net117994, net121110, net121136,
         net121144, net121143, net121526, net121576, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n58, n59, n60, n61, n62, n63, n64,
         n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80,
         n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95, n96,
         n98, n99, n100, n101, n102, n103, n104, n106, n107, n108, n109, n110,
         n111, n112, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n287, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n447), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n446), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n445), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n444), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n443), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n442), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n441), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n440), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n439), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n438), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n437), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n436), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n435), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n434), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n433), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n432), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n431), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n430), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n429), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n428), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n427), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n426), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n425), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n424), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n423), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n422), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n421), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n420), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n419), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n418), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n417), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n416), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n415), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n414), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n413), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n412), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n411), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n410), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n409), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n408), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n407), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n406), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n405), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n404), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n403), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n402), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n401), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n400), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n399), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n398), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n397), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n396), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n395), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n394), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n393), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n392), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n391), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n390), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n389), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n388), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n387), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n386), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n385), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n384), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n383), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n382), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n381), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n380), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n379), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n378), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n377), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n376), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n375), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n374), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n373), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n372), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n371), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n370), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n369), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n368), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n367), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n366), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n365), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n364), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n363), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n362), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n361), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n360), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n359), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n358), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n357), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n356), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n355), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n354), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n353), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n352), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n351), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n350), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n349), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n348), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n347), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n346), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n345), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n344), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n343), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n342), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n341), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n340), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n339), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n338), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n337), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n336), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n335), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n334), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n333), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n332), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n331), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n330), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n329), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n328), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n327), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n326), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n325), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n324), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n323), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n322), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n321), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n320), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n319), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n318), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n317), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n316), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n315), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n314), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n313), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n312), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n311), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n310), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n309), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n308), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n307), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n306), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n305), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n304), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n303), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n302), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n301), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n300), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n299), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n298), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n297), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n296), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n294), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n292), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n291), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n290), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n289), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n288), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(net121576), .B(net90935), .Y(n56) );
  OAI21X1 U50 ( .A(n648), .B(n723), .C(n567), .Y(n288) );
  OAI21X1 U52 ( .A(n648), .B(n722), .C(n565), .Y(n289) );
  OAI21X1 U54 ( .A(n648), .B(n721), .C(n563), .Y(n290) );
  OAI21X1 U56 ( .A(n648), .B(n720), .C(n561), .Y(n291) );
  OAI21X1 U58 ( .A(n648), .B(n719), .C(n559), .Y(n292) );
  OAI21X1 U62 ( .A(n723), .B(n711), .C(n557), .Y(n293) );
  OAI21X1 U64 ( .A(n722), .B(n711), .C(n555), .Y(n294) );
  OAI21X1 U66 ( .A(n721), .B(n711), .C(n553), .Y(n295) );
  OAI21X1 U68 ( .A(n720), .B(n711), .C(n551), .Y(n296) );
  OAI21X1 U70 ( .A(n719), .B(n711), .C(n549), .Y(n297) );
  OAI21X1 U74 ( .A(n723), .B(n709), .C(n547), .Y(n298) );
  OAI21X1 U76 ( .A(n722), .B(n709), .C(n545), .Y(n299) );
  OAI21X1 U78 ( .A(n721), .B(n709), .C(n543), .Y(n300) );
  OAI21X1 U80 ( .A(n720), .B(n709), .C(n541), .Y(n301) );
  OAI21X1 U82 ( .A(n719), .B(n709), .C(n539), .Y(n302) );
  OAI21X1 U86 ( .A(n723), .B(n707), .C(n537), .Y(n303) );
  OAI21X1 U88 ( .A(n722), .B(n707), .C(n535), .Y(n304) );
  OAI21X1 U90 ( .A(n721), .B(n707), .C(n533), .Y(n305) );
  OAI21X1 U92 ( .A(n720), .B(n707), .C(n531), .Y(n306) );
  OAI21X1 U94 ( .A(n719), .B(n707), .C(n529), .Y(n307) );
  OAI21X1 U98 ( .A(n723), .B(n705), .C(n527), .Y(n308) );
  OAI21X1 U100 ( .A(n722), .B(n705), .C(n525), .Y(n309) );
  OAI21X1 U102 ( .A(n721), .B(n705), .C(n523), .Y(n310) );
  OAI21X1 U104 ( .A(n720), .B(n705), .C(n521), .Y(n311) );
  OAI21X1 U106 ( .A(n719), .B(n705), .C(n519), .Y(n312) );
  OAI21X1 U110 ( .A(n723), .B(n703), .C(n517), .Y(n313) );
  OAI21X1 U112 ( .A(n722), .B(n703), .C(n515), .Y(n314) );
  OAI21X1 U114 ( .A(n721), .B(n703), .C(n513), .Y(n315) );
  OAI21X1 U116 ( .A(n720), .B(n703), .C(n511), .Y(n316) );
  OAI21X1 U118 ( .A(n719), .B(n703), .C(n509), .Y(n317) );
  OAI21X1 U122 ( .A(n723), .B(n701), .C(n507), .Y(n318) );
  OAI21X1 U124 ( .A(n722), .B(n701), .C(n505), .Y(n319) );
  OAI21X1 U126 ( .A(n721), .B(n701), .C(n503), .Y(n320) );
  OAI21X1 U128 ( .A(n720), .B(n701), .C(n501), .Y(n321) );
  OAI21X1 U130 ( .A(n719), .B(n701), .C(n499), .Y(n322) );
  OAI21X1 U134 ( .A(n723), .B(n699), .C(n497), .Y(n323) );
  OAI21X1 U136 ( .A(n722), .B(n699), .C(n495), .Y(n324) );
  OAI21X1 U138 ( .A(n721), .B(n699), .C(n493), .Y(n325) );
  OAI21X1 U140 ( .A(n720), .B(n699), .C(n491), .Y(n326) );
  OAI21X1 U142 ( .A(n719), .B(n699), .C(n489), .Y(n327) );
  NAND3X1 U146 ( .A(net89359), .B(n115), .C(net89223), .Y(n114) );
  OAI21X1 U147 ( .A(n723), .B(n696), .C(n487), .Y(n328) );
  OAI21X1 U149 ( .A(n722), .B(n696), .C(n485), .Y(n329) );
  OAI21X1 U151 ( .A(n721), .B(n696), .C(n483), .Y(n330) );
  OAI21X1 U153 ( .A(n720), .B(n696), .C(n481), .Y(n331) );
  OAI21X1 U155 ( .A(n719), .B(n696), .C(n479), .Y(n332) );
  OAI21X1 U159 ( .A(n723), .B(n694), .C(n477), .Y(n333) );
  OAI21X1 U161 ( .A(n722), .B(n694), .C(n475), .Y(n334) );
  OAI21X1 U163 ( .A(n721), .B(n694), .C(n473), .Y(n335) );
  OAI21X1 U165 ( .A(n720), .B(n694), .C(n471), .Y(n336) );
  OAI21X1 U167 ( .A(n719), .B(n694), .C(n469), .Y(n337) );
  OAI21X1 U171 ( .A(n723), .B(n693), .C(n467), .Y(n338) );
  OAI21X1 U173 ( .A(n722), .B(n693), .C(n465), .Y(n339) );
  OAI21X1 U175 ( .A(n721), .B(n693), .C(n463), .Y(n340) );
  OAI21X1 U177 ( .A(n720), .B(n693), .C(n461), .Y(n341) );
  OAI21X1 U179 ( .A(n719), .B(n693), .C(n459), .Y(n342) );
  OAI21X1 U183 ( .A(n723), .B(n691), .C(n457), .Y(n343) );
  OAI21X1 U185 ( .A(n722), .B(n691), .C(n455), .Y(n344) );
  OAI21X1 U187 ( .A(n721), .B(n691), .C(n453), .Y(n345) );
  OAI21X1 U189 ( .A(n720), .B(n691), .C(n451), .Y(n346) );
  OAI21X1 U191 ( .A(n719), .B(n691), .C(n449), .Y(n347) );
  OAI21X1 U195 ( .A(n723), .B(n689), .C(n287), .Y(n348) );
  OAI21X1 U197 ( .A(n722), .B(n689), .C(n284), .Y(n349) );
  OAI21X1 U199 ( .A(n721), .B(n689), .C(n282), .Y(n350) );
  OAI21X1 U201 ( .A(n720), .B(n689), .C(n280), .Y(n351) );
  OAI21X1 U203 ( .A(n719), .B(n689), .C(n278), .Y(n352) );
  OAI21X1 U207 ( .A(n723), .B(n687), .C(n276), .Y(n353) );
  OAI21X1 U209 ( .A(n722), .B(n687), .C(n274), .Y(n354) );
  OAI21X1 U211 ( .A(n721), .B(n687), .C(n272), .Y(n355) );
  OAI21X1 U213 ( .A(n720), .B(n687), .C(n270), .Y(n356) );
  OAI21X1 U215 ( .A(n719), .B(n687), .C(n268), .Y(n357) );
  OAI21X1 U219 ( .A(n723), .B(n684), .C(n266), .Y(n358) );
  OAI21X1 U221 ( .A(n722), .B(n684), .C(n264), .Y(n359) );
  OAI21X1 U223 ( .A(n721), .B(n684), .C(n262), .Y(n360) );
  OAI21X1 U225 ( .A(n720), .B(n684), .C(n260), .Y(n361) );
  OAI21X1 U227 ( .A(n719), .B(n684), .C(n258), .Y(n362) );
  OAI21X1 U231 ( .A(n723), .B(n682), .C(n256), .Y(n363) );
  OAI21X1 U233 ( .A(n722), .B(n682), .C(n254), .Y(n364) );
  OAI21X1 U235 ( .A(n721), .B(n682), .C(n252), .Y(n365) );
  OAI21X1 U237 ( .A(n720), .B(n682), .C(n250), .Y(n366) );
  OAI21X1 U239 ( .A(n719), .B(n682), .C(n248), .Y(n367) );
  NAND3X1 U243 ( .A(n115), .B(net89361), .C(net89223), .Y(n172) );
  OAI21X1 U244 ( .A(n723), .B(n681), .C(n246), .Y(n368) );
  OAI21X1 U246 ( .A(n722), .B(n681), .C(n244), .Y(n369) );
  OAI21X1 U248 ( .A(n721), .B(n681), .C(n242), .Y(n370) );
  OAI21X1 U250 ( .A(n720), .B(n681), .C(n240), .Y(n371) );
  OAI21X1 U252 ( .A(n719), .B(n681), .C(n238), .Y(n372) );
  OAI21X1 U256 ( .A(n723), .B(n679), .C(n236), .Y(n373) );
  OAI21X1 U258 ( .A(n722), .B(n679), .C(n234), .Y(n374) );
  OAI21X1 U260 ( .A(n721), .B(n679), .C(n232), .Y(n375) );
  OAI21X1 U262 ( .A(n720), .B(n679), .C(n230), .Y(n376) );
  OAI21X1 U264 ( .A(n719), .B(n679), .C(n227), .Y(n377) );
  OAI21X1 U268 ( .A(n723), .B(n676), .C(n225), .Y(n378) );
  OAI21X1 U270 ( .A(n722), .B(n676), .C(n223), .Y(n379) );
  OAI21X1 U272 ( .A(n721), .B(n676), .C(n221), .Y(n380) );
  OAI21X1 U274 ( .A(n720), .B(n676), .C(n219), .Y(n381) );
  OAI21X1 U276 ( .A(n719), .B(n676), .C(n217), .Y(n382) );
  OAI21X1 U280 ( .A(n723), .B(n675), .C(n215), .Y(n383) );
  OAI21X1 U282 ( .A(n722), .B(n675), .C(n213), .Y(n384) );
  OAI21X1 U284 ( .A(n721), .B(n675), .C(n211), .Y(n385) );
  OAI21X1 U286 ( .A(n720), .B(n675), .C(n209), .Y(n386) );
  OAI21X1 U288 ( .A(n719), .B(n675), .C(n207), .Y(n387) );
  OAI21X1 U292 ( .A(n723), .B(n672), .C(n205), .Y(n388) );
  OAI21X1 U294 ( .A(n722), .B(n672), .C(n203), .Y(n389) );
  OAI21X1 U296 ( .A(n721), .B(n672), .C(n201), .Y(n390) );
  OAI21X1 U298 ( .A(n720), .B(n672), .C(n199), .Y(n391) );
  OAI21X1 U300 ( .A(n719), .B(n672), .C(n197), .Y(n392) );
  OAI21X1 U304 ( .A(n723), .B(n671), .C(n195), .Y(n393) );
  OAI21X1 U306 ( .A(n722), .B(n671), .C(n193), .Y(n394) );
  OAI21X1 U308 ( .A(n721), .B(n671), .C(n191), .Y(n395) );
  OAI21X1 U310 ( .A(n720), .B(n671), .C(n189), .Y(n396) );
  OAI21X1 U312 ( .A(n719), .B(n671), .C(n187), .Y(n397) );
  OAI21X1 U316 ( .A(n723), .B(n669), .C(n185), .Y(n398) );
  OAI21X1 U318 ( .A(n722), .B(n669), .C(n183), .Y(n399) );
  OAI21X1 U320 ( .A(n721), .B(n669), .C(n181), .Y(n400) );
  OAI21X1 U322 ( .A(n720), .B(n669), .C(n179), .Y(n401) );
  OAI21X1 U324 ( .A(n719), .B(n669), .C(n177), .Y(n402) );
  OAI21X1 U328 ( .A(n723), .B(n667), .C(n175), .Y(n403) );
  OAI21X1 U330 ( .A(n722), .B(n667), .C(n173), .Y(n404) );
  OAI21X1 U332 ( .A(n721), .B(n667), .C(n170), .Y(n405) );
  OAI21X1 U334 ( .A(n720), .B(n667), .C(n168), .Y(n406) );
  OAI21X1 U336 ( .A(n719), .B(n667), .C(n166), .Y(n407) );
  NAND3X1 U340 ( .A(n115), .B(net89225), .C(net89359), .Y(n229) );
  OAI21X1 U341 ( .A(n723), .B(n665), .C(n164), .Y(n408) );
  OAI21X1 U343 ( .A(n722), .B(n665), .C(n162), .Y(n409) );
  OAI21X1 U345 ( .A(n721), .B(n665), .C(n160), .Y(n410) );
  OAI21X1 U347 ( .A(n720), .B(n665), .C(n158), .Y(n411) );
  OAI21X1 U349 ( .A(n719), .B(n665), .C(n156), .Y(n412) );
  NOR3X1 U353 ( .A(net89783), .B(net102546), .C(net89515), .Y(n57) );
  OAI21X1 U354 ( .A(n723), .B(n663), .C(n154), .Y(n413) );
  OAI21X1 U356 ( .A(n722), .B(n663), .C(n152), .Y(n414) );
  OAI21X1 U358 ( .A(n721), .B(n663), .C(n150), .Y(n415) );
  OAI21X1 U360 ( .A(n720), .B(n663), .C(n148), .Y(n416) );
  OAI21X1 U362 ( .A(n719), .B(n663), .C(n146), .Y(n417) );
  NOR3X1 U366 ( .A(net89783), .B(net103275), .C(net89515), .Y(n65) );
  OAI21X1 U367 ( .A(n723), .B(n661), .C(n144), .Y(n418) );
  OAI21X1 U369 ( .A(n722), .B(n661), .C(n142), .Y(n419) );
  OAI21X1 U371 ( .A(n721), .B(n661), .C(n140), .Y(n420) );
  OAI21X1 U373 ( .A(n720), .B(n661), .C(n138), .Y(n421) );
  OAI21X1 U375 ( .A(n719), .B(n661), .C(n136), .Y(n422) );
  NOR3X1 U379 ( .A(net102831), .B(net89781), .C(net89515), .Y(n73) );
  OAI21X1 U380 ( .A(n723), .B(n659), .C(n134), .Y(n423) );
  OAI21X1 U382 ( .A(n722), .B(n659), .C(n132), .Y(n424) );
  OAI21X1 U384 ( .A(n721), .B(n659), .C(n130), .Y(n425) );
  OAI21X1 U386 ( .A(n720), .B(n659), .C(n128), .Y(n426) );
  OAI21X1 U388 ( .A(n719), .B(n659), .C(n126), .Y(n427) );
  NOR3X1 U392 ( .A(net103275), .B(net89775), .C(net89515), .Y(n81) );
  OAI21X1 U393 ( .A(n723), .B(n657), .C(n124), .Y(n428) );
  OAI21X1 U395 ( .A(n722), .B(n657), .C(n122), .Y(n429) );
  OAI21X1 U397 ( .A(n721), .B(n657), .C(n120), .Y(n430) );
  OAI21X1 U399 ( .A(n720), .B(n657), .C(n118), .Y(n431) );
  OAI21X1 U401 ( .A(n719), .B(n657), .C(n116), .Y(n432) );
  NOR3X1 U405 ( .A(net102831), .B(net89513), .C(net89783), .Y(n89) );
  OAI21X1 U406 ( .A(n723), .B(n655), .C(n111), .Y(n433) );
  OAI21X1 U408 ( .A(n722), .B(n655), .C(n109), .Y(n434) );
  OAI21X1 U410 ( .A(n721), .B(n655), .C(n107), .Y(n435) );
  OAI21X1 U412 ( .A(n720), .B(n655), .C(n104), .Y(n436) );
  OAI21X1 U414 ( .A(n719), .B(n655), .C(n102), .Y(n437) );
  NOR3X1 U418 ( .A(net102825), .B(net89513), .C(net89783), .Y(n97) );
  OAI21X1 U419 ( .A(n723), .B(n653), .C(n100), .Y(n438) );
  OAI21X1 U421 ( .A(n722), .B(n653), .C(n98), .Y(n439) );
  OAI21X1 U423 ( .A(n721), .B(n653), .C(n95), .Y(n440) );
  OAI21X1 U425 ( .A(n720), .B(n653), .C(n93), .Y(n441) );
  OAI21X1 U427 ( .A(n719), .B(n653), .C(n91), .Y(n442) );
  NOR3X1 U431 ( .A(net89777), .B(net89513), .C(net102831), .Y(n105) );
  OAI21X1 U432 ( .A(n723), .B(n651), .C(n88), .Y(n443) );
  OAI21X1 U435 ( .A(n722), .B(n651), .C(n86), .Y(n444) );
  OAI21X1 U438 ( .A(n721), .B(n651), .C(n84), .Y(n445) );
  OAI21X1 U441 ( .A(n720), .B(n651), .C(n82), .Y(n446) );
  OAI21X1 U444 ( .A(n719), .B(n651), .C(n79), .Y(n447) );
  NOR3X1 U448 ( .A(net89775), .B(net89513), .C(net103275), .Y(n113) );
  NAND3X1 U449 ( .A(net89361), .B(net89225), .C(n115), .Y(n286) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n115) );
  INVX2 U3 ( .A(n583), .Y(n723) );
  INVX2 U4 ( .A(n582), .Y(n722) );
  INVX2 U5 ( .A(n581), .Y(n721) );
  INVX2 U6 ( .A(n580), .Y(n720) );
  INVX2 U7 ( .A(n579), .Y(n719) );
  INVX1 U8 ( .A(\mem<9><2> ), .Y(n860) );
  INVX1 U9 ( .A(\mem<8><2> ), .Y(n861) );
  INVX1 U10 ( .A(\mem<11><2> ), .Y(n862) );
  INVX1 U11 ( .A(\mem<8><1> ), .Y(n800) );
  INVX1 U12 ( .A(\mem<5><1> ), .Y(n791) );
  INVX1 U13 ( .A(\mem<4><1> ), .Y(n792) );
  INVX1 U14 ( .A(\mem<7><1> ), .Y(n793) );
  INVX1 U15 ( .A(\mem<15><2> ), .Y(n868) );
  INVX1 U16 ( .A(\mem<14><2> ), .Y(n869) );
  INVX1 U17 ( .A(\mem<13><2> ), .Y(n866) );
  INVX1 U18 ( .A(\mem<12><2> ), .Y(n867) );
  INVX1 U19 ( .A(\mem<10><2> ), .Y(n863) );
  INVX1 U20 ( .A(\mem<7><2> ), .Y(n854) );
  INVX1 U21 ( .A(\mem<6><2> ), .Y(n855) );
  INVX1 U22 ( .A(\mem<0><2> ), .Y(n847) );
  INVX1 U23 ( .A(\mem<1><2> ), .Y(n846) );
  INVX1 U24 ( .A(\mem<2><2> ), .Y(n849) );
  INVX1 U25 ( .A(\mem<3><2> ), .Y(n848) );
  INVX1 U26 ( .A(\mem<4><2> ), .Y(n853) );
  INVX1 U27 ( .A(\mem<5><2> ), .Y(n852) );
  INVX1 U28 ( .A(\mem<21><2> ), .Y(n880) );
  INVX1 U29 ( .A(\mem<20><2> ), .Y(n881) );
  INVX1 U30 ( .A(\mem<16><2> ), .Y(n876) );
  INVX1 U31 ( .A(\mem<17><2> ), .Y(n875) );
  INVX1 U32 ( .A(\mem<22><2> ), .Y(n883) );
  INVX1 U33 ( .A(\mem<23><2> ), .Y(n882) );
  INVX1 U34 ( .A(\mem<29><2> ), .Y(n894) );
  INVX1 U35 ( .A(\mem<28><2> ), .Y(n895) );
  INVX1 U36 ( .A(\mem<24><2> ), .Y(n889) );
  INVX1 U37 ( .A(\mem<25><2> ), .Y(n888) );
  INVX1 U38 ( .A(\mem<26><2> ), .Y(n891) );
  INVX1 U39 ( .A(\mem<27><2> ), .Y(n890) );
  INVX1 U40 ( .A(\mem<30><2> ), .Y(n897) );
  INVX1 U41 ( .A(\mem<31><2> ), .Y(n896) );
  INVX1 U42 ( .A(\mem<15><1> ), .Y(n806) );
  INVX1 U43 ( .A(\mem<14><1> ), .Y(n807) );
  INVX1 U44 ( .A(\mem<12><3> ), .Y(n925) );
  INVX1 U45 ( .A(\mem<13><3> ), .Y(n924) );
  INVX1 U46 ( .A(\mem<9><3> ), .Y(n920) );
  INVX1 U47 ( .A(\mem<8><3> ), .Y(n921) );
  INVX1 U48 ( .A(\mem<15><3> ), .Y(n926) );
  INVX1 U49 ( .A(\mem<14><3> ), .Y(n927) );
  INVX1 U51 ( .A(\mem<3><3> ), .Y(n908) );
  INVX1 U53 ( .A(\mem<2><3> ), .Y(n909) );
  INVX1 U55 ( .A(\mem<4><3> ), .Y(n913) );
  INVX1 U57 ( .A(\mem<5><3> ), .Y(n912) );
  INVX1 U59 ( .A(\mem<7><3> ), .Y(n914) );
  INVX1 U60 ( .A(\mem<6><3> ), .Y(n915) );
  INVX1 U61 ( .A(\mem<0><3> ), .Y(n907) );
  INVX1 U63 ( .A(\mem<1><3> ), .Y(n906) );
  INVX1 U65 ( .A(\mem<17><3> ), .Y(n934) );
  INVX1 U67 ( .A(\mem<16><3> ), .Y(n935) );
  INVX1 U69 ( .A(\mem<22><3> ), .Y(n943) );
  INVX1 U71 ( .A(\mem<23><3> ), .Y(n942) );
  INVX1 U72 ( .A(\mem<20><3> ), .Y(n941) );
  INVX1 U73 ( .A(\mem<21><3> ), .Y(n940) );
  INVX1 U75 ( .A(\mem<18><3> ), .Y(n937) );
  INVX1 U77 ( .A(\mem<19><3> ), .Y(n936) );
  INVX1 U79 ( .A(\mem<31><3> ), .Y(n956) );
  INVX1 U81 ( .A(\mem<30><3> ), .Y(n957) );
  INVX1 U83 ( .A(\mem<27><3> ), .Y(n950) );
  INVX1 U84 ( .A(\mem<26><3> ), .Y(n951) );
  INVX1 U85 ( .A(\mem<24><3> ), .Y(n949) );
  INVX1 U87 ( .A(\mem<25><3> ), .Y(n948) );
  INVX1 U89 ( .A(\mem<28><3> ), .Y(n955) );
  INVX1 U91 ( .A(\mem<29><3> ), .Y(n954) );
  INVX1 U93 ( .A(\mem<13><4> ), .Y(n51) );
  INVX1 U95 ( .A(\mem<12><4> ), .Y(n50) );
  INVX1 U96 ( .A(\mem<7><4> ), .Y(n62) );
  INVX1 U97 ( .A(\mem<6><4> ), .Y(n61) );
  INVX1 U99 ( .A(\mem<2><4> ), .Y(n68) );
  INVX1 U101 ( .A(\mem<3><4> ), .Y(n69) );
  INVX1 U103 ( .A(\mem<1><4> ), .Y(n71) );
  INVX1 U105 ( .A(\mem<0><4> ), .Y(n70) );
  INVX1 U107 ( .A(\mem<4><4> ), .Y(n63) );
  INVX1 U108 ( .A(\mem<5><4> ), .Y(n64) );
  INVX1 U109 ( .A(\mem<31><4> ), .Y(n20) );
  INVX1 U111 ( .A(\mem<30><4> ), .Y(n19) );
  INVX1 U113 ( .A(\mem<27><4> ), .Y(n26) );
  INVX1 U115 ( .A(\mem<26><4> ), .Y(n25) );
  INVX1 U117 ( .A(\mem<24><4> ), .Y(n27) );
  INVX1 U119 ( .A(\mem<25><4> ), .Y(n28) );
  INVX1 U120 ( .A(\mem<28><4> ), .Y(n21) );
  INVX1 U121 ( .A(\mem<29><4> ), .Y(n22) );
  INVX1 U123 ( .A(\mem<23><4> ), .Y(n34) );
  INVX1 U125 ( .A(\mem<22><4> ), .Y(n33) );
  INVX1 U127 ( .A(\mem<16><4> ), .Y(n41) );
  INVX1 U129 ( .A(\mem<17><4> ), .Y(n42) );
  INVX1 U131 ( .A(\mem<18><4> ), .Y(n39) );
  INVX1 U132 ( .A(\mem<19><4> ), .Y(n40) );
  INVX1 U133 ( .A(\mem<20><4> ), .Y(n35) );
  INVX1 U135 ( .A(\mem<21><4> ), .Y(n36) );
  INVX1 U137 ( .A(\mem<13><0> ), .Y(n743) );
  INVX1 U139 ( .A(\mem<12><0> ), .Y(n744) );
  INVX1 U141 ( .A(\mem<8><0> ), .Y(n739) );
  INVX1 U143 ( .A(\mem<9><0> ), .Y(n738) );
  INVX1 U144 ( .A(\mem<14><0> ), .Y(n746) );
  INVX1 U145 ( .A(\mem<15><0> ), .Y(n745) );
  INVX1 U148 ( .A(\mem<0><0> ), .Y(n725) );
  INVX1 U150 ( .A(\mem<1><0> ), .Y(n724) );
  INVX1 U152 ( .A(\mem<4><0> ), .Y(n731) );
  INVX1 U154 ( .A(\mem<5><0> ), .Y(n730) );
  INVX1 U156 ( .A(\mem<6><0> ), .Y(n733) );
  INVX1 U157 ( .A(\mem<7><0> ), .Y(n732) );
  INVX1 U158 ( .A(\mem<2><0> ), .Y(n727) );
  INVX1 U160 ( .A(\mem<3><0> ), .Y(n726) );
  INVX1 U162 ( .A(\mem<29><0> ), .Y(n773) );
  INVX1 U164 ( .A(\mem<28><0> ), .Y(n774) );
  INVX1 U166 ( .A(\mem<27><0> ), .Y(n769) );
  INVX1 U168 ( .A(\mem<26><0> ), .Y(n770) );
  INVX1 U169 ( .A(\mem<25><0> ), .Y(n767) );
  INVX1 U170 ( .A(\mem<24><0> ), .Y(n768) );
  INVX1 U172 ( .A(\mem<31><0> ), .Y(n775) );
  INVX1 U174 ( .A(\mem<30><0> ), .Y(n776) );
  INVX1 U176 ( .A(\mem<21><0> ), .Y(n759) );
  INVX1 U178 ( .A(\mem<20><0> ), .Y(n760) );
  INVX1 U180 ( .A(\mem<17><0> ), .Y(n753) );
  INVX1 U181 ( .A(\mem<16><0> ), .Y(n754) );
  INVX1 U182 ( .A(\mem<18><0> ), .Y(n756) );
  INVX1 U184 ( .A(\mem<19><0> ), .Y(n755) );
  INVX1 U186 ( .A(\mem<22><0> ), .Y(n762) );
  INVX1 U188 ( .A(\mem<23><0> ), .Y(n761) );
  INVX1 U190 ( .A(\mem<23><1> ), .Y(n821) );
  INVX1 U192 ( .A(\mem<22><1> ), .Y(n822) );
  INVX1 U193 ( .A(\mem<16><1> ), .Y(n814) );
  INVX1 U194 ( .A(\mem<17><1> ), .Y(n813) );
  INVX1 U196 ( .A(\mem<18><1> ), .Y(n816) );
  INVX1 U198 ( .A(\mem<19><1> ), .Y(n815) );
  INVX1 U200 ( .A(\mem<20><1> ), .Y(n820) );
  INVX1 U202 ( .A(\mem<21><1> ), .Y(n819) );
  INVX1 U204 ( .A(\mem<31><1> ), .Y(n835) );
  INVX1 U205 ( .A(\mem<30><1> ), .Y(n836) );
  INVX1 U206 ( .A(\mem<26><1> ), .Y(n830) );
  INVX1 U208 ( .A(\mem<27><1> ), .Y(n829) );
  INVX1 U210 ( .A(\mem<24><1> ), .Y(n828) );
  INVX1 U212 ( .A(\mem<25><1> ), .Y(n827) );
  INVX1 U214 ( .A(\mem<28><1> ), .Y(n834) );
  INVX1 U216 ( .A(\mem<29><1> ), .Y(n833) );
  INVX1 U217 ( .A(\mem<2><1> ), .Y(n788) );
  INVX1 U218 ( .A(\mem<3><1> ), .Y(n787) );
  INVX1 U220 ( .A(\mem<0><1> ), .Y(n786) );
  INVX1 U222 ( .A(\mem<1><1> ), .Y(n785) );
  INVX1 U224 ( .A(\mem<9><1> ), .Y(n799) );
  INVX1 U226 ( .A(\mem<6><1> ), .Y(n794) );
  INVX1 U228 ( .A(rst), .Y(net90935) );
  AND2X2 U229 ( .A(n6), .B(n10), .Y(\data_out<4> ) );
  AND2X2 U230 ( .A(n9), .B(net90935), .Y(n6) );
  MUX2X1 U232 ( .B(n11), .A(n12), .S(net89223), .Y(n10) );
  MUX2X1 U234 ( .B(n43), .A(n44), .S(net89359), .Y(n11) );
  MUX2X1 U236 ( .B(n55), .A(n58), .S(net89513), .Y(n43) );
  MUX2X1 U238 ( .B(n67), .A(n66), .S(net89783), .Y(n55) );
  MUX2X1 U240 ( .B(n68), .A(n69), .S(net90241), .Y(n67) );
  INVX8 U241 ( .A(net90255), .Y(net90241) );
  MUX2X1 U242 ( .B(n70), .A(n71), .S(net90249), .Y(n66) );
  INVX8 U245 ( .A(net90251), .Y(net90249) );
  INVX8 U247 ( .A(N11), .Y(net89783) );
  MUX2X1 U249 ( .B(n59), .A(n60), .S(net89779), .Y(n58) );
  MUX2X1 U251 ( .B(n63), .A(n64), .S(net90241), .Y(n59) );
  MUX2X1 U253 ( .B(n61), .A(n62), .S(net90243), .Y(n60) );
  INVX8 U254 ( .A(net90251), .Y(net90243) );
  INVX8 U255 ( .A(net89783), .Y(net89779) );
  INVX8 U257 ( .A(net89515), .Y(net89513) );
  MUX2X1 U259 ( .B(n45), .A(n46), .S(net89513), .Y(n44) );
  MUX2X1 U261 ( .B(n52), .A(n7), .S(net89783), .Y(n45) );
  INVX1 U263 ( .A(n1), .Y(n52) );
  MUX2X1 U265 ( .B(\mem<11><4> ), .A(\mem<10><4> ), .S(net121144), .Y(n1) );
  INVX1 U266 ( .A(net121143), .Y(net121144) );
  AND2X2 U267 ( .A(n2), .B(n3), .Y(n7) );
  NAND2X1 U269 ( .A(n53), .B(net117994), .Y(n2) );
  INVX1 U271 ( .A(\mem<8><4> ), .Y(n53) );
  INVX1 U273 ( .A(net121110), .Y(net117994) );
  NAND2X1 U275 ( .A(n54), .B(net90247), .Y(n3) );
  INVX1 U277 ( .A(\mem<9><4> ), .Y(n54) );
  INVX8 U278 ( .A(net90251), .Y(net90247) );
  MUX2X1 U279 ( .B(n47), .A(n8), .S(net89779), .Y(n46) );
  MUX2X1 U281 ( .B(n50), .A(n51), .S(net90239), .Y(n47) );
  INVX8 U283 ( .A(net90255), .Y(net90239) );
  AND2X2 U285 ( .A(n4), .B(n5), .Y(n8) );
  NAND2X1 U287 ( .A(n48), .B(net102839), .Y(n4) );
  INVX1 U289 ( .A(\mem<14><4> ), .Y(n48) );
  INVX1 U290 ( .A(net102545), .Y(net102839) );
  NAND2X1 U291 ( .A(n49), .B(net90239), .Y(n5) );
  INVX1 U293 ( .A(\mem<15><4> ), .Y(n49) );
  INVX8 U295 ( .A(net89361), .Y(net89359) );
  MUX2X1 U297 ( .B(n13), .A(n14), .S(net89359), .Y(n12) );
  MUX2X1 U299 ( .B(n29), .A(n30), .S(net89513), .Y(n13) );
  MUX2X1 U301 ( .B(n37), .A(n38), .S(net89777), .Y(n29) );
  MUX2X1 U302 ( .B(n41), .A(n42), .S(net90239), .Y(n37) );
  MUX2X1 U303 ( .B(n39), .A(n40), .S(net90241), .Y(n38) );
  INVX8 U305 ( .A(net89783), .Y(net89777) );
  MUX2X1 U307 ( .B(n31), .A(n32), .S(net89775), .Y(n30) );
  MUX2X1 U309 ( .B(n35), .A(n36), .S(net90241), .Y(n31) );
  MUX2X1 U311 ( .B(n33), .A(n34), .S(net90245), .Y(n32) );
  INVX8 U313 ( .A(net90251), .Y(net90245) );
  INVX8 U314 ( .A(net89783), .Y(net89775) );
  MUX2X1 U315 ( .B(n15), .A(n16), .S(net89513), .Y(n14) );
  MUX2X1 U317 ( .B(n23), .A(n24), .S(net89781), .Y(n15) );
  MUX2X1 U319 ( .B(n27), .A(n28), .S(net90249), .Y(n23) );
  MUX2X1 U321 ( .B(n25), .A(n26), .S(net90239), .Y(n24) );
  INVX8 U323 ( .A(net89783), .Y(net89781) );
  MUX2X1 U325 ( .B(n17), .A(n18), .S(net89781), .Y(n16) );
  MUX2X1 U326 ( .B(n21), .A(n22), .S(net90239), .Y(n17) );
  MUX2X1 U327 ( .B(n19), .A(n20), .S(net90241), .Y(n18) );
  INVX8 U329 ( .A(net89225), .Y(net89223) );
  INVX1 U331 ( .A(write), .Y(n9) );
  AND2X2 U333 ( .A(n6), .B(net85891), .Y(\data_out<3> ) );
  AND2X2 U335 ( .A(n6), .B(net86080), .Y(\data_out<0> ) );
  AND2X2 U337 ( .A(n6), .B(net85954), .Y(\data_out<2> ) );
  AND2X2 U338 ( .A(n573), .B(n574), .Y(n72) );
  AND2X2 U339 ( .A(n571), .B(n569), .Y(n74) );
  AND2X2 U342 ( .A(n712), .B(n713), .Y(n75) );
  AND2X2 U344 ( .A(n715), .B(n716), .Y(n76) );
  AND2X2 U346 ( .A(n717), .B(n718), .Y(n77) );
  AND2X2 U348 ( .A(\mem<0><4> ), .B(n585), .Y(n78) );
  INVX1 U350 ( .A(n78), .Y(n79) );
  AND2X2 U351 ( .A(\mem<0><3> ), .B(n585), .Y(n80) );
  INVX1 U352 ( .A(n80), .Y(n82) );
  AND2X2 U355 ( .A(\mem<0><2> ), .B(n585), .Y(n83) );
  INVX1 U357 ( .A(n83), .Y(n84) );
  AND2X2 U359 ( .A(\mem<0><1> ), .B(n585), .Y(n85) );
  INVX1 U361 ( .A(n85), .Y(n86) );
  AND2X2 U363 ( .A(\mem<0><0> ), .B(n585), .Y(n87) );
  INVX1 U364 ( .A(n87), .Y(n88) );
  AND2X2 U365 ( .A(\mem<1><4> ), .B(n587), .Y(n90) );
  INVX1 U368 ( .A(n90), .Y(n91) );
  AND2X2 U370 ( .A(\mem<1><3> ), .B(n587), .Y(n92) );
  INVX1 U372 ( .A(n92), .Y(n93) );
  AND2X2 U374 ( .A(\mem<1><2> ), .B(n587), .Y(n94) );
  INVX1 U376 ( .A(n94), .Y(n95) );
  AND2X2 U377 ( .A(\mem<1><1> ), .B(n587), .Y(n96) );
  INVX1 U378 ( .A(n96), .Y(n98) );
  AND2X2 U381 ( .A(\mem<1><0> ), .B(n587), .Y(n99) );
  INVX1 U383 ( .A(n99), .Y(n100) );
  AND2X2 U385 ( .A(\mem<2><4> ), .B(n589), .Y(n101) );
  INVX1 U387 ( .A(n101), .Y(n102) );
  AND2X2 U389 ( .A(\mem<2><3> ), .B(n589), .Y(n103) );
  INVX1 U390 ( .A(n103), .Y(n104) );
  AND2X2 U391 ( .A(\mem<2><2> ), .B(n589), .Y(n106) );
  INVX1 U394 ( .A(n106), .Y(n107) );
  AND2X2 U396 ( .A(\mem<2><1> ), .B(n589), .Y(n108) );
  INVX1 U398 ( .A(n108), .Y(n109) );
  AND2X2 U400 ( .A(\mem<2><0> ), .B(n589), .Y(n110) );
  INVX1 U402 ( .A(n110), .Y(n111) );
  AND2X2 U403 ( .A(\mem<3><4> ), .B(n591), .Y(n112) );
  INVX1 U404 ( .A(n112), .Y(n116) );
  AND2X2 U407 ( .A(\mem<3><3> ), .B(n591), .Y(n117) );
  INVX1 U409 ( .A(n117), .Y(n118) );
  AND2X2 U411 ( .A(\mem<3><2> ), .B(n591), .Y(n119) );
  INVX1 U413 ( .A(n119), .Y(n120) );
  AND2X2 U415 ( .A(\mem<3><1> ), .B(n591), .Y(n121) );
  INVX1 U416 ( .A(n121), .Y(n122) );
  AND2X2 U417 ( .A(\mem<3><0> ), .B(n591), .Y(n123) );
  INVX1 U420 ( .A(n123), .Y(n124) );
  AND2X2 U422 ( .A(\mem<4><4> ), .B(n593), .Y(n125) );
  INVX1 U424 ( .A(n125), .Y(n126) );
  AND2X2 U426 ( .A(\mem<4><3> ), .B(n593), .Y(n127) );
  INVX1 U428 ( .A(n127), .Y(n128) );
  AND2X2 U429 ( .A(\mem<4><2> ), .B(n593), .Y(n129) );
  INVX1 U430 ( .A(n129), .Y(n130) );
  AND2X2 U433 ( .A(\mem<4><1> ), .B(n593), .Y(n131) );
  INVX1 U434 ( .A(n131), .Y(n132) );
  AND2X2 U436 ( .A(\mem<4><0> ), .B(n593), .Y(n133) );
  INVX1 U437 ( .A(n133), .Y(n134) );
  AND2X2 U439 ( .A(\mem<5><4> ), .B(n595), .Y(n135) );
  INVX1 U440 ( .A(n135), .Y(n136) );
  AND2X2 U442 ( .A(\mem<5><3> ), .B(n595), .Y(n137) );
  INVX1 U443 ( .A(n137), .Y(n138) );
  AND2X2 U445 ( .A(\mem<5><2> ), .B(n595), .Y(n139) );
  INVX1 U446 ( .A(n139), .Y(n140) );
  AND2X2 U447 ( .A(\mem<5><1> ), .B(n595), .Y(n141) );
  INVX1 U451 ( .A(n141), .Y(n142) );
  AND2X2 U452 ( .A(\mem<5><0> ), .B(n595), .Y(n143) );
  INVX1 U453 ( .A(n143), .Y(n144) );
  AND2X2 U454 ( .A(\mem<6><4> ), .B(n597), .Y(n145) );
  INVX1 U455 ( .A(n145), .Y(n146) );
  AND2X2 U456 ( .A(\mem<6><3> ), .B(n597), .Y(n147) );
  INVX1 U457 ( .A(n147), .Y(n148) );
  AND2X2 U458 ( .A(\mem<6><2> ), .B(n597), .Y(n149) );
  INVX1 U459 ( .A(n149), .Y(n150) );
  AND2X2 U460 ( .A(\mem<6><1> ), .B(n597), .Y(n151) );
  INVX1 U461 ( .A(n151), .Y(n152) );
  AND2X2 U462 ( .A(\mem<6><0> ), .B(n597), .Y(n153) );
  INVX1 U463 ( .A(n153), .Y(n154) );
  AND2X2 U464 ( .A(\mem<7><4> ), .B(n599), .Y(n155) );
  INVX1 U465 ( .A(n155), .Y(n156) );
  AND2X2 U466 ( .A(\mem<7><3> ), .B(n599), .Y(n157) );
  INVX1 U467 ( .A(n157), .Y(n158) );
  AND2X2 U468 ( .A(\mem<7><2> ), .B(n599), .Y(n159) );
  INVX1 U469 ( .A(n159), .Y(n160) );
  AND2X2 U470 ( .A(\mem<7><1> ), .B(n599), .Y(n161) );
  INVX1 U471 ( .A(n161), .Y(n162) );
  AND2X2 U472 ( .A(\mem<7><0> ), .B(n599), .Y(n163) );
  INVX1 U473 ( .A(n163), .Y(n164) );
  AND2X2 U474 ( .A(\mem<8><4> ), .B(n601), .Y(n165) );
  INVX1 U475 ( .A(n165), .Y(n166) );
  AND2X2 U476 ( .A(\mem<8><3> ), .B(n601), .Y(n167) );
  INVX1 U477 ( .A(n167), .Y(n168) );
  AND2X2 U478 ( .A(\mem<8><2> ), .B(n601), .Y(n169) );
  INVX1 U479 ( .A(n169), .Y(n170) );
  AND2X2 U480 ( .A(\mem<8><1> ), .B(n601), .Y(n171) );
  INVX1 U481 ( .A(n171), .Y(n173) );
  AND2X2 U482 ( .A(\mem<8><0> ), .B(n601), .Y(n174) );
  INVX1 U483 ( .A(n174), .Y(n175) );
  AND2X2 U484 ( .A(\mem<9><4> ), .B(n603), .Y(n176) );
  INVX1 U485 ( .A(n176), .Y(n177) );
  AND2X2 U486 ( .A(\mem<9><3> ), .B(n603), .Y(n178) );
  INVX1 U487 ( .A(n178), .Y(n179) );
  AND2X2 U488 ( .A(\mem<9><2> ), .B(n603), .Y(n180) );
  INVX1 U489 ( .A(n180), .Y(n181) );
  AND2X2 U490 ( .A(\mem<9><1> ), .B(n603), .Y(n182) );
  INVX1 U491 ( .A(n182), .Y(n183) );
  AND2X2 U492 ( .A(\mem<9><0> ), .B(n603), .Y(n184) );
  INVX1 U493 ( .A(n184), .Y(n185) );
  AND2X2 U494 ( .A(\mem<10><4> ), .B(n605), .Y(n186) );
  INVX1 U495 ( .A(n186), .Y(n187) );
  AND2X2 U496 ( .A(\mem<10><3> ), .B(n605), .Y(n188) );
  INVX1 U497 ( .A(n188), .Y(n189) );
  AND2X2 U498 ( .A(\mem<10><2> ), .B(n605), .Y(n190) );
  INVX1 U499 ( .A(n190), .Y(n191) );
  AND2X2 U500 ( .A(\mem<10><1> ), .B(n605), .Y(n192) );
  INVX1 U501 ( .A(n192), .Y(n193) );
  AND2X2 U502 ( .A(\mem<10><0> ), .B(n605), .Y(n194) );
  INVX1 U503 ( .A(n194), .Y(n195) );
  AND2X2 U504 ( .A(\mem<11><4> ), .B(n607), .Y(n196) );
  INVX1 U505 ( .A(n196), .Y(n197) );
  AND2X2 U506 ( .A(\mem<11><3> ), .B(n607), .Y(n198) );
  INVX1 U507 ( .A(n198), .Y(n199) );
  AND2X2 U508 ( .A(\mem<11><2> ), .B(n607), .Y(n200) );
  INVX1 U509 ( .A(n200), .Y(n201) );
  AND2X2 U510 ( .A(\mem<11><1> ), .B(n607), .Y(n202) );
  INVX1 U511 ( .A(n202), .Y(n203) );
  AND2X2 U512 ( .A(\mem<11><0> ), .B(n607), .Y(n204) );
  INVX1 U513 ( .A(n204), .Y(n205) );
  AND2X2 U514 ( .A(\mem<12><4> ), .B(n609), .Y(n206) );
  INVX1 U515 ( .A(n206), .Y(n207) );
  AND2X2 U516 ( .A(\mem<12><3> ), .B(n609), .Y(n208) );
  INVX1 U517 ( .A(n208), .Y(n209) );
  AND2X2 U518 ( .A(\mem<12><2> ), .B(n609), .Y(n210) );
  INVX1 U519 ( .A(n210), .Y(n211) );
  AND2X2 U520 ( .A(\mem<12><1> ), .B(n609), .Y(n212) );
  INVX1 U521 ( .A(n212), .Y(n213) );
  AND2X2 U522 ( .A(\mem<12><0> ), .B(n609), .Y(n214) );
  INVX1 U523 ( .A(n214), .Y(n215) );
  AND2X2 U524 ( .A(\mem<13><4> ), .B(n611), .Y(n216) );
  INVX1 U525 ( .A(n216), .Y(n217) );
  AND2X2 U526 ( .A(\mem<13><3> ), .B(n611), .Y(n218) );
  INVX1 U527 ( .A(n218), .Y(n219) );
  AND2X2 U528 ( .A(\mem<13><2> ), .B(n611), .Y(n220) );
  INVX1 U529 ( .A(n220), .Y(n221) );
  AND2X2 U530 ( .A(\mem<13><1> ), .B(n611), .Y(n222) );
  INVX1 U531 ( .A(n222), .Y(n223) );
  AND2X2 U532 ( .A(\mem<13><0> ), .B(n611), .Y(n224) );
  INVX1 U533 ( .A(n224), .Y(n225) );
  AND2X2 U534 ( .A(\mem<14><4> ), .B(n613), .Y(n226) );
  INVX1 U535 ( .A(n226), .Y(n227) );
  AND2X2 U536 ( .A(\mem<14><3> ), .B(n613), .Y(n228) );
  INVX1 U537 ( .A(n228), .Y(n230) );
  AND2X2 U538 ( .A(\mem<14><2> ), .B(n613), .Y(n231) );
  INVX1 U539 ( .A(n231), .Y(n232) );
  AND2X2 U540 ( .A(\mem<14><1> ), .B(n613), .Y(n233) );
  INVX1 U541 ( .A(n233), .Y(n234) );
  AND2X2 U542 ( .A(\mem<14><0> ), .B(n613), .Y(n235) );
  INVX1 U543 ( .A(n235), .Y(n236) );
  AND2X2 U544 ( .A(\mem<15><4> ), .B(n615), .Y(n237) );
  INVX1 U545 ( .A(n237), .Y(n238) );
  AND2X2 U546 ( .A(\mem<15><3> ), .B(n615), .Y(n239) );
  INVX1 U547 ( .A(n239), .Y(n240) );
  AND2X2 U548 ( .A(\mem<15><2> ), .B(n615), .Y(n241) );
  INVX1 U549 ( .A(n241), .Y(n242) );
  AND2X2 U550 ( .A(\mem<15><1> ), .B(n615), .Y(n243) );
  INVX1 U551 ( .A(n243), .Y(n244) );
  AND2X2 U552 ( .A(\mem<15><0> ), .B(n615), .Y(n245) );
  INVX1 U553 ( .A(n245), .Y(n246) );
  AND2X2 U554 ( .A(\mem<16><4> ), .B(n617), .Y(n247) );
  INVX1 U555 ( .A(n247), .Y(n248) );
  AND2X2 U556 ( .A(\mem<16><3> ), .B(n617), .Y(n249) );
  INVX1 U557 ( .A(n249), .Y(n250) );
  AND2X2 U558 ( .A(\mem<16><2> ), .B(n617), .Y(n251) );
  INVX1 U559 ( .A(n251), .Y(n252) );
  AND2X2 U560 ( .A(\mem<16><1> ), .B(n617), .Y(n253) );
  INVX1 U561 ( .A(n253), .Y(n254) );
  AND2X2 U562 ( .A(\mem<16><0> ), .B(n617), .Y(n255) );
  INVX1 U563 ( .A(n255), .Y(n256) );
  AND2X2 U564 ( .A(\mem<17><4> ), .B(n619), .Y(n257) );
  INVX1 U565 ( .A(n257), .Y(n258) );
  AND2X2 U566 ( .A(\mem<17><3> ), .B(n619), .Y(n259) );
  INVX1 U567 ( .A(n259), .Y(n260) );
  AND2X2 U568 ( .A(\mem<17><2> ), .B(n619), .Y(n261) );
  INVX1 U569 ( .A(n261), .Y(n262) );
  AND2X2 U570 ( .A(\mem<17><1> ), .B(n619), .Y(n263) );
  INVX1 U571 ( .A(n263), .Y(n264) );
  AND2X2 U572 ( .A(\mem<17><0> ), .B(n619), .Y(n265) );
  INVX1 U573 ( .A(n265), .Y(n266) );
  AND2X2 U574 ( .A(\mem<18><4> ), .B(n621), .Y(n267) );
  INVX1 U575 ( .A(n267), .Y(n268) );
  AND2X2 U576 ( .A(\mem<18><3> ), .B(n621), .Y(n269) );
  INVX1 U577 ( .A(n269), .Y(n270) );
  AND2X2 U578 ( .A(\mem<18><2> ), .B(n621), .Y(n271) );
  INVX1 U579 ( .A(n271), .Y(n272) );
  AND2X2 U580 ( .A(\mem<18><1> ), .B(n621), .Y(n273) );
  INVX1 U581 ( .A(n273), .Y(n274) );
  AND2X2 U582 ( .A(\mem<18><0> ), .B(n621), .Y(n275) );
  INVX1 U583 ( .A(n275), .Y(n276) );
  AND2X2 U584 ( .A(\mem<19><4> ), .B(n623), .Y(n277) );
  INVX1 U585 ( .A(n277), .Y(n278) );
  AND2X2 U586 ( .A(\mem<19><3> ), .B(n623), .Y(n279) );
  INVX1 U587 ( .A(n279), .Y(n280) );
  AND2X2 U588 ( .A(\mem<19><2> ), .B(n623), .Y(n281) );
  INVX1 U589 ( .A(n281), .Y(n282) );
  AND2X2 U590 ( .A(\mem<19><1> ), .B(n623), .Y(n283) );
  INVX1 U591 ( .A(n283), .Y(n284) );
  AND2X2 U592 ( .A(\mem<19><0> ), .B(n623), .Y(n285) );
  INVX1 U593 ( .A(n285), .Y(n287) );
  AND2X2 U594 ( .A(\mem<20><4> ), .B(n625), .Y(n448) );
  INVX1 U595 ( .A(n448), .Y(n449) );
  AND2X2 U596 ( .A(\mem<20><3> ), .B(n625), .Y(n450) );
  INVX1 U597 ( .A(n450), .Y(n451) );
  AND2X2 U598 ( .A(\mem<20><2> ), .B(n625), .Y(n452) );
  INVX1 U599 ( .A(n452), .Y(n453) );
  AND2X2 U600 ( .A(\mem<20><1> ), .B(n625), .Y(n454) );
  INVX1 U601 ( .A(n454), .Y(n455) );
  AND2X2 U602 ( .A(\mem<20><0> ), .B(n625), .Y(n456) );
  INVX1 U603 ( .A(n456), .Y(n457) );
  AND2X2 U604 ( .A(\mem<21><4> ), .B(n627), .Y(n458) );
  INVX1 U605 ( .A(n458), .Y(n459) );
  AND2X2 U606 ( .A(\mem<21><3> ), .B(n627), .Y(n460) );
  INVX1 U607 ( .A(n460), .Y(n461) );
  AND2X2 U608 ( .A(\mem<21><2> ), .B(n627), .Y(n462) );
  INVX1 U609 ( .A(n462), .Y(n463) );
  AND2X2 U610 ( .A(\mem<21><1> ), .B(n627), .Y(n464) );
  INVX1 U611 ( .A(n464), .Y(n465) );
  AND2X2 U612 ( .A(\mem<21><0> ), .B(n627), .Y(n466) );
  INVX1 U613 ( .A(n466), .Y(n467) );
  AND2X2 U614 ( .A(\mem<22><4> ), .B(n629), .Y(n468) );
  INVX1 U615 ( .A(n468), .Y(n469) );
  AND2X2 U616 ( .A(\mem<22><3> ), .B(n629), .Y(n470) );
  INVX1 U617 ( .A(n470), .Y(n471) );
  AND2X2 U618 ( .A(\mem<22><2> ), .B(n629), .Y(n472) );
  INVX1 U619 ( .A(n472), .Y(n473) );
  AND2X2 U620 ( .A(\mem<22><1> ), .B(n629), .Y(n474) );
  INVX1 U621 ( .A(n474), .Y(n475) );
  AND2X2 U622 ( .A(\mem<22><0> ), .B(n629), .Y(n476) );
  INVX1 U623 ( .A(n476), .Y(n477) );
  AND2X2 U624 ( .A(\mem<23><4> ), .B(n631), .Y(n478) );
  INVX1 U625 ( .A(n478), .Y(n479) );
  AND2X2 U626 ( .A(\mem<23><3> ), .B(n631), .Y(n480) );
  INVX1 U627 ( .A(n480), .Y(n481) );
  AND2X2 U628 ( .A(\mem<23><2> ), .B(n631), .Y(n482) );
  INVX1 U629 ( .A(n482), .Y(n483) );
  AND2X2 U630 ( .A(\mem<23><1> ), .B(n631), .Y(n484) );
  INVX1 U631 ( .A(n484), .Y(n485) );
  AND2X2 U632 ( .A(\mem<23><0> ), .B(n631), .Y(n486) );
  INVX1 U633 ( .A(n486), .Y(n487) );
  AND2X2 U634 ( .A(\mem<24><4> ), .B(n633), .Y(n488) );
  INVX1 U635 ( .A(n488), .Y(n489) );
  AND2X2 U636 ( .A(\mem<24><3> ), .B(n633), .Y(n490) );
  INVX1 U637 ( .A(n490), .Y(n491) );
  AND2X2 U638 ( .A(\mem<24><2> ), .B(n633), .Y(n492) );
  INVX1 U639 ( .A(n492), .Y(n493) );
  AND2X2 U640 ( .A(\mem<24><1> ), .B(n633), .Y(n494) );
  INVX1 U641 ( .A(n494), .Y(n495) );
  AND2X2 U642 ( .A(\mem<24><0> ), .B(n633), .Y(n496) );
  INVX1 U643 ( .A(n496), .Y(n497) );
  AND2X2 U644 ( .A(\mem<25><4> ), .B(n635), .Y(n498) );
  INVX1 U645 ( .A(n498), .Y(n499) );
  AND2X2 U646 ( .A(\mem<25><3> ), .B(n635), .Y(n500) );
  INVX1 U647 ( .A(n500), .Y(n501) );
  AND2X2 U648 ( .A(\mem<25><2> ), .B(n635), .Y(n502) );
  INVX1 U649 ( .A(n502), .Y(n503) );
  AND2X2 U650 ( .A(\mem<25><1> ), .B(n635), .Y(n504) );
  INVX1 U651 ( .A(n504), .Y(n505) );
  AND2X2 U652 ( .A(\mem<25><0> ), .B(n635), .Y(n506) );
  INVX1 U653 ( .A(n506), .Y(n507) );
  AND2X2 U654 ( .A(\mem<26><4> ), .B(n637), .Y(n508) );
  INVX1 U655 ( .A(n508), .Y(n509) );
  AND2X2 U656 ( .A(\mem<26><3> ), .B(n637), .Y(n510) );
  INVX1 U657 ( .A(n510), .Y(n511) );
  AND2X2 U658 ( .A(\mem<26><2> ), .B(n637), .Y(n512) );
  INVX1 U659 ( .A(n512), .Y(n513) );
  AND2X2 U660 ( .A(\mem<26><1> ), .B(n637), .Y(n514) );
  INVX1 U661 ( .A(n514), .Y(n515) );
  AND2X2 U662 ( .A(\mem<26><0> ), .B(n637), .Y(n516) );
  INVX1 U663 ( .A(n516), .Y(n517) );
  AND2X2 U664 ( .A(\mem<27><4> ), .B(n639), .Y(n518) );
  INVX1 U665 ( .A(n518), .Y(n519) );
  AND2X2 U666 ( .A(\mem<27><3> ), .B(n639), .Y(n520) );
  INVX1 U667 ( .A(n520), .Y(n521) );
  AND2X2 U668 ( .A(\mem<27><2> ), .B(n639), .Y(n522) );
  INVX1 U669 ( .A(n522), .Y(n523) );
  AND2X2 U670 ( .A(\mem<27><1> ), .B(n639), .Y(n524) );
  INVX1 U671 ( .A(n524), .Y(n525) );
  AND2X2 U672 ( .A(\mem<27><0> ), .B(n639), .Y(n526) );
  INVX1 U673 ( .A(n526), .Y(n527) );
  AND2X2 U674 ( .A(\mem<28><4> ), .B(n641), .Y(n528) );
  INVX1 U675 ( .A(n528), .Y(n529) );
  AND2X2 U676 ( .A(\mem<28><3> ), .B(n641), .Y(n530) );
  INVX1 U677 ( .A(n530), .Y(n531) );
  AND2X2 U678 ( .A(\mem<28><2> ), .B(n641), .Y(n532) );
  INVX1 U679 ( .A(n532), .Y(n533) );
  AND2X2 U680 ( .A(\mem<28><1> ), .B(n641), .Y(n534) );
  INVX1 U681 ( .A(n534), .Y(n535) );
  AND2X2 U682 ( .A(\mem<28><0> ), .B(n641), .Y(n536) );
  INVX1 U683 ( .A(n536), .Y(n537) );
  AND2X2 U684 ( .A(\mem<29><4> ), .B(n643), .Y(n538) );
  INVX1 U685 ( .A(n538), .Y(n539) );
  AND2X2 U686 ( .A(\mem<29><3> ), .B(n643), .Y(n540) );
  INVX1 U687 ( .A(n540), .Y(n541) );
  AND2X2 U688 ( .A(\mem<29><2> ), .B(n643), .Y(n542) );
  INVX1 U689 ( .A(n542), .Y(n543) );
  AND2X2 U690 ( .A(\mem<29><1> ), .B(n643), .Y(n544) );
  INVX1 U691 ( .A(n544), .Y(n545) );
  AND2X2 U692 ( .A(\mem<29><0> ), .B(n643), .Y(n546) );
  INVX1 U693 ( .A(n546), .Y(n547) );
  AND2X2 U694 ( .A(\mem<30><4> ), .B(n645), .Y(n548) );
  INVX1 U695 ( .A(n548), .Y(n549) );
  AND2X2 U696 ( .A(\mem<30><3> ), .B(n645), .Y(n550) );
  INVX1 U697 ( .A(n550), .Y(n551) );
  AND2X2 U698 ( .A(\mem<30><2> ), .B(n645), .Y(n552) );
  INVX1 U699 ( .A(n552), .Y(n553) );
  AND2X2 U700 ( .A(\mem<30><1> ), .B(n645), .Y(n554) );
  INVX1 U701 ( .A(n554), .Y(n555) );
  AND2X2 U702 ( .A(\mem<30><0> ), .B(n645), .Y(n556) );
  INVX1 U703 ( .A(n556), .Y(n557) );
  AND2X2 U704 ( .A(\mem<31><4> ), .B(n647), .Y(n558) );
  INVX1 U705 ( .A(n558), .Y(n559) );
  AND2X2 U706 ( .A(\mem<31><3> ), .B(n647), .Y(n560) );
  INVX1 U707 ( .A(n560), .Y(n561) );
  AND2X2 U708 ( .A(\mem<31><2> ), .B(n647), .Y(n562) );
  INVX1 U709 ( .A(n562), .Y(n563) );
  AND2X2 U710 ( .A(\mem<31><1> ), .B(n647), .Y(n564) );
  INVX1 U711 ( .A(n564), .Y(n565) );
  AND2X2 U712 ( .A(\mem<31><0> ), .B(n647), .Y(n566) );
  INVX1 U713 ( .A(n566), .Y(n567) );
  AND2X2 U714 ( .A(net89511), .B(n872), .Y(n568) );
  INVX1 U715 ( .A(n568), .Y(n569) );
  AND2X2 U716 ( .A(n873), .B(net102667), .Y(n570) );
  INVX1 U717 ( .A(n570), .Y(n571) );
  AND2X1 U718 ( .A(n845), .B(net90935), .Y(n572) );
  INVX1 U719 ( .A(net121526), .Y(net121576) );
  INVX1 U720 ( .A(write), .Y(net121526) );
  INVX1 U721 ( .A(net90251), .Y(net121136) );
  MUX2X1 U722 ( .B(n825), .A(n826), .S(net89515), .Y(n842) );
  INVX1 U723 ( .A(net90255), .Y(net121143) );
  MUX2X1 U724 ( .B(n863), .A(n862), .S(net121110), .Y(n864) );
  MUX2X1 U725 ( .B(n924), .A(n925), .S(net117994), .Y(n929) );
  MUX2X1 U726 ( .B(n918), .A(n919), .S(net89515), .Y(n933) );
  MUX2X1 U727 ( .B(n870), .A(n871), .S(net89783), .Y(n872) );
  INVX1 U728 ( .A(net90251), .Y(net121110) );
  MUX2X1 U729 ( .B(n861), .A(n860), .S(net102545), .Y(n865) );
  NAND2X1 U730 ( .A(n878), .B(net121144), .Y(n573) );
  NAND2X1 U731 ( .A(n877), .B(net121136), .Y(n574) );
  INVX1 U732 ( .A(\mem<18><2> ), .Y(n878) );
  INVX1 U733 ( .A(\mem<19><2> ), .Y(n877) );
  MUX2X1 U734 ( .B(n850), .A(n851), .S(net89783), .Y(n859) );
  INVX1 U735 ( .A(net102846), .Y(net117952) );
  MUX2X1 U736 ( .B(n902), .A(n903), .S(net89361), .Y(n904) );
  BUFX2 U737 ( .A(n286), .Y(n575) );
  INVX1 U738 ( .A(n575), .Y(n966) );
  BUFX2 U739 ( .A(n229), .Y(n576) );
  INVX1 U740 ( .A(n576), .Y(n967) );
  BUFX2 U741 ( .A(n172), .Y(n577) );
  INVX1 U742 ( .A(n577), .Y(n968) );
  BUFX2 U743 ( .A(n114), .Y(n578) );
  INVX1 U744 ( .A(n578), .Y(n969) );
  AND2X1 U745 ( .A(\data_in<4> ), .B(n56), .Y(n579) );
  AND2X1 U746 ( .A(\data_in<3> ), .B(n56), .Y(n580) );
  AND2X1 U747 ( .A(\data_in<2> ), .B(n56), .Y(n581) );
  AND2X1 U748 ( .A(\data_in<1> ), .B(n56), .Y(n582) );
  AND2X1 U749 ( .A(\data_in<0> ), .B(n56), .Y(n583) );
  AND2X1 U750 ( .A(n650), .B(n56), .Y(n584) );
  INVX1 U751 ( .A(n584), .Y(n585) );
  AND2X1 U752 ( .A(n652), .B(n56), .Y(n586) );
  INVX1 U753 ( .A(n586), .Y(n587) );
  AND2X1 U754 ( .A(n654), .B(n56), .Y(n588) );
  INVX1 U755 ( .A(n588), .Y(n589) );
  AND2X1 U756 ( .A(n656), .B(n56), .Y(n590) );
  INVX1 U757 ( .A(n590), .Y(n591) );
  AND2X1 U758 ( .A(n658), .B(n56), .Y(n592) );
  INVX1 U759 ( .A(n592), .Y(n593) );
  AND2X1 U760 ( .A(n660), .B(n56), .Y(n594) );
  INVX1 U761 ( .A(n594), .Y(n595) );
  AND2X1 U762 ( .A(n662), .B(n56), .Y(n596) );
  INVX1 U763 ( .A(n596), .Y(n597) );
  AND2X1 U764 ( .A(n664), .B(n56), .Y(n598) );
  INVX1 U765 ( .A(n598), .Y(n599) );
  AND2X1 U766 ( .A(n666), .B(n56), .Y(n600) );
  INVX1 U767 ( .A(n600), .Y(n601) );
  AND2X1 U768 ( .A(n668), .B(n56), .Y(n602) );
  INVX1 U769 ( .A(n602), .Y(n603) );
  AND2X1 U770 ( .A(n670), .B(n56), .Y(n604) );
  INVX1 U771 ( .A(n604), .Y(n605) );
  AND2X1 U772 ( .A(n673), .B(n56), .Y(n606) );
  INVX1 U773 ( .A(n606), .Y(n607) );
  AND2X1 U774 ( .A(n674), .B(n56), .Y(n608) );
  INVX1 U775 ( .A(n608), .Y(n609) );
  AND2X1 U776 ( .A(n677), .B(n56), .Y(n610) );
  INVX1 U777 ( .A(n610), .Y(n611) );
  AND2X1 U778 ( .A(n678), .B(n56), .Y(n612) );
  INVX1 U779 ( .A(n612), .Y(n613) );
  AND2X1 U780 ( .A(n680), .B(n56), .Y(n614) );
  INVX1 U781 ( .A(n614), .Y(n615) );
  AND2X1 U782 ( .A(n683), .B(n56), .Y(n616) );
  INVX1 U783 ( .A(n616), .Y(n617) );
  AND2X1 U784 ( .A(n685), .B(n56), .Y(n618) );
  INVX1 U785 ( .A(n618), .Y(n619) );
  AND2X1 U786 ( .A(n686), .B(n56), .Y(n620) );
  INVX1 U787 ( .A(n620), .Y(n621) );
  AND2X1 U788 ( .A(n688), .B(n56), .Y(n622) );
  INVX1 U789 ( .A(n622), .Y(n623) );
  AND2X1 U790 ( .A(n690), .B(n56), .Y(n624) );
  INVX1 U791 ( .A(n624), .Y(n625) );
  AND2X1 U792 ( .A(n692), .B(n56), .Y(n626) );
  INVX1 U793 ( .A(n626), .Y(n627) );
  AND2X1 U794 ( .A(n695), .B(n56), .Y(n628) );
  INVX1 U795 ( .A(n628), .Y(n629) );
  AND2X1 U796 ( .A(n697), .B(n56), .Y(n630) );
  INVX1 U797 ( .A(n630), .Y(n631) );
  AND2X1 U798 ( .A(n698), .B(n56), .Y(n632) );
  INVX1 U799 ( .A(n632), .Y(n633) );
  AND2X1 U800 ( .A(n700), .B(n56), .Y(n634) );
  INVX1 U801 ( .A(n634), .Y(n635) );
  AND2X1 U802 ( .A(n702), .B(n56), .Y(n636) );
  INVX1 U803 ( .A(n636), .Y(n637) );
  AND2X1 U804 ( .A(n704), .B(n56), .Y(n638) );
  INVX1 U805 ( .A(n638), .Y(n639) );
  AND2X1 U806 ( .A(n706), .B(n56), .Y(n640) );
  INVX1 U807 ( .A(n640), .Y(n641) );
  AND2X1 U808 ( .A(n708), .B(n56), .Y(n642) );
  INVX1 U809 ( .A(n642), .Y(n643) );
  AND2X1 U810 ( .A(n710), .B(n56), .Y(n644) );
  INVX1 U811 ( .A(n644), .Y(n645) );
  AND2X1 U812 ( .A(n649), .B(n56), .Y(n646) );
  INVX1 U813 ( .A(n646), .Y(n647) );
  INVX1 U814 ( .A(n649), .Y(n648) );
  AND2X1 U815 ( .A(n57), .B(n969), .Y(n649) );
  AND2X1 U816 ( .A(n966), .B(n113), .Y(n650) );
  INVX1 U817 ( .A(n650), .Y(n651) );
  AND2X1 U818 ( .A(n966), .B(n105), .Y(n652) );
  INVX1 U819 ( .A(n652), .Y(n653) );
  AND2X1 U820 ( .A(n966), .B(n97), .Y(n654) );
  INVX1 U821 ( .A(n654), .Y(n655) );
  AND2X1 U822 ( .A(n966), .B(n89), .Y(n656) );
  INVX1 U823 ( .A(n656), .Y(n657) );
  AND2X1 U824 ( .A(n966), .B(n81), .Y(n658) );
  INVX1 U825 ( .A(n658), .Y(n659) );
  AND2X1 U826 ( .A(n966), .B(n73), .Y(n660) );
  INVX1 U827 ( .A(n660), .Y(n661) );
  AND2X1 U828 ( .A(n966), .B(n65), .Y(n662) );
  INVX1 U829 ( .A(n662), .Y(n663) );
  AND2X1 U830 ( .A(n966), .B(n57), .Y(n664) );
  INVX1 U831 ( .A(n664), .Y(n665) );
  AND2X1 U832 ( .A(n967), .B(n113), .Y(n666) );
  INVX1 U833 ( .A(n666), .Y(n667) );
  AND2X1 U834 ( .A(n967), .B(n105), .Y(n668) );
  INVX1 U835 ( .A(n668), .Y(n669) );
  AND2X1 U836 ( .A(n967), .B(n97), .Y(n670) );
  INVX1 U837 ( .A(n670), .Y(n671) );
  INVX1 U838 ( .A(n673), .Y(n672) );
  AND2X1 U839 ( .A(n967), .B(n89), .Y(n673) );
  AND2X1 U840 ( .A(n967), .B(n81), .Y(n674) );
  INVX1 U841 ( .A(n674), .Y(n675) );
  INVX1 U842 ( .A(n677), .Y(n676) );
  AND2X1 U843 ( .A(n967), .B(n73), .Y(n677) );
  AND2X1 U844 ( .A(n967), .B(n65), .Y(n678) );
  INVX1 U845 ( .A(n678), .Y(n679) );
  AND2X1 U846 ( .A(n967), .B(n57), .Y(n680) );
  INVX1 U847 ( .A(n680), .Y(n681) );
  INVX1 U848 ( .A(n683), .Y(n682) );
  AND2X1 U849 ( .A(n968), .B(n113), .Y(n683) );
  INVX1 U850 ( .A(n685), .Y(n684) );
  AND2X1 U851 ( .A(n968), .B(n105), .Y(n685) );
  AND2X1 U852 ( .A(n968), .B(n97), .Y(n686) );
  INVX1 U853 ( .A(n686), .Y(n687) );
  AND2X1 U854 ( .A(n968), .B(n89), .Y(n688) );
  INVX1 U855 ( .A(n688), .Y(n689) );
  AND2X1 U856 ( .A(n968), .B(n81), .Y(n690) );
  INVX1 U857 ( .A(n690), .Y(n691) );
  AND2X1 U858 ( .A(n968), .B(n73), .Y(n692) );
  INVX1 U859 ( .A(n692), .Y(n693) );
  INVX1 U860 ( .A(n695), .Y(n694) );
  AND2X1 U861 ( .A(n968), .B(n65), .Y(n695) );
  INVX1 U862 ( .A(n697), .Y(n696) );
  AND2X1 U863 ( .A(n968), .B(n57), .Y(n697) );
  AND2X1 U864 ( .A(n113), .B(n969), .Y(n698) );
  INVX1 U865 ( .A(n698), .Y(n699) );
  AND2X1 U866 ( .A(n105), .B(n969), .Y(n700) );
  INVX1 U867 ( .A(n700), .Y(n701) );
  AND2X1 U868 ( .A(n97), .B(n969), .Y(n702) );
  INVX1 U869 ( .A(n702), .Y(n703) );
  AND2X1 U870 ( .A(n89), .B(n969), .Y(n704) );
  INVX1 U871 ( .A(n704), .Y(n705) );
  AND2X1 U872 ( .A(n81), .B(n969), .Y(n706) );
  INVX1 U873 ( .A(n706), .Y(n707) );
  AND2X1 U874 ( .A(n73), .B(n969), .Y(n708) );
  INVX1 U875 ( .A(n708), .Y(n709) );
  AND2X1 U876 ( .A(n65), .B(n969), .Y(n710) );
  INVX1 U877 ( .A(n710), .Y(n711) );
  INVX1 U878 ( .A(net102831), .Y(net103275) );
  MUX2X1 U879 ( .B(n846), .A(n847), .S(net121144), .Y(n851) );
  INVX1 U880 ( .A(net121143), .Y(net102846) );
  INVX1 U881 ( .A(net102546), .Y(net102837) );
  INVX1 U882 ( .A(net102837), .Y(net102831) );
  INVX1 U883 ( .A(net90255), .Y(net102825) );
  MUX2X1 U884 ( .B(n757), .A(n758), .S(net89783), .Y(n766) );
  INVX8 U885 ( .A(N10), .Y(net90251) );
  INVX4 U886 ( .A(N10), .Y(net90255) );
  INVX1 U887 ( .A(net89511), .Y(net102667) );
  MUX2X1 U888 ( .B(n771), .A(n772), .S(net89783), .Y(n780) );
  MUX2X1 U889 ( .B(n783), .A(n784), .S(net89225), .Y(net86080) );
  NAND2X1 U890 ( .A(n805), .B(net90251), .Y(n712) );
  NAND2X1 U891 ( .A(n804), .B(net121136), .Y(n713) );
  INVX1 U892 ( .A(\mem<12><1> ), .Y(n805) );
  INVX1 U893 ( .A(\mem<13><1> ), .Y(n804) );
  MUX2X1 U894 ( .B(n808), .A(n75), .S(net89783), .Y(n809) );
  MUX2X1 U895 ( .B(n799), .A(n800), .S(net90255), .Y(n803) );
  INVX1 U896 ( .A(net90255), .Y(net102545) );
  INVX1 U897 ( .A(net102545), .Y(net102546) );
  INVX1 U898 ( .A(n714), .Y(n922) );
  MUX2X1 U899 ( .B(n724), .A(n725), .S(net90255), .Y(n729) );
  MUX2X1 U900 ( .B(\mem<11><3> ), .A(\mem<10><3> ), .S(net102839), .Y(n714) );
  NAND2X1 U901 ( .A(n741), .B(net96102), .Y(n715) );
  NAND2X1 U902 ( .A(n740), .B(net90245), .Y(n716) );
  INVX1 U903 ( .A(net90243), .Y(net96102) );
  INVX1 U904 ( .A(\mem<10><0> ), .Y(n741) );
  INVX1 U905 ( .A(\mem<11><0> ), .Y(n740) );
  NAND2X1 U906 ( .A(n802), .B(net102846), .Y(n717) );
  NAND2X1 U907 ( .A(n801), .B(net90243), .Y(n718) );
  INVX1 U908 ( .A(\mem<10><1> ), .Y(n802) );
  INVX1 U909 ( .A(\mem<11><1> ), .Y(n801) );
  INVX8 U910 ( .A(net89515), .Y(net89511) );
  INVX8 U911 ( .A(N12), .Y(net89515) );
  INVX8 U912 ( .A(N13), .Y(net89361) );
  INVX8 U913 ( .A(N14), .Y(net89225) );
  MUX2X1 U914 ( .B(n727), .A(n726), .S(net90247), .Y(n728) );
  MUX2X1 U915 ( .B(n729), .A(n728), .S(net89775), .Y(n737) );
  MUX2X1 U916 ( .B(n731), .A(n730), .S(net90243), .Y(n735) );
  MUX2X1 U917 ( .B(n733), .A(n732), .S(net121136), .Y(n734) );
  MUX2X1 U918 ( .B(n735), .A(n734), .S(net89777), .Y(n736) );
  MUX2X1 U919 ( .B(n737), .A(n736), .S(net89511), .Y(n752) );
  MUX2X1 U920 ( .B(n739), .A(n738), .S(net90249), .Y(n742) );
  MUX2X1 U921 ( .B(n742), .A(n76), .S(net89775), .Y(n750) );
  MUX2X1 U922 ( .B(n744), .A(n743), .S(net90243), .Y(n748) );
  MUX2X1 U923 ( .B(n746), .A(n745), .S(net90239), .Y(n747) );
  MUX2X1 U924 ( .B(n748), .A(n747), .S(net89775), .Y(n749) );
  MUX2X1 U925 ( .B(n750), .A(n749), .S(net89511), .Y(n751) );
  MUX2X1 U926 ( .B(n752), .A(n751), .S(net89359), .Y(n784) );
  MUX2X1 U927 ( .B(n754), .A(n753), .S(net90247), .Y(n758) );
  MUX2X1 U928 ( .B(n756), .A(n755), .S(net90243), .Y(n757) );
  MUX2X1 U929 ( .B(n760), .A(n759), .S(net90245), .Y(n764) );
  MUX2X1 U930 ( .B(n762), .A(n761), .S(net90247), .Y(n763) );
  MUX2X1 U931 ( .B(n764), .A(n763), .S(net89777), .Y(n765) );
  MUX2X1 U932 ( .B(n766), .A(n765), .S(net89511), .Y(n782) );
  MUX2X1 U933 ( .B(n768), .A(n767), .S(net90249), .Y(n772) );
  MUX2X1 U934 ( .B(n770), .A(n769), .S(net90247), .Y(n771) );
  MUX2X1 U935 ( .B(n774), .A(n773), .S(net90247), .Y(n778) );
  MUX2X1 U936 ( .B(n776), .A(n775), .S(net90247), .Y(n777) );
  MUX2X1 U937 ( .B(n778), .A(n777), .S(net89781), .Y(n779) );
  MUX2X1 U938 ( .B(n780), .A(n779), .S(net89511), .Y(n781) );
  MUX2X1 U939 ( .B(n782), .A(n781), .S(net89359), .Y(n783) );
  MUX2X1 U940 ( .B(n786), .A(n785), .S(net90249), .Y(n790) );
  MUX2X1 U941 ( .B(n788), .A(n787), .S(net90249), .Y(n789) );
  MUX2X1 U942 ( .B(n790), .A(n789), .S(net89777), .Y(n798) );
  MUX2X1 U943 ( .B(n792), .A(n791), .S(net90247), .Y(n796) );
  MUX2X1 U944 ( .B(n794), .A(n793), .S(net90247), .Y(n795) );
  MUX2X1 U945 ( .B(n796), .A(n795), .S(net89777), .Y(n797) );
  MUX2X1 U946 ( .B(n798), .A(n797), .S(net89511), .Y(n812) );
  MUX2X1 U947 ( .B(n803), .A(n77), .S(net89777), .Y(n810) );
  MUX2X1 U948 ( .B(n807), .A(n806), .S(net90243), .Y(n808) );
  MUX2X1 U949 ( .B(n810), .A(n809), .S(net89511), .Y(n811) );
  MUX2X1 U950 ( .B(n812), .A(n811), .S(net89359), .Y(n844) );
  MUX2X1 U951 ( .B(n814), .A(n813), .S(net90245), .Y(n818) );
  MUX2X1 U952 ( .B(n816), .A(n815), .S(net90243), .Y(n817) );
  MUX2X1 U953 ( .B(n818), .A(n817), .S(net89775), .Y(n826) );
  MUX2X1 U954 ( .B(n820), .A(n819), .S(net90243), .Y(n824) );
  MUX2X1 U955 ( .B(n822), .A(n821), .S(net90243), .Y(n823) );
  MUX2X1 U956 ( .B(n824), .A(n823), .S(net89775), .Y(n825) );
  MUX2X1 U957 ( .B(n828), .A(n827), .S(net90245), .Y(n832) );
  MUX2X1 U958 ( .B(n830), .A(n829), .S(net90247), .Y(n831) );
  MUX2X1 U959 ( .B(n832), .A(n831), .S(net89781), .Y(n840) );
  MUX2X1 U960 ( .B(n834), .A(n833), .S(net90245), .Y(n838) );
  MUX2X1 U961 ( .B(n836), .A(n835), .S(net90243), .Y(n837) );
  MUX2X1 U962 ( .B(n838), .A(n837), .S(net89775), .Y(n839) );
  MUX2X1 U963 ( .B(n840), .A(n839), .S(net89511), .Y(n841) );
  MUX2X1 U964 ( .B(n842), .A(n841), .S(net89359), .Y(n843) );
  MUX2X1 U965 ( .B(n844), .A(n843), .S(net89223), .Y(n845) );
  AND2X2 U966 ( .A(net121526), .B(n572), .Y(\data_out<1> ) );
  MUX2X1 U967 ( .B(n849), .A(n848), .S(net90249), .Y(n850) );
  MUX2X1 U968 ( .B(n853), .A(n852), .S(net90241), .Y(n857) );
  MUX2X1 U969 ( .B(n855), .A(n854), .S(net90247), .Y(n856) );
  MUX2X1 U970 ( .B(n857), .A(n856), .S(net89775), .Y(n858) );
  MUX2X1 U971 ( .B(n859), .A(n858), .S(net89511), .Y(n874) );
  MUX2X1 U972 ( .B(n865), .A(n864), .S(net89781), .Y(n873) );
  MUX2X1 U973 ( .B(n867), .A(n866), .S(net90245), .Y(n871) );
  MUX2X1 U974 ( .B(n869), .A(n868), .S(net90249), .Y(n870) );
  MUX2X1 U975 ( .B(n874), .A(n74), .S(net89359), .Y(n905) );
  MUX2X1 U976 ( .B(n876), .A(n875), .S(net90245), .Y(n879) );
  MUX2X1 U977 ( .B(n879), .A(n72), .S(net89781), .Y(n887) );
  MUX2X1 U978 ( .B(n881), .A(n880), .S(net90243), .Y(n885) );
  MUX2X1 U979 ( .B(n883), .A(n882), .S(net90245), .Y(n884) );
  MUX2X1 U980 ( .B(n885), .A(n884), .S(net89777), .Y(n886) );
  MUX2X1 U981 ( .B(n887), .A(n886), .S(net89511), .Y(n903) );
  MUX2X1 U982 ( .B(n889), .A(n888), .S(net90239), .Y(n893) );
  MUX2X1 U983 ( .B(n891), .A(n890), .S(net90241), .Y(n892) );
  MUX2X1 U984 ( .B(n893), .A(n892), .S(net89775), .Y(n901) );
  MUX2X1 U985 ( .B(n895), .A(n894), .S(net90245), .Y(n899) );
  MUX2X1 U986 ( .B(n897), .A(n896), .S(net90241), .Y(n898) );
  MUX2X1 U987 ( .B(n899), .A(n898), .S(net89777), .Y(n900) );
  MUX2X1 U988 ( .B(n901), .A(n900), .S(net89511), .Y(n902) );
  MUX2X1 U989 ( .B(n905), .A(n904), .S(net89223), .Y(net85954) );
  MUX2X1 U990 ( .B(n907), .A(n906), .S(net90239), .Y(n911) );
  MUX2X1 U991 ( .B(n909), .A(n908), .S(net90239), .Y(n910) );
  MUX2X1 U992 ( .B(n911), .A(n910), .S(net89779), .Y(n919) );
  MUX2X1 U993 ( .B(n913), .A(n912), .S(net90239), .Y(n917) );
  MUX2X1 U994 ( .B(n915), .A(n914), .S(net90241), .Y(n916) );
  MUX2X1 U995 ( .B(n917), .A(n916), .S(net89779), .Y(n918) );
  MUX2X1 U996 ( .B(n921), .A(n920), .S(net90241), .Y(n923) );
  MUX2X1 U997 ( .B(n923), .A(n922), .S(net89779), .Y(n931) );
  MUX2X1 U998 ( .B(n927), .A(n926), .S(net90241), .Y(n928) );
  MUX2X1 U999 ( .B(n929), .A(n928), .S(net89779), .Y(n930) );
  MUX2X1 U1000 ( .B(n931), .A(n930), .S(net89513), .Y(n932) );
  MUX2X1 U1001 ( .B(n933), .A(n932), .S(net89359), .Y(n965) );
  MUX2X1 U1002 ( .B(n935), .A(n934), .S(net90239), .Y(n939) );
  MUX2X1 U1003 ( .B(n937), .A(n936), .S(net117952), .Y(n938) );
  MUX2X1 U1004 ( .B(n939), .A(n938), .S(net89779), .Y(n947) );
  MUX2X1 U1005 ( .B(n941), .A(n940), .S(net90247), .Y(n945) );
  MUX2X1 U1006 ( .B(n943), .A(n942), .S(net102837), .Y(n944) );
  MUX2X1 U1007 ( .B(n945), .A(n944), .S(net89779), .Y(n946) );
  MUX2X1 U1008 ( .B(n947), .A(n946), .S(net89513), .Y(n963) );
  MUX2X1 U1009 ( .B(n949), .A(n948), .S(net90245), .Y(n953) );
  MUX2X1 U1010 ( .B(n951), .A(n950), .S(net90239), .Y(n952) );
  MUX2X1 U1011 ( .B(n953), .A(n952), .S(net89779), .Y(n961) );
  MUX2X1 U1012 ( .B(n955), .A(n954), .S(net90239), .Y(n959) );
  MUX2X1 U1013 ( .B(n957), .A(n956), .S(net102825), .Y(n958) );
  MUX2X1 U1014 ( .B(n959), .A(n958), .S(net89779), .Y(n960) );
  MUX2X1 U1015 ( .B(n961), .A(n960), .S(net89513), .Y(n962) );
  MUX2X1 U1016 ( .B(n963), .A(n962), .S(net89359), .Y(n964) );
  MUX2X1 U1017 ( .B(n965), .A(n964), .S(net89223), .Y(net85891) );
endmodule


module memc_Size1_1 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , N17, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n92), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n91), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n90), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n89), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n88), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n87), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n86), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n85), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n84), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n83), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n82), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n81), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n80), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n79), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n78), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n77), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n76), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n75), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n74), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n73), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n72), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n71), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n70), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n69), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n68), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n67), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n66), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n65), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n64), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n63), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n62), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n61), .CLK(clk), .Q(\mem<31><0> ) );
  INVX1 U2 ( .A(n163), .Y(n151) );
  INVX1 U3 ( .A(n150), .Y(N17) );
  INVX1 U4 ( .A(N12), .Y(n165) );
  INVX1 U5 ( .A(n169), .Y(n2) );
  AND2X1 U6 ( .A(n161), .B(n96), .Y(n117) );
  INVX1 U7 ( .A(n160), .Y(n152) );
  INVX2 U8 ( .A(n5), .Y(n157) );
  INVX2 U9 ( .A(n1), .Y(n156) );
  INVX4 U10 ( .A(n3), .Y(n187) );
  NOR3X1 U11 ( .A(n4), .B(n103), .C(n2), .Y(n1) );
  INVX1 U12 ( .A(n167), .Y(n4) );
  NOR3X1 U13 ( .A(n169), .B(n9), .C(n4), .Y(n3) );
  INVX1 U14 ( .A(n169), .Y(n168) );
  NOR3X1 U15 ( .A(n167), .B(n9), .C(N14), .Y(n5) );
  INVX1 U16 ( .A(n167), .Y(n166) );
  INVX1 U17 ( .A(N13), .Y(n167) );
  INVX1 U18 ( .A(N14), .Y(n169) );
  OR2X2 U19 ( .A(n98), .B(write), .Y(n6) );
  INVX1 U20 ( .A(n6), .Y(\data_out<0> ) );
  OR2X2 U21 ( .A(n100), .B(n94), .Y(n8) );
  OR2X2 U22 ( .A(\addr<5> ), .B(n8), .Y(n9) );
  INVX1 U23 ( .A(n9), .Y(n10) );
  AND2X2 U24 ( .A(n119), .B(n59), .Y(n11) );
  INVX1 U25 ( .A(n11), .Y(n12) );
  AND2X2 U26 ( .A(n115), .B(n59), .Y(n13) );
  INVX1 U27 ( .A(n13), .Y(n14) );
  AND2X2 U28 ( .A(n104), .B(n59), .Y(n15) );
  INVX1 U29 ( .A(n15), .Y(n16) );
  AND2X2 U30 ( .A(n106), .B(n59), .Y(n17) );
  INVX1 U31 ( .A(n17), .Y(n18) );
  AND2X2 U32 ( .A(n108), .B(n59), .Y(n19) );
  INVX1 U33 ( .A(n19), .Y(n20) );
  AND2X2 U34 ( .A(n110), .B(n59), .Y(n21) );
  INVX1 U35 ( .A(n21), .Y(n22) );
  AND2X2 U36 ( .A(n112), .B(n59), .Y(n23) );
  INVX1 U37 ( .A(n23), .Y(n24) );
  AND2X2 U38 ( .A(n117), .B(n59), .Y(n25) );
  INVX1 U39 ( .A(n25), .Y(n26) );
  AND2X2 U40 ( .A(n119), .B(n60), .Y(n27) );
  INVX1 U41 ( .A(n27), .Y(n28) );
  AND2X2 U42 ( .A(n115), .B(n60), .Y(n29) );
  INVX1 U43 ( .A(n29), .Y(n30) );
  AND2X2 U44 ( .A(n104), .B(n60), .Y(n31) );
  INVX1 U45 ( .A(n31), .Y(n32) );
  AND2X2 U46 ( .A(n106), .B(n60), .Y(n33) );
  INVX1 U47 ( .A(n33), .Y(n34) );
  AND2X2 U48 ( .A(n108), .B(n60), .Y(n35) );
  INVX1 U49 ( .A(n35), .Y(n36) );
  AND2X2 U50 ( .A(n110), .B(n60), .Y(n37) );
  INVX1 U51 ( .A(n37), .Y(n38) );
  AND2X2 U52 ( .A(n112), .B(n60), .Y(n39) );
  INVX1 U53 ( .A(n39), .Y(n40) );
  AND2X2 U54 ( .A(n117), .B(n60), .Y(n41) );
  INVX1 U55 ( .A(n41), .Y(n42) );
  AND2X2 U56 ( .A(n119), .B(n93), .Y(n43) );
  INVX1 U57 ( .A(n43), .Y(n44) );
  AND2X2 U58 ( .A(n115), .B(n93), .Y(n45) );
  INVX1 U59 ( .A(n45), .Y(n46) );
  AND2X2 U60 ( .A(n104), .B(n93), .Y(n47) );
  INVX1 U61 ( .A(n47), .Y(n48) );
  AND2X2 U62 ( .A(n106), .B(n93), .Y(n49) );
  INVX1 U63 ( .A(n49), .Y(n50) );
  AND2X2 U64 ( .A(n108), .B(n93), .Y(n51) );
  INVX1 U65 ( .A(n51), .Y(n52) );
  AND2X2 U66 ( .A(n110), .B(n93), .Y(n53) );
  INVX1 U67 ( .A(n53), .Y(n54) );
  AND2X2 U68 ( .A(n112), .B(n93), .Y(n55) );
  INVX1 U69 ( .A(n55), .Y(n56) );
  AND2X2 U70 ( .A(n117), .B(n93), .Y(n57) );
  INVX1 U71 ( .A(n57), .Y(n58) );
  AND2X2 U72 ( .A(\data_in<0> ), .B(n3), .Y(n59) );
  AND2X2 U73 ( .A(\data_in<0> ), .B(n5), .Y(n60) );
  AND2X2 U74 ( .A(\data_in<0> ), .B(n1), .Y(n93) );
  INVX1 U75 ( .A(n165), .Y(n164) );
  INVX1 U76 ( .A(n163), .Y(n162) );
  INVX1 U77 ( .A(n161), .Y(n160) );
  INVX2 U78 ( .A(n154), .Y(n155) );
  OR2X1 U79 ( .A(n102), .B(n99), .Y(n94) );
  OR2X1 U80 ( .A(n162), .B(n164), .Y(n95) );
  INVX1 U81 ( .A(n95), .Y(n96) );
  AND2X1 U82 ( .A(N17), .B(n159), .Y(n97) );
  INVX1 U83 ( .A(n97), .Y(n98) );
  INVX1 U84 ( .A(n159), .Y(n99) );
  INVX1 U85 ( .A(write), .Y(n100) );
  INVX1 U86 ( .A(rst), .Y(n159) );
  AND2X1 U87 ( .A(n164), .B(n162), .Y(n101) );
  OR2X1 U88 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n102) );
  INVX1 U89 ( .A(n10), .Y(n103) );
  INVX1 U90 ( .A(n105), .Y(n104) );
  BUFX2 U91 ( .A(n199), .Y(n105) );
  INVX1 U92 ( .A(n107), .Y(n106) );
  BUFX2 U93 ( .A(n201), .Y(n107) );
  INVX1 U94 ( .A(n109), .Y(n108) );
  BUFX2 U95 ( .A(n203), .Y(n109) );
  INVX1 U96 ( .A(n111), .Y(n110) );
  BUFX2 U97 ( .A(n205), .Y(n111) );
  INVX1 U98 ( .A(n113), .Y(n112) );
  BUFX2 U99 ( .A(n207), .Y(n113) );
  INVX1 U100 ( .A(n115), .Y(n114) );
  AND2X1 U101 ( .A(n161), .B(n101), .Y(n115) );
  INVX1 U102 ( .A(n117), .Y(n116) );
  INVX1 U103 ( .A(n119), .Y(n118) );
  AND2X1 U104 ( .A(n160), .B(n101), .Y(n119) );
  INVX1 U105 ( .A(N11), .Y(n163) );
  MUX2X1 U106 ( .B(n121), .A(n122), .S(n151), .Y(n120) );
  MUX2X1 U107 ( .B(n124), .A(n125), .S(n151), .Y(n123) );
  MUX2X1 U108 ( .B(n127), .A(n128), .S(n151), .Y(n126) );
  MUX2X1 U109 ( .B(n130), .A(n131), .S(n151), .Y(n129) );
  MUX2X1 U110 ( .B(n133), .A(n134), .S(n166), .Y(n132) );
  MUX2X1 U111 ( .B(n136), .A(n137), .S(n151), .Y(n135) );
  MUX2X1 U112 ( .B(n139), .A(n140), .S(n151), .Y(n138) );
  MUX2X1 U113 ( .B(n142), .A(n143), .S(n151), .Y(n141) );
  MUX2X1 U114 ( .B(n145), .A(n146), .S(n151), .Y(n144) );
  MUX2X1 U115 ( .B(n148), .A(n149), .S(n166), .Y(n147) );
  MUX2X1 U116 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n153), .Y(n122) );
  MUX2X1 U117 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n153), .Y(n121) );
  MUX2X1 U118 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n153), .Y(n125) );
  MUX2X1 U119 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n153), .Y(n124) );
  MUX2X1 U120 ( .B(n123), .A(n120), .S(n164), .Y(n134) );
  MUX2X1 U121 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n153), .Y(n128) );
  MUX2X1 U122 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n153), .Y(n127) );
  MUX2X1 U123 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n153), .Y(n131) );
  MUX2X1 U124 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n153), .Y(n130) );
  MUX2X1 U125 ( .B(n129), .A(n126), .S(n164), .Y(n133) );
  MUX2X1 U126 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n153), .Y(n137) );
  MUX2X1 U127 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n153), .Y(n136) );
  MUX2X1 U128 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n153), .Y(n140) );
  MUX2X1 U129 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n153), .Y(n139) );
  MUX2X1 U130 ( .B(n138), .A(n135), .S(n164), .Y(n149) );
  MUX2X1 U131 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n153), .Y(n143) );
  MUX2X1 U132 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n153), .Y(n142) );
  MUX2X1 U133 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n153), .Y(n146) );
  MUX2X1 U134 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n153), .Y(n145) );
  MUX2X1 U135 ( .B(n144), .A(n141), .S(n164), .Y(n148) );
  MUX2X1 U136 ( .B(n147), .A(n132), .S(n168), .Y(n150) );
  INVX8 U137 ( .A(n152), .Y(n153) );
  INVX1 U138 ( .A(n177), .Y(n154) );
  INVX1 U139 ( .A(N10), .Y(n161) );
  AND2X2 U140 ( .A(\data_in<0> ), .B(n154), .Y(n158) );
  INVX8 U141 ( .A(n158), .Y(n179) );
  NAND3X1 U142 ( .A(n168), .B(n166), .C(n10), .Y(n177) );
  OAI21X1 U143 ( .A(n155), .B(n118), .C(\mem<31><0> ), .Y(n170) );
  OAI21X1 U144 ( .A(n179), .B(n118), .C(n170), .Y(n61) );
  OAI21X1 U145 ( .A(n114), .B(n155), .C(\mem<30><0> ), .Y(n171) );
  OAI21X1 U146 ( .A(n114), .B(n179), .C(n171), .Y(n62) );
  NAND3X1 U147 ( .A(n160), .B(n164), .C(n163), .Y(n199) );
  OAI21X1 U148 ( .A(n105), .B(n155), .C(\mem<29><0> ), .Y(n172) );
  OAI21X1 U149 ( .A(n105), .B(n179), .C(n172), .Y(n63) );
  NAND3X1 U150 ( .A(n164), .B(n163), .C(n161), .Y(n201) );
  OAI21X1 U151 ( .A(n107), .B(n155), .C(\mem<28><0> ), .Y(n173) );
  OAI21X1 U152 ( .A(n107), .B(n179), .C(n173), .Y(n64) );
  NAND3X1 U153 ( .A(n160), .B(n162), .C(n165), .Y(n203) );
  OAI21X1 U154 ( .A(n109), .B(n155), .C(\mem<27><0> ), .Y(n174) );
  OAI21X1 U155 ( .A(n109), .B(n179), .C(n174), .Y(n65) );
  NAND3X1 U156 ( .A(n165), .B(n162), .C(n161), .Y(n205) );
  OAI21X1 U157 ( .A(n111), .B(n155), .C(\mem<26><0> ), .Y(n175) );
  OAI21X1 U158 ( .A(n111), .B(n179), .C(n175), .Y(n66) );
  NAND3X1 U159 ( .A(n160), .B(n165), .C(n163), .Y(n207) );
  OAI21X1 U160 ( .A(n113), .B(n155), .C(\mem<25><0> ), .Y(n176) );
  OAI21X1 U161 ( .A(n113), .B(n179), .C(n176), .Y(n67) );
  OAI21X1 U162 ( .A(n116), .B(n155), .C(\mem<24><0> ), .Y(n178) );
  OAI21X1 U163 ( .A(n116), .B(n179), .C(n178), .Y(n68) );
  OAI21X1 U164 ( .A(n187), .B(n118), .C(\mem<23><0> ), .Y(n180) );
  NAND2X1 U165 ( .A(n12), .B(n180), .Y(n69) );
  OAI21X1 U166 ( .A(n187), .B(n114), .C(\mem<22><0> ), .Y(n181) );
  NAND2X1 U167 ( .A(n14), .B(n181), .Y(n70) );
  OAI21X1 U168 ( .A(n187), .B(n105), .C(\mem<21><0> ), .Y(n182) );
  NAND2X1 U169 ( .A(n16), .B(n182), .Y(n71) );
  OAI21X1 U170 ( .A(n187), .B(n107), .C(\mem<20><0> ), .Y(n183) );
  NAND2X1 U171 ( .A(n18), .B(n183), .Y(n72) );
  OAI21X1 U172 ( .A(n187), .B(n109), .C(\mem<19><0> ), .Y(n184) );
  NAND2X1 U173 ( .A(n20), .B(n184), .Y(n73) );
  OAI21X1 U174 ( .A(n187), .B(n111), .C(\mem<18><0> ), .Y(n185) );
  NAND2X1 U175 ( .A(n22), .B(n185), .Y(n74) );
  OAI21X1 U176 ( .A(n187), .B(n113), .C(\mem<17><0> ), .Y(n186) );
  NAND2X1 U177 ( .A(n24), .B(n186), .Y(n75) );
  OAI21X1 U178 ( .A(n187), .B(n116), .C(\mem<16><0> ), .Y(n188) );
  NAND2X1 U179 ( .A(n26), .B(n188), .Y(n76) );
  OAI21X1 U180 ( .A(n157), .B(n118), .C(\mem<15><0> ), .Y(n189) );
  NAND2X1 U181 ( .A(n28), .B(n189), .Y(n77) );
  OAI21X1 U182 ( .A(n157), .B(n114), .C(\mem<14><0> ), .Y(n190) );
  NAND2X1 U183 ( .A(n30), .B(n190), .Y(n78) );
  OAI21X1 U184 ( .A(n157), .B(n105), .C(\mem<13><0> ), .Y(n191) );
  NAND2X1 U185 ( .A(n32), .B(n191), .Y(n79) );
  OAI21X1 U186 ( .A(n157), .B(n107), .C(\mem<12><0> ), .Y(n192) );
  NAND2X1 U187 ( .A(n34), .B(n192), .Y(n80) );
  OAI21X1 U188 ( .A(n157), .B(n109), .C(\mem<11><0> ), .Y(n193) );
  NAND2X1 U189 ( .A(n36), .B(n193), .Y(n81) );
  OAI21X1 U190 ( .A(n157), .B(n111), .C(\mem<10><0> ), .Y(n194) );
  NAND2X1 U191 ( .A(n38), .B(n194), .Y(n82) );
  OAI21X1 U192 ( .A(n157), .B(n113), .C(\mem<9><0> ), .Y(n195) );
  NAND2X1 U193 ( .A(n40), .B(n195), .Y(n83) );
  OAI21X1 U194 ( .A(n157), .B(n116), .C(\mem<8><0> ), .Y(n196) );
  NAND2X1 U195 ( .A(n42), .B(n196), .Y(n84) );
  OAI21X1 U196 ( .A(n156), .B(n118), .C(\mem<7><0> ), .Y(n197) );
  NAND2X1 U197 ( .A(n44), .B(n197), .Y(n85) );
  OAI21X1 U198 ( .A(n156), .B(n114), .C(\mem<6><0> ), .Y(n198) );
  NAND2X1 U199 ( .A(n46), .B(n198), .Y(n86) );
  OAI21X1 U200 ( .A(n156), .B(n105), .C(\mem<5><0> ), .Y(n200) );
  NAND2X1 U201 ( .A(n48), .B(n200), .Y(n87) );
  OAI21X1 U202 ( .A(n156), .B(n107), .C(\mem<4><0> ), .Y(n202) );
  NAND2X1 U203 ( .A(n50), .B(n202), .Y(n88) );
  OAI21X1 U204 ( .A(n156), .B(n109), .C(\mem<3><0> ), .Y(n204) );
  NAND2X1 U205 ( .A(n52), .B(n204), .Y(n89) );
  OAI21X1 U206 ( .A(n156), .B(n111), .C(\mem<2><0> ), .Y(n206) );
  NAND2X1 U207 ( .A(n54), .B(n206), .Y(n90) );
  OAI21X1 U208 ( .A(n156), .B(n113), .C(\mem<1><0> ), .Y(n208) );
  NAND2X1 U209 ( .A(n56), .B(n208), .Y(n91) );
  OAI21X1 U210 ( .A(n156), .B(n116), .C(\mem<0><0> ), .Y(n209) );
  NAND2X1 U211 ( .A(n58), .B(n209), .Y(n92) );
endmodule


module memv_1 ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , N28, n39, n42, n46, n49, n52, n55, n58, n61, n64, n67,
         n70, n73, n76, n79, n82, n85, n88, n90, n91, n92, n94, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n113, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n132, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n151, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n188, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n206, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n224,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n243, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n261, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n279, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n297, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n316, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n334, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n352, n355, n356, n357, n358, n359, n361, n363, n364, n365,
         n366, n367, n368, n370, n371, n372, n373, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n43,
         n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60, n62, n63,
         n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81, n83, n84,
         n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149, n150,
         n152, n169, n171, n187, n189, n205, n207, n223, n225, n241, n242,
         n244, n260, n262, n278, n280, n296, n298, n314, n315, n317, n333,
         n335, n351, n353, n354, n360, n362, n369, n374, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n633), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n632), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n631), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n630), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n629), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n628), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n627), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n626), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n625), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n624), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n623), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n622), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n621), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n620), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n619), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n618), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n617), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n616), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n615), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n614), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n613), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n612), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n611), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n610), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n609), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n608), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n607), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n606), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n605), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n604), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n603), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n602), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n601), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n600), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n599), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n598), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n597), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n596), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n595), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n594), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n593), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n592), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n591), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n590), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n589), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n588), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n587), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n586), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n585), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n584), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n583), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n582), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n581), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n580), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n579), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n578), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n577), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n576), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n575), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n574), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n573), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n572), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n571), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n570), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n569), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n568), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n567), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n566), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n565), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n564), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n563), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n562), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n561), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n560), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n559), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n558), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n557), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n556), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n555), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n554), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n553), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n552), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n551), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n550), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n549), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n548), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n547), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n546), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n545), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n544), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n543), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n542), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n541), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n540), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n539), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n538), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n537), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n536), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n535), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n534), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n533), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n532), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n531), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n530), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n529), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n528), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n527), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n526), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n525), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n524), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n523), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n522), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n521), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n520), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n519), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n518), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n517), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n516), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n515), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n514), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n513), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n512), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n511), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n510), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n509), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n508), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n507), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n506), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n505), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n504), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n503), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n502), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n501), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n500), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n499), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n498), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n497), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n496), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n495), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n494), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n493), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n492), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n491), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n490), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n489), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n488), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n487), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n486), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n485), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n484), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n483), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n482), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n481), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n480), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n479), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n478), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n477), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n476), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n475), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n474), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n473), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n472), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n471), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n470), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n469), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n468), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n467), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n466), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n465), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n464), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n463), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n462), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n461), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n460), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n459), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n458), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n457), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n456), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n455), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n454), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n453), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n452), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n451), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n450), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n449), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n448), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n447), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n446), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n445), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n444), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n443), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n442), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n441), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n440), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n439), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n438), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n437), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n436), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n435), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n434), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n433), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n432), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n431), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n430), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n429), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n428), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n427), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n426), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n425), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n424), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n423), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n422), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n421), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n420), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n419), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n418), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n417), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n416), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n415), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n414), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n413), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n412), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n411), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n410), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n409), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n408), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n407), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n406), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n405), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n404), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n403), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n402), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n401), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n400), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n399), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n398), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n397), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n396), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n395), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n394), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n393), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n392), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n391), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n390), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n389), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n388), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n387), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n386), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n385), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n384), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n383), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n382), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n381), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n380), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n379), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n378), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U5 ( .A(N23), .B(n998), .Y(n111) );
  AND2X2 U6 ( .A(N21), .B(n995), .Y(n355) );
  AND2X2 U7 ( .A(N21), .B(n996), .Y(n364) );
  AND2X2 U8 ( .A(n993), .B(n926), .Y(n356) );
  AND2X2 U9 ( .A(n993), .B(n992), .Y(n358) );
  OAI21X1 U49 ( .A(n962), .B(n991), .C(n42), .Y(n378) );
  OAI21X1 U50 ( .A(n45), .B(n989), .C(\mem<255> ), .Y(n42) );
  OAI21X1 U51 ( .A(n641), .B(n959), .C(n46), .Y(n379) );
  OAI21X1 U52 ( .A(n990), .B(n43), .C(\mem<254> ), .Y(n46) );
  OAI21X1 U53 ( .A(n991), .B(n958), .C(n49), .Y(n380) );
  OAI21X1 U54 ( .A(n990), .B(n40), .C(\mem<253> ), .Y(n49) );
  OAI21X1 U55 ( .A(n641), .B(n957), .C(n52), .Y(n381) );
  OAI21X1 U56 ( .A(n990), .B(n37), .C(\mem<252> ), .Y(n52) );
  OAI21X1 U57 ( .A(n641), .B(n955), .C(n55), .Y(n382) );
  OAI21X1 U58 ( .A(n990), .B(n35), .C(\mem<251> ), .Y(n55) );
  OAI21X1 U59 ( .A(n641), .B(n953), .C(n58), .Y(n383) );
  OAI21X1 U60 ( .A(n990), .B(n33), .C(\mem<250> ), .Y(n58) );
  OAI21X1 U61 ( .A(n641), .B(n951), .C(n61), .Y(n384) );
  OAI21X1 U62 ( .A(n990), .B(n31), .C(\mem<249> ), .Y(n61) );
  OAI21X1 U63 ( .A(n641), .B(n949), .C(n64), .Y(n385) );
  OAI21X1 U64 ( .A(n990), .B(n29), .C(\mem<248> ), .Y(n64) );
  OAI21X1 U65 ( .A(n991), .B(n948), .C(n67), .Y(n386) );
  OAI21X1 U66 ( .A(n990), .B(n27), .C(\mem<247> ), .Y(n67) );
  OAI21X1 U67 ( .A(n991), .B(n947), .C(n70), .Y(n387) );
  OAI21X1 U68 ( .A(n989), .B(n25), .C(\mem<246> ), .Y(n70) );
  OAI21X1 U69 ( .A(n991), .B(n946), .C(n73), .Y(n388) );
  OAI21X1 U70 ( .A(n989), .B(n23), .C(\mem<245> ), .Y(n73) );
  OAI21X1 U71 ( .A(n991), .B(n945), .C(n76), .Y(n389) );
  OAI21X1 U72 ( .A(n989), .B(n21), .C(\mem<244> ), .Y(n76) );
  OAI21X1 U73 ( .A(n991), .B(n944), .C(n79), .Y(n390) );
  OAI21X1 U74 ( .A(n989), .B(n19), .C(\mem<243> ), .Y(n79) );
  OAI21X1 U75 ( .A(n991), .B(n943), .C(n82), .Y(n391) );
  OAI21X1 U76 ( .A(n989), .B(n17), .C(\mem<242> ), .Y(n82) );
  OAI21X1 U77 ( .A(n991), .B(n942), .C(n85), .Y(n392) );
  OAI21X1 U78 ( .A(n989), .B(n15), .C(\mem<241> ), .Y(n85) );
  OAI21X1 U79 ( .A(n991), .B(n939), .C(n88), .Y(n393) );
  OAI21X1 U80 ( .A(n989), .B(n13), .C(\mem<240> ), .Y(n88) );
  OAI21X1 U83 ( .A(n962), .B(n637), .C(n94), .Y(n394) );
  OAI21X1 U84 ( .A(n45), .B(n988), .C(\mem<239> ), .Y(n94) );
  OAI21X1 U85 ( .A(n960), .B(n637), .C(n96), .Y(n395) );
  OAI21X1 U86 ( .A(n43), .B(n988), .C(\mem<238> ), .Y(n96) );
  OAI21X1 U87 ( .A(n958), .B(n637), .C(n97), .Y(n396) );
  OAI21X1 U88 ( .A(n40), .B(n988), .C(\mem<237> ), .Y(n97) );
  OAI21X1 U89 ( .A(n957), .B(n637), .C(n98), .Y(n397) );
  OAI21X1 U90 ( .A(n37), .B(n988), .C(\mem<236> ), .Y(n98) );
  OAI21X1 U91 ( .A(n956), .B(n637), .C(n99), .Y(n398) );
  OAI21X1 U92 ( .A(n35), .B(n988), .C(\mem<235> ), .Y(n99) );
  OAI21X1 U93 ( .A(n954), .B(n637), .C(n100), .Y(n399) );
  OAI21X1 U94 ( .A(n33), .B(n988), .C(\mem<234> ), .Y(n100) );
  OAI21X1 U95 ( .A(n952), .B(n637), .C(n101), .Y(n400) );
  OAI21X1 U96 ( .A(n31), .B(n988), .C(\mem<233> ), .Y(n101) );
  OAI21X1 U97 ( .A(n950), .B(n637), .C(n102), .Y(n401) );
  OAI21X1 U98 ( .A(n29), .B(n988), .C(\mem<232> ), .Y(n102) );
  OAI21X1 U99 ( .A(n948), .B(n637), .C(n103), .Y(n402) );
  OAI21X1 U100 ( .A(n27), .B(n987), .C(\mem<231> ), .Y(n103) );
  OAI21X1 U101 ( .A(n947), .B(n637), .C(n104), .Y(n403) );
  OAI21X1 U102 ( .A(n25), .B(n987), .C(\mem<230> ), .Y(n104) );
  OAI21X1 U103 ( .A(n946), .B(n637), .C(n105), .Y(n404) );
  OAI21X1 U104 ( .A(n23), .B(n987), .C(\mem<229> ), .Y(n105) );
  OAI21X1 U105 ( .A(n945), .B(n637), .C(n106), .Y(n405) );
  OAI21X1 U106 ( .A(n21), .B(n987), .C(\mem<228> ), .Y(n106) );
  OAI21X1 U107 ( .A(n944), .B(n637), .C(n107), .Y(n406) );
  OAI21X1 U108 ( .A(n19), .B(n987), .C(\mem<227> ), .Y(n107) );
  OAI21X1 U109 ( .A(n943), .B(n637), .C(n108), .Y(n407) );
  OAI21X1 U110 ( .A(n17), .B(n987), .C(\mem<226> ), .Y(n108) );
  OAI21X1 U111 ( .A(n942), .B(n637), .C(n109), .Y(n408) );
  OAI21X1 U112 ( .A(n15), .B(n987), .C(\mem<225> ), .Y(n109) );
  OAI21X1 U113 ( .A(n939), .B(n637), .C(n110), .Y(n409) );
  OAI21X1 U114 ( .A(n13), .B(n987), .C(\mem<224> ), .Y(n110) );
  OAI21X1 U117 ( .A(n962), .B(n374), .C(n113), .Y(n410) );
  OAI21X1 U118 ( .A(n45), .B(n986), .C(\mem<223> ), .Y(n113) );
  OAI21X1 U119 ( .A(n960), .B(n374), .C(n115), .Y(n411) );
  OAI21X1 U120 ( .A(n43), .B(n986), .C(\mem<222> ), .Y(n115) );
  OAI21X1 U121 ( .A(n958), .B(n374), .C(n116), .Y(n412) );
  OAI21X1 U122 ( .A(n40), .B(n986), .C(\mem<221> ), .Y(n116) );
  OAI21X1 U123 ( .A(n957), .B(n374), .C(n117), .Y(n413) );
  OAI21X1 U124 ( .A(n37), .B(n986), .C(\mem<220> ), .Y(n117) );
  OAI21X1 U125 ( .A(n956), .B(n374), .C(n118), .Y(n414) );
  OAI21X1 U126 ( .A(n35), .B(n986), .C(\mem<219> ), .Y(n118) );
  OAI21X1 U127 ( .A(n954), .B(n374), .C(n119), .Y(n415) );
  OAI21X1 U128 ( .A(n33), .B(n986), .C(\mem<218> ), .Y(n119) );
  OAI21X1 U129 ( .A(n952), .B(n374), .C(n120), .Y(n416) );
  OAI21X1 U130 ( .A(n31), .B(n986), .C(\mem<217> ), .Y(n120) );
  OAI21X1 U131 ( .A(n950), .B(n374), .C(n121), .Y(n417) );
  OAI21X1 U132 ( .A(n29), .B(n986), .C(\mem<216> ), .Y(n121) );
  OAI21X1 U133 ( .A(n948), .B(n374), .C(n122), .Y(n418) );
  OAI21X1 U134 ( .A(n27), .B(n986), .C(\mem<215> ), .Y(n122) );
  OAI21X1 U135 ( .A(n947), .B(n374), .C(n123), .Y(n419) );
  OAI21X1 U136 ( .A(n25), .B(n986), .C(\mem<214> ), .Y(n123) );
  OAI21X1 U137 ( .A(n946), .B(n374), .C(n124), .Y(n420) );
  OAI21X1 U138 ( .A(n23), .B(n986), .C(\mem<213> ), .Y(n124) );
  OAI21X1 U139 ( .A(n945), .B(n374), .C(n125), .Y(n421) );
  OAI21X1 U140 ( .A(n21), .B(n986), .C(\mem<212> ), .Y(n125) );
  OAI21X1 U141 ( .A(n944), .B(n374), .C(n126), .Y(n422) );
  OAI21X1 U142 ( .A(n19), .B(n986), .C(\mem<211> ), .Y(n126) );
  OAI21X1 U143 ( .A(n943), .B(n374), .C(n127), .Y(n423) );
  OAI21X1 U144 ( .A(n17), .B(n986), .C(\mem<210> ), .Y(n127) );
  OAI21X1 U145 ( .A(n942), .B(n374), .C(n128), .Y(n424) );
  OAI21X1 U146 ( .A(n15), .B(n986), .C(\mem<209> ), .Y(n128) );
  OAI21X1 U147 ( .A(n939), .B(n374), .C(n129), .Y(n425) );
  OAI21X1 U148 ( .A(n13), .B(n986), .C(\mem<208> ), .Y(n129) );
  OAI21X1 U151 ( .A(n962), .B(n362), .C(n132), .Y(n426) );
  OAI21X1 U152 ( .A(n45), .B(n985), .C(\mem<207> ), .Y(n132) );
  OAI21X1 U153 ( .A(n960), .B(n362), .C(n134), .Y(n427) );
  OAI21X1 U154 ( .A(n43), .B(n985), .C(\mem<206> ), .Y(n134) );
  OAI21X1 U155 ( .A(n958), .B(n362), .C(n135), .Y(n428) );
  OAI21X1 U156 ( .A(n40), .B(n985), .C(\mem<205> ), .Y(n135) );
  OAI21X1 U157 ( .A(n957), .B(n362), .C(n136), .Y(n429) );
  OAI21X1 U158 ( .A(n37), .B(n985), .C(\mem<204> ), .Y(n136) );
  OAI21X1 U159 ( .A(n956), .B(n362), .C(n137), .Y(n430) );
  OAI21X1 U160 ( .A(n35), .B(n985), .C(\mem<203> ), .Y(n137) );
  OAI21X1 U161 ( .A(n954), .B(n362), .C(n138), .Y(n431) );
  OAI21X1 U162 ( .A(n33), .B(n985), .C(\mem<202> ), .Y(n138) );
  OAI21X1 U163 ( .A(n952), .B(n362), .C(n139), .Y(n432) );
  OAI21X1 U164 ( .A(n31), .B(n985), .C(\mem<201> ), .Y(n139) );
  OAI21X1 U165 ( .A(n950), .B(n362), .C(n140), .Y(n433) );
  OAI21X1 U166 ( .A(n29), .B(n985), .C(\mem<200> ), .Y(n140) );
  OAI21X1 U167 ( .A(n948), .B(n362), .C(n141), .Y(n434) );
  OAI21X1 U168 ( .A(n27), .B(n985), .C(\mem<199> ), .Y(n141) );
  OAI21X1 U169 ( .A(n947), .B(n362), .C(n142), .Y(n435) );
  OAI21X1 U170 ( .A(n25), .B(n985), .C(\mem<198> ), .Y(n142) );
  OAI21X1 U171 ( .A(n946), .B(n362), .C(n143), .Y(n436) );
  OAI21X1 U172 ( .A(n23), .B(n985), .C(\mem<197> ), .Y(n143) );
  OAI21X1 U173 ( .A(n945), .B(n362), .C(n144), .Y(n437) );
  OAI21X1 U174 ( .A(n21), .B(n985), .C(\mem<196> ), .Y(n144) );
  OAI21X1 U175 ( .A(n944), .B(n362), .C(n145), .Y(n438) );
  OAI21X1 U176 ( .A(n19), .B(n985), .C(\mem<195> ), .Y(n145) );
  OAI21X1 U177 ( .A(n943), .B(n362), .C(n146), .Y(n439) );
  OAI21X1 U178 ( .A(n17), .B(n985), .C(\mem<194> ), .Y(n146) );
  OAI21X1 U179 ( .A(n942), .B(n362), .C(n147), .Y(n440) );
  OAI21X1 U180 ( .A(n15), .B(n985), .C(\mem<193> ), .Y(n147) );
  OAI21X1 U181 ( .A(n939), .B(n362), .C(n148), .Y(n441) );
  OAI21X1 U182 ( .A(n13), .B(n985), .C(\mem<192> ), .Y(n148) );
  OAI21X1 U185 ( .A(n962), .B(n354), .C(n151), .Y(n442) );
  OAI21X1 U186 ( .A(n45), .B(n984), .C(\mem<191> ), .Y(n151) );
  OAI21X1 U187 ( .A(n960), .B(n354), .C(n153), .Y(n443) );
  OAI21X1 U188 ( .A(n43), .B(n984), .C(\mem<190> ), .Y(n153) );
  OAI21X1 U189 ( .A(n958), .B(n354), .C(n154), .Y(n444) );
  OAI21X1 U190 ( .A(n40), .B(n984), .C(\mem<189> ), .Y(n154) );
  OAI21X1 U191 ( .A(n957), .B(n354), .C(n155), .Y(n445) );
  OAI21X1 U192 ( .A(n37), .B(n984), .C(\mem<188> ), .Y(n155) );
  OAI21X1 U193 ( .A(n956), .B(n354), .C(n156), .Y(n446) );
  OAI21X1 U194 ( .A(n35), .B(n984), .C(\mem<187> ), .Y(n156) );
  OAI21X1 U195 ( .A(n954), .B(n354), .C(n157), .Y(n447) );
  OAI21X1 U196 ( .A(n33), .B(n984), .C(\mem<186> ), .Y(n157) );
  OAI21X1 U197 ( .A(n952), .B(n354), .C(n158), .Y(n448) );
  OAI21X1 U198 ( .A(n31), .B(n984), .C(\mem<185> ), .Y(n158) );
  OAI21X1 U199 ( .A(n950), .B(n354), .C(n159), .Y(n449) );
  OAI21X1 U200 ( .A(n29), .B(n984), .C(\mem<184> ), .Y(n159) );
  OAI21X1 U201 ( .A(n948), .B(n354), .C(n160), .Y(n450) );
  OAI21X1 U202 ( .A(n27), .B(n983), .C(\mem<183> ), .Y(n160) );
  OAI21X1 U203 ( .A(n947), .B(n354), .C(n161), .Y(n451) );
  OAI21X1 U204 ( .A(n25), .B(n983), .C(\mem<182> ), .Y(n161) );
  OAI21X1 U205 ( .A(n946), .B(n354), .C(n162), .Y(n452) );
  OAI21X1 U206 ( .A(n23), .B(n983), .C(\mem<181> ), .Y(n162) );
  OAI21X1 U207 ( .A(n945), .B(n354), .C(n163), .Y(n453) );
  OAI21X1 U208 ( .A(n21), .B(n983), .C(\mem<180> ), .Y(n163) );
  OAI21X1 U209 ( .A(n944), .B(n354), .C(n164), .Y(n454) );
  OAI21X1 U210 ( .A(n19), .B(n983), .C(\mem<179> ), .Y(n164) );
  OAI21X1 U211 ( .A(n943), .B(n354), .C(n165), .Y(n455) );
  OAI21X1 U212 ( .A(n17), .B(n983), .C(\mem<178> ), .Y(n165) );
  OAI21X1 U213 ( .A(n942), .B(n354), .C(n166), .Y(n456) );
  OAI21X1 U214 ( .A(n15), .B(n983), .C(\mem<177> ), .Y(n166) );
  OAI21X1 U215 ( .A(n939), .B(n354), .C(n167), .Y(n457) );
  OAI21X1 U216 ( .A(n13), .B(n983), .C(\mem<176> ), .Y(n167) );
  OAI21X1 U219 ( .A(n962), .B(n333), .C(n170), .Y(n458) );
  OAI21X1 U220 ( .A(n45), .B(n982), .C(\mem<175> ), .Y(n170) );
  OAI21X1 U221 ( .A(n960), .B(n333), .C(n172), .Y(n459) );
  OAI21X1 U222 ( .A(n43), .B(n982), .C(\mem<174> ), .Y(n172) );
  OAI21X1 U223 ( .A(n958), .B(n333), .C(n173), .Y(n460) );
  OAI21X1 U224 ( .A(n40), .B(n982), .C(\mem<173> ), .Y(n173) );
  OAI21X1 U225 ( .A(n957), .B(n333), .C(n174), .Y(n461) );
  OAI21X1 U226 ( .A(n37), .B(n982), .C(\mem<172> ), .Y(n174) );
  OAI21X1 U227 ( .A(n956), .B(n333), .C(n175), .Y(n462) );
  OAI21X1 U228 ( .A(n35), .B(n982), .C(\mem<171> ), .Y(n175) );
  OAI21X1 U229 ( .A(n954), .B(n333), .C(n176), .Y(n463) );
  OAI21X1 U230 ( .A(n33), .B(n982), .C(\mem<170> ), .Y(n176) );
  OAI21X1 U231 ( .A(n952), .B(n333), .C(n177), .Y(n464) );
  OAI21X1 U232 ( .A(n31), .B(n982), .C(\mem<169> ), .Y(n177) );
  OAI21X1 U233 ( .A(n950), .B(n333), .C(n178), .Y(n465) );
  OAI21X1 U234 ( .A(n29), .B(n982), .C(\mem<168> ), .Y(n178) );
  OAI21X1 U235 ( .A(n948), .B(n333), .C(n179), .Y(n466) );
  OAI21X1 U236 ( .A(n27), .B(n981), .C(\mem<167> ), .Y(n179) );
  OAI21X1 U237 ( .A(n947), .B(n333), .C(n180), .Y(n467) );
  OAI21X1 U238 ( .A(n25), .B(n981), .C(\mem<166> ), .Y(n180) );
  OAI21X1 U239 ( .A(n946), .B(n333), .C(n181), .Y(n468) );
  OAI21X1 U240 ( .A(n23), .B(n981), .C(\mem<165> ), .Y(n181) );
  OAI21X1 U241 ( .A(n945), .B(n333), .C(n182), .Y(n469) );
  OAI21X1 U242 ( .A(n21), .B(n981), .C(\mem<164> ), .Y(n182) );
  OAI21X1 U243 ( .A(n944), .B(n333), .C(n183), .Y(n470) );
  OAI21X1 U244 ( .A(n19), .B(n981), .C(\mem<163> ), .Y(n183) );
  OAI21X1 U245 ( .A(n943), .B(n333), .C(n184), .Y(n471) );
  OAI21X1 U246 ( .A(n17), .B(n981), .C(\mem<162> ), .Y(n184) );
  OAI21X1 U247 ( .A(n942), .B(n333), .C(n185), .Y(n472) );
  OAI21X1 U248 ( .A(n15), .B(n981), .C(\mem<161> ), .Y(n185) );
  OAI21X1 U249 ( .A(n939), .B(n333), .C(n186), .Y(n473) );
  OAI21X1 U250 ( .A(n13), .B(n981), .C(\mem<160> ), .Y(n186) );
  OAI21X1 U253 ( .A(n962), .B(n298), .C(n188), .Y(n474) );
  OAI21X1 U254 ( .A(n45), .B(n980), .C(\mem<159> ), .Y(n188) );
  OAI21X1 U255 ( .A(n960), .B(n298), .C(n190), .Y(n475) );
  OAI21X1 U256 ( .A(n43), .B(n980), .C(\mem<158> ), .Y(n190) );
  OAI21X1 U257 ( .A(n958), .B(n298), .C(n191), .Y(n476) );
  OAI21X1 U258 ( .A(n40), .B(n980), .C(\mem<157> ), .Y(n191) );
  OAI21X1 U259 ( .A(n957), .B(n298), .C(n192), .Y(n477) );
  OAI21X1 U260 ( .A(n37), .B(n980), .C(\mem<156> ), .Y(n192) );
  OAI21X1 U261 ( .A(n956), .B(n298), .C(n193), .Y(n478) );
  OAI21X1 U262 ( .A(n35), .B(n980), .C(\mem<155> ), .Y(n193) );
  OAI21X1 U263 ( .A(n954), .B(n298), .C(n194), .Y(n479) );
  OAI21X1 U264 ( .A(n33), .B(n980), .C(\mem<154> ), .Y(n194) );
  OAI21X1 U265 ( .A(n952), .B(n298), .C(n195), .Y(n480) );
  OAI21X1 U266 ( .A(n31), .B(n980), .C(\mem<153> ), .Y(n195) );
  OAI21X1 U267 ( .A(n950), .B(n298), .C(n196), .Y(n481) );
  OAI21X1 U268 ( .A(n29), .B(n980), .C(\mem<152> ), .Y(n196) );
  OAI21X1 U269 ( .A(n948), .B(n298), .C(n197), .Y(n482) );
  OAI21X1 U270 ( .A(n27), .B(n979), .C(\mem<151> ), .Y(n197) );
  OAI21X1 U271 ( .A(n947), .B(n298), .C(n198), .Y(n483) );
  OAI21X1 U272 ( .A(n25), .B(n979), .C(\mem<150> ), .Y(n198) );
  OAI21X1 U273 ( .A(n946), .B(n298), .C(n199), .Y(n484) );
  OAI21X1 U274 ( .A(n23), .B(n979), .C(\mem<149> ), .Y(n199) );
  OAI21X1 U275 ( .A(n945), .B(n298), .C(n200), .Y(n485) );
  OAI21X1 U276 ( .A(n21), .B(n979), .C(\mem<148> ), .Y(n200) );
  OAI21X1 U277 ( .A(n944), .B(n298), .C(n201), .Y(n486) );
  OAI21X1 U278 ( .A(n19), .B(n979), .C(\mem<147> ), .Y(n201) );
  OAI21X1 U279 ( .A(n943), .B(n298), .C(n202), .Y(n487) );
  OAI21X1 U280 ( .A(n17), .B(n979), .C(\mem<146> ), .Y(n202) );
  OAI21X1 U281 ( .A(n942), .B(n298), .C(n203), .Y(n488) );
  OAI21X1 U282 ( .A(n15), .B(n979), .C(\mem<145> ), .Y(n203) );
  OAI21X1 U283 ( .A(n939), .B(n298), .C(n204), .Y(n489) );
  OAI21X1 U284 ( .A(n13), .B(n979), .C(\mem<144> ), .Y(n204) );
  OAI21X1 U287 ( .A(n962), .B(n262), .C(n206), .Y(n490) );
  OAI21X1 U288 ( .A(n45), .B(n978), .C(\mem<143> ), .Y(n206) );
  OAI21X1 U289 ( .A(n960), .B(n262), .C(n208), .Y(n491) );
  OAI21X1 U290 ( .A(n43), .B(n978), .C(\mem<142> ), .Y(n208) );
  OAI21X1 U291 ( .A(n958), .B(n262), .C(n209), .Y(n492) );
  OAI21X1 U292 ( .A(n40), .B(n978), .C(\mem<141> ), .Y(n209) );
  OAI21X1 U293 ( .A(n957), .B(n262), .C(n210), .Y(n493) );
  OAI21X1 U294 ( .A(n37), .B(n978), .C(\mem<140> ), .Y(n210) );
  OAI21X1 U295 ( .A(n956), .B(n262), .C(n211), .Y(n494) );
  OAI21X1 U296 ( .A(n35), .B(n978), .C(\mem<139> ), .Y(n211) );
  OAI21X1 U297 ( .A(n954), .B(n262), .C(n212), .Y(n495) );
  OAI21X1 U298 ( .A(n33), .B(n978), .C(\mem<138> ), .Y(n212) );
  OAI21X1 U299 ( .A(n952), .B(n262), .C(n213), .Y(n496) );
  OAI21X1 U300 ( .A(n31), .B(n978), .C(\mem<137> ), .Y(n213) );
  OAI21X1 U301 ( .A(n950), .B(n262), .C(n214), .Y(n497) );
  OAI21X1 U302 ( .A(n29), .B(n978), .C(\mem<136> ), .Y(n214) );
  OAI21X1 U303 ( .A(n948), .B(n262), .C(n215), .Y(n498) );
  OAI21X1 U304 ( .A(n27), .B(n977), .C(\mem<135> ), .Y(n215) );
  OAI21X1 U305 ( .A(n947), .B(n262), .C(n216), .Y(n499) );
  OAI21X1 U306 ( .A(n25), .B(n977), .C(\mem<134> ), .Y(n216) );
  OAI21X1 U307 ( .A(n946), .B(n262), .C(n217), .Y(n500) );
  OAI21X1 U308 ( .A(n23), .B(n977), .C(\mem<133> ), .Y(n217) );
  OAI21X1 U309 ( .A(n945), .B(n262), .C(n218), .Y(n501) );
  OAI21X1 U310 ( .A(n21), .B(n977), .C(\mem<132> ), .Y(n218) );
  OAI21X1 U311 ( .A(n944), .B(n262), .C(n219), .Y(n502) );
  OAI21X1 U312 ( .A(n19), .B(n977), .C(\mem<131> ), .Y(n219) );
  OAI21X1 U313 ( .A(n943), .B(n262), .C(n220), .Y(n503) );
  OAI21X1 U314 ( .A(n17), .B(n977), .C(\mem<130> ), .Y(n220) );
  OAI21X1 U315 ( .A(n942), .B(n262), .C(n221), .Y(n504) );
  OAI21X1 U316 ( .A(n15), .B(n977), .C(\mem<129> ), .Y(n221) );
  OAI21X1 U317 ( .A(n939), .B(n262), .C(n222), .Y(n505) );
  OAI21X1 U318 ( .A(n13), .B(n977), .C(\mem<128> ), .Y(n222) );
  OAI21X1 U321 ( .A(n961), .B(n241), .C(n224), .Y(n506) );
  OAI21X1 U322 ( .A(n45), .B(n975), .C(\mem<127> ), .Y(n224) );
  OAI21X1 U323 ( .A(n960), .B(n241), .C(n226), .Y(n507) );
  OAI21X1 U324 ( .A(n43), .B(n975), .C(\mem<126> ), .Y(n226) );
  OAI21X1 U325 ( .A(n958), .B(n976), .C(n227), .Y(n508) );
  OAI21X1 U326 ( .A(n40), .B(n975), .C(\mem<125> ), .Y(n227) );
  OAI21X1 U327 ( .A(n957), .B(n976), .C(n228), .Y(n509) );
  OAI21X1 U328 ( .A(n37), .B(n975), .C(\mem<124> ), .Y(n228) );
  OAI21X1 U329 ( .A(n956), .B(n241), .C(n229), .Y(n510) );
  OAI21X1 U330 ( .A(n35), .B(n975), .C(\mem<123> ), .Y(n229) );
  OAI21X1 U331 ( .A(n954), .B(n241), .C(n230), .Y(n511) );
  OAI21X1 U332 ( .A(n33), .B(n975), .C(\mem<122> ), .Y(n230) );
  OAI21X1 U333 ( .A(n952), .B(n241), .C(n231), .Y(n512) );
  OAI21X1 U334 ( .A(n31), .B(n975), .C(\mem<121> ), .Y(n231) );
  OAI21X1 U335 ( .A(n950), .B(n241), .C(n232), .Y(n513) );
  OAI21X1 U336 ( .A(n29), .B(n975), .C(\mem<120> ), .Y(n232) );
  OAI21X1 U337 ( .A(n948), .B(n976), .C(n233), .Y(n514) );
  OAI21X1 U338 ( .A(n27), .B(n975), .C(\mem<119> ), .Y(n233) );
  OAI21X1 U339 ( .A(n947), .B(n976), .C(n234), .Y(n515) );
  OAI21X1 U340 ( .A(n25), .B(n975), .C(\mem<118> ), .Y(n234) );
  OAI21X1 U341 ( .A(n946), .B(n976), .C(n235), .Y(n516) );
  OAI21X1 U342 ( .A(n23), .B(n975), .C(\mem<117> ), .Y(n235) );
  OAI21X1 U343 ( .A(n945), .B(n976), .C(n236), .Y(n517) );
  OAI21X1 U344 ( .A(n21), .B(n975), .C(\mem<116> ), .Y(n236) );
  OAI21X1 U345 ( .A(n944), .B(n976), .C(n237), .Y(n518) );
  OAI21X1 U346 ( .A(n19), .B(n975), .C(\mem<115> ), .Y(n237) );
  OAI21X1 U347 ( .A(n943), .B(n976), .C(n238), .Y(n519) );
  OAI21X1 U348 ( .A(n17), .B(n975), .C(\mem<114> ), .Y(n238) );
  OAI21X1 U349 ( .A(n942), .B(n976), .C(n239), .Y(n520) );
  OAI21X1 U350 ( .A(n15), .B(n975), .C(\mem<113> ), .Y(n239) );
  OAI21X1 U351 ( .A(n939), .B(n976), .C(n240), .Y(n521) );
  OAI21X1 U352 ( .A(n13), .B(n975), .C(\mem<112> ), .Y(n240) );
  OAI21X1 U355 ( .A(n961), .B(n223), .C(n243), .Y(n522) );
  OAI21X1 U356 ( .A(n45), .B(n973), .C(\mem<111> ), .Y(n243) );
  OAI21X1 U357 ( .A(n959), .B(n223), .C(n245), .Y(n523) );
  OAI21X1 U358 ( .A(n43), .B(n973), .C(\mem<110> ), .Y(n245) );
  OAI21X1 U359 ( .A(n958), .B(n974), .C(n246), .Y(n524) );
  OAI21X1 U360 ( .A(n40), .B(n973), .C(\mem<109> ), .Y(n246) );
  OAI21X1 U361 ( .A(n957), .B(n974), .C(n247), .Y(n525) );
  OAI21X1 U362 ( .A(n37), .B(n973), .C(\mem<108> ), .Y(n247) );
  OAI21X1 U363 ( .A(n955), .B(n223), .C(n248), .Y(n526) );
  OAI21X1 U364 ( .A(n35), .B(n973), .C(\mem<107> ), .Y(n248) );
  OAI21X1 U365 ( .A(n953), .B(n223), .C(n249), .Y(n527) );
  OAI21X1 U366 ( .A(n33), .B(n973), .C(\mem<106> ), .Y(n249) );
  OAI21X1 U367 ( .A(n951), .B(n223), .C(n250), .Y(n528) );
  OAI21X1 U368 ( .A(n31), .B(n973), .C(\mem<105> ), .Y(n250) );
  OAI21X1 U369 ( .A(n949), .B(n223), .C(n251), .Y(n529) );
  OAI21X1 U370 ( .A(n29), .B(n973), .C(\mem<104> ), .Y(n251) );
  OAI21X1 U371 ( .A(n948), .B(n974), .C(n252), .Y(n530) );
  OAI21X1 U372 ( .A(n27), .B(n973), .C(\mem<103> ), .Y(n252) );
  OAI21X1 U373 ( .A(n947), .B(n974), .C(n253), .Y(n531) );
  OAI21X1 U374 ( .A(n25), .B(n973), .C(\mem<102> ), .Y(n253) );
  OAI21X1 U375 ( .A(n946), .B(n974), .C(n254), .Y(n532) );
  OAI21X1 U376 ( .A(n23), .B(n973), .C(\mem<101> ), .Y(n254) );
  OAI21X1 U377 ( .A(n945), .B(n974), .C(n255), .Y(n533) );
  OAI21X1 U378 ( .A(n21), .B(n973), .C(\mem<100> ), .Y(n255) );
  OAI21X1 U379 ( .A(n944), .B(n974), .C(n256), .Y(n534) );
  OAI21X1 U380 ( .A(n19), .B(n973), .C(\mem<99> ), .Y(n256) );
  OAI21X1 U381 ( .A(n943), .B(n974), .C(n257), .Y(n535) );
  OAI21X1 U382 ( .A(n17), .B(n973), .C(\mem<98> ), .Y(n257) );
  OAI21X1 U383 ( .A(n942), .B(n974), .C(n258), .Y(n536) );
  OAI21X1 U384 ( .A(n15), .B(n973), .C(\mem<97> ), .Y(n258) );
  OAI21X1 U385 ( .A(n939), .B(n974), .C(n259), .Y(n537) );
  OAI21X1 U386 ( .A(n13), .B(n973), .C(\mem<96> ), .Y(n259) );
  OAI21X1 U389 ( .A(n961), .B(n205), .C(n261), .Y(n538) );
  OAI21X1 U390 ( .A(n45), .B(n971), .C(\mem<95> ), .Y(n261) );
  OAI21X1 U391 ( .A(n959), .B(n205), .C(n263), .Y(n539) );
  OAI21X1 U392 ( .A(n43), .B(n971), .C(\mem<94> ), .Y(n263) );
  OAI21X1 U393 ( .A(n958), .B(n972), .C(n264), .Y(n540) );
  OAI21X1 U394 ( .A(n40), .B(n971), .C(\mem<93> ), .Y(n264) );
  OAI21X1 U395 ( .A(n957), .B(n972), .C(n265), .Y(n541) );
  OAI21X1 U396 ( .A(n37), .B(n971), .C(\mem<92> ), .Y(n265) );
  OAI21X1 U397 ( .A(n955), .B(n205), .C(n266), .Y(n542) );
  OAI21X1 U398 ( .A(n35), .B(n971), .C(\mem<91> ), .Y(n266) );
  OAI21X1 U399 ( .A(n953), .B(n205), .C(n267), .Y(n543) );
  OAI21X1 U400 ( .A(n33), .B(n971), .C(\mem<90> ), .Y(n267) );
  OAI21X1 U401 ( .A(n951), .B(n205), .C(n268), .Y(n544) );
  OAI21X1 U402 ( .A(n31), .B(n971), .C(\mem<89> ), .Y(n268) );
  OAI21X1 U403 ( .A(n949), .B(n205), .C(n269), .Y(n545) );
  OAI21X1 U404 ( .A(n29), .B(n971), .C(\mem<88> ), .Y(n269) );
  OAI21X1 U405 ( .A(n948), .B(n972), .C(n270), .Y(n546) );
  OAI21X1 U406 ( .A(n27), .B(n971), .C(\mem<87> ), .Y(n270) );
  OAI21X1 U407 ( .A(n947), .B(n972), .C(n271), .Y(n547) );
  OAI21X1 U408 ( .A(n25), .B(n971), .C(\mem<86> ), .Y(n271) );
  OAI21X1 U409 ( .A(n946), .B(n972), .C(n272), .Y(n548) );
  OAI21X1 U410 ( .A(n23), .B(n971), .C(\mem<85> ), .Y(n272) );
  OAI21X1 U411 ( .A(n945), .B(n972), .C(n273), .Y(n549) );
  OAI21X1 U412 ( .A(n21), .B(n971), .C(\mem<84> ), .Y(n273) );
  OAI21X1 U413 ( .A(n944), .B(n972), .C(n274), .Y(n550) );
  OAI21X1 U414 ( .A(n19), .B(n971), .C(\mem<83> ), .Y(n274) );
  OAI21X1 U415 ( .A(n943), .B(n972), .C(n275), .Y(n551) );
  OAI21X1 U416 ( .A(n17), .B(n971), .C(\mem<82> ), .Y(n275) );
  OAI21X1 U417 ( .A(n942), .B(n972), .C(n276), .Y(n552) );
  OAI21X1 U418 ( .A(n15), .B(n971), .C(\mem<81> ), .Y(n276) );
  OAI21X1 U419 ( .A(n939), .B(n972), .C(n277), .Y(n553) );
  OAI21X1 U420 ( .A(n13), .B(n971), .C(\mem<80> ), .Y(n277) );
  OAI21X1 U423 ( .A(n961), .B(n187), .C(n279), .Y(n554) );
  OAI21X1 U424 ( .A(n45), .B(n969), .C(\mem<79> ), .Y(n279) );
  OAI21X1 U425 ( .A(n959), .B(n187), .C(n281), .Y(n555) );
  OAI21X1 U426 ( .A(n43), .B(n969), .C(\mem<78> ), .Y(n281) );
  OAI21X1 U427 ( .A(n958), .B(n970), .C(n282), .Y(n556) );
  OAI21X1 U428 ( .A(n40), .B(n969), .C(\mem<77> ), .Y(n282) );
  OAI21X1 U429 ( .A(n957), .B(n970), .C(n283), .Y(n557) );
  OAI21X1 U430 ( .A(n37), .B(n969), .C(\mem<76> ), .Y(n283) );
  OAI21X1 U431 ( .A(n955), .B(n187), .C(n284), .Y(n558) );
  OAI21X1 U432 ( .A(n35), .B(n969), .C(\mem<75> ), .Y(n284) );
  OAI21X1 U433 ( .A(n953), .B(n187), .C(n285), .Y(n559) );
  OAI21X1 U434 ( .A(n33), .B(n969), .C(\mem<74> ), .Y(n285) );
  OAI21X1 U435 ( .A(n951), .B(n187), .C(n286), .Y(n560) );
  OAI21X1 U436 ( .A(n31), .B(n969), .C(\mem<73> ), .Y(n286) );
  OAI21X1 U437 ( .A(n949), .B(n187), .C(n287), .Y(n561) );
  OAI21X1 U438 ( .A(n29), .B(n969), .C(\mem<72> ), .Y(n287) );
  OAI21X1 U439 ( .A(n948), .B(n970), .C(n288), .Y(n562) );
  OAI21X1 U440 ( .A(n27), .B(n969), .C(\mem<71> ), .Y(n288) );
  OAI21X1 U441 ( .A(n947), .B(n970), .C(n289), .Y(n563) );
  OAI21X1 U442 ( .A(n25), .B(n969), .C(\mem<70> ), .Y(n289) );
  OAI21X1 U443 ( .A(n946), .B(n970), .C(n290), .Y(n564) );
  OAI21X1 U444 ( .A(n23), .B(n969), .C(\mem<69> ), .Y(n290) );
  OAI21X1 U445 ( .A(n945), .B(n970), .C(n291), .Y(n565) );
  OAI21X1 U446 ( .A(n21), .B(n969), .C(\mem<68> ), .Y(n291) );
  OAI21X1 U447 ( .A(n944), .B(n970), .C(n292), .Y(n566) );
  OAI21X1 U448 ( .A(n19), .B(n969), .C(\mem<67> ), .Y(n292) );
  OAI21X1 U449 ( .A(n943), .B(n970), .C(n293), .Y(n567) );
  OAI21X1 U450 ( .A(n17), .B(n969), .C(\mem<66> ), .Y(n293) );
  OAI21X1 U451 ( .A(n942), .B(n970), .C(n294), .Y(n568) );
  OAI21X1 U452 ( .A(n15), .B(n969), .C(\mem<65> ), .Y(n294) );
  OAI21X1 U453 ( .A(n939), .B(n970), .C(n295), .Y(n569) );
  OAI21X1 U454 ( .A(n13), .B(n969), .C(\mem<64> ), .Y(n295) );
  OAI21X1 U458 ( .A(n961), .B(n169), .C(n297), .Y(n570) );
  OAI21X1 U459 ( .A(n45), .B(n967), .C(\mem<63> ), .Y(n297) );
  OAI21X1 U460 ( .A(n959), .B(n169), .C(n299), .Y(n571) );
  OAI21X1 U461 ( .A(n43), .B(n967), .C(\mem<62> ), .Y(n299) );
  OAI21X1 U462 ( .A(n958), .B(n968), .C(n300), .Y(n572) );
  OAI21X1 U463 ( .A(n40), .B(n967), .C(\mem<61> ), .Y(n300) );
  OAI21X1 U464 ( .A(n957), .B(n968), .C(n301), .Y(n573) );
  OAI21X1 U465 ( .A(n37), .B(n967), .C(\mem<60> ), .Y(n301) );
  OAI21X1 U466 ( .A(n955), .B(n169), .C(n302), .Y(n574) );
  OAI21X1 U467 ( .A(n35), .B(n967), .C(\mem<59> ), .Y(n302) );
  OAI21X1 U468 ( .A(n953), .B(n169), .C(n303), .Y(n575) );
  OAI21X1 U469 ( .A(n33), .B(n967), .C(\mem<58> ), .Y(n303) );
  OAI21X1 U470 ( .A(n951), .B(n169), .C(n304), .Y(n576) );
  OAI21X1 U471 ( .A(n31), .B(n967), .C(\mem<57> ), .Y(n304) );
  OAI21X1 U472 ( .A(n949), .B(n169), .C(n305), .Y(n577) );
  OAI21X1 U473 ( .A(n29), .B(n967), .C(\mem<56> ), .Y(n305) );
  OAI21X1 U474 ( .A(n948), .B(n968), .C(n306), .Y(n578) );
  OAI21X1 U475 ( .A(n27), .B(n967), .C(\mem<55> ), .Y(n306) );
  OAI21X1 U476 ( .A(n947), .B(n968), .C(n307), .Y(n579) );
  OAI21X1 U477 ( .A(n25), .B(n967), .C(\mem<54> ), .Y(n307) );
  OAI21X1 U478 ( .A(n946), .B(n968), .C(n308), .Y(n580) );
  OAI21X1 U479 ( .A(n23), .B(n967), .C(\mem<53> ), .Y(n308) );
  OAI21X1 U480 ( .A(n945), .B(n968), .C(n309), .Y(n581) );
  OAI21X1 U481 ( .A(n21), .B(n967), .C(\mem<52> ), .Y(n309) );
  OAI21X1 U482 ( .A(n944), .B(n968), .C(n310), .Y(n582) );
  OAI21X1 U483 ( .A(n19), .B(n967), .C(\mem<51> ), .Y(n310) );
  OAI21X1 U484 ( .A(n943), .B(n968), .C(n311), .Y(n583) );
  OAI21X1 U485 ( .A(n17), .B(n967), .C(\mem<50> ), .Y(n311) );
  OAI21X1 U486 ( .A(n942), .B(n968), .C(n312), .Y(n584) );
  OAI21X1 U487 ( .A(n15), .B(n967), .C(\mem<49> ), .Y(n312) );
  OAI21X1 U488 ( .A(n939), .B(n968), .C(n313), .Y(n585) );
  OAI21X1 U489 ( .A(n13), .B(n967), .C(\mem<48> ), .Y(n313) );
  OAI21X1 U492 ( .A(n961), .B(n150), .C(n316), .Y(n586) );
  OAI21X1 U493 ( .A(n45), .B(n965), .C(\mem<47> ), .Y(n316) );
  OAI21X1 U494 ( .A(n959), .B(n150), .C(n318), .Y(n587) );
  OAI21X1 U495 ( .A(n43), .B(n965), .C(\mem<46> ), .Y(n318) );
  OAI21X1 U496 ( .A(n958), .B(n966), .C(n319), .Y(n588) );
  OAI21X1 U497 ( .A(n40), .B(n965), .C(\mem<45> ), .Y(n319) );
  OAI21X1 U498 ( .A(n957), .B(n966), .C(n320), .Y(n589) );
  OAI21X1 U499 ( .A(n37), .B(n965), .C(\mem<44> ), .Y(n320) );
  OAI21X1 U500 ( .A(n955), .B(n150), .C(n321), .Y(n590) );
  OAI21X1 U501 ( .A(n35), .B(n965), .C(\mem<43> ), .Y(n321) );
  OAI21X1 U502 ( .A(n953), .B(n150), .C(n322), .Y(n591) );
  OAI21X1 U503 ( .A(n33), .B(n965), .C(\mem<42> ), .Y(n322) );
  OAI21X1 U504 ( .A(n951), .B(n150), .C(n323), .Y(n592) );
  OAI21X1 U505 ( .A(n31), .B(n965), .C(\mem<41> ), .Y(n323) );
  OAI21X1 U506 ( .A(n949), .B(n150), .C(n324), .Y(n593) );
  OAI21X1 U507 ( .A(n29), .B(n965), .C(\mem<40> ), .Y(n324) );
  OAI21X1 U508 ( .A(n948), .B(n966), .C(n325), .Y(n594) );
  OAI21X1 U509 ( .A(n27), .B(n965), .C(\mem<39> ), .Y(n325) );
  OAI21X1 U510 ( .A(n947), .B(n966), .C(n326), .Y(n595) );
  OAI21X1 U511 ( .A(n25), .B(n965), .C(\mem<38> ), .Y(n326) );
  OAI21X1 U512 ( .A(n946), .B(n966), .C(n327), .Y(n596) );
  OAI21X1 U513 ( .A(n23), .B(n965), .C(\mem<37> ), .Y(n327) );
  OAI21X1 U514 ( .A(n945), .B(n966), .C(n328), .Y(n597) );
  OAI21X1 U515 ( .A(n21), .B(n965), .C(\mem<36> ), .Y(n328) );
  OAI21X1 U516 ( .A(n944), .B(n966), .C(n329), .Y(n598) );
  OAI21X1 U517 ( .A(n19), .B(n965), .C(\mem<35> ), .Y(n329) );
  OAI21X1 U518 ( .A(n943), .B(n966), .C(n330), .Y(n599) );
  OAI21X1 U519 ( .A(n17), .B(n965), .C(\mem<34> ), .Y(n330) );
  OAI21X1 U520 ( .A(n942), .B(n966), .C(n331), .Y(n600) );
  OAI21X1 U521 ( .A(n15), .B(n965), .C(\mem<33> ), .Y(n331) );
  OAI21X1 U522 ( .A(n939), .B(n966), .C(n332), .Y(n601) );
  OAI21X1 U523 ( .A(n13), .B(n965), .C(\mem<32> ), .Y(n332) );
  OAI21X1 U526 ( .A(n961), .B(n133), .C(n334), .Y(n602) );
  OAI21X1 U527 ( .A(n45), .B(n963), .C(\mem<31> ), .Y(n334) );
  OAI21X1 U528 ( .A(n959), .B(n133), .C(n336), .Y(n603) );
  OAI21X1 U529 ( .A(n43), .B(n963), .C(\mem<30> ), .Y(n336) );
  OAI21X1 U530 ( .A(n958), .B(n964), .C(n337), .Y(n604) );
  OAI21X1 U531 ( .A(n40), .B(n963), .C(\mem<29> ), .Y(n337) );
  OAI21X1 U532 ( .A(n957), .B(n964), .C(n338), .Y(n605) );
  OAI21X1 U533 ( .A(n37), .B(n963), .C(\mem<28> ), .Y(n338) );
  OAI21X1 U534 ( .A(n955), .B(n133), .C(n339), .Y(n606) );
  OAI21X1 U535 ( .A(n35), .B(n963), .C(\mem<27> ), .Y(n339) );
  OAI21X1 U536 ( .A(n953), .B(n133), .C(n340), .Y(n607) );
  OAI21X1 U537 ( .A(n33), .B(n963), .C(\mem<26> ), .Y(n340) );
  OAI21X1 U538 ( .A(n951), .B(n133), .C(n341), .Y(n608) );
  OAI21X1 U539 ( .A(n31), .B(n963), .C(\mem<25> ), .Y(n341) );
  OAI21X1 U540 ( .A(n949), .B(n133), .C(n342), .Y(n609) );
  OAI21X1 U541 ( .A(n29), .B(n963), .C(\mem<24> ), .Y(n342) );
  OAI21X1 U542 ( .A(n948), .B(n964), .C(n343), .Y(n610) );
  OAI21X1 U543 ( .A(n27), .B(n963), .C(\mem<23> ), .Y(n343) );
  OAI21X1 U544 ( .A(n947), .B(n964), .C(n344), .Y(n611) );
  OAI21X1 U545 ( .A(n25), .B(n963), .C(\mem<22> ), .Y(n344) );
  OAI21X1 U546 ( .A(n946), .B(n964), .C(n345), .Y(n612) );
  OAI21X1 U547 ( .A(n23), .B(n963), .C(\mem<21> ), .Y(n345) );
  OAI21X1 U548 ( .A(n945), .B(n964), .C(n346), .Y(n613) );
  OAI21X1 U549 ( .A(n21), .B(n963), .C(\mem<20> ), .Y(n346) );
  OAI21X1 U550 ( .A(n944), .B(n964), .C(n347), .Y(n614) );
  OAI21X1 U551 ( .A(n19), .B(n963), .C(\mem<19> ), .Y(n347) );
  OAI21X1 U552 ( .A(n943), .B(n964), .C(n348), .Y(n615) );
  OAI21X1 U553 ( .A(n17), .B(n963), .C(\mem<18> ), .Y(n348) );
  OAI21X1 U554 ( .A(n942), .B(n964), .C(n349), .Y(n616) );
  OAI21X1 U555 ( .A(n15), .B(n963), .C(\mem<17> ), .Y(n349) );
  OAI21X1 U556 ( .A(n939), .B(n964), .C(n350), .Y(n617) );
  OAI21X1 U557 ( .A(n13), .B(n963), .C(\mem<16> ), .Y(n350) );
  OAI21X1 U561 ( .A(n961), .B(n78), .C(n352), .Y(n618) );
  OAI21X1 U562 ( .A(n45), .B(n940), .C(\mem<15> ), .Y(n352) );
  OAI21X1 U565 ( .A(n959), .B(n78), .C(n357), .Y(n619) );
  OAI21X1 U566 ( .A(n43), .B(n940), .C(\mem<14> ), .Y(n357) );
  OAI21X1 U569 ( .A(n958), .B(n941), .C(n359), .Y(n620) );
  OAI21X1 U570 ( .A(n40), .B(n940), .C(\mem<13> ), .Y(n359) );
  OAI21X1 U573 ( .A(n957), .B(n941), .C(n361), .Y(n621) );
  OAI21X1 U574 ( .A(n37), .B(n940), .C(\mem<12> ), .Y(n361) );
  OAI21X1 U577 ( .A(n955), .B(n78), .C(n363), .Y(n622) );
  OAI21X1 U578 ( .A(n35), .B(n940), .C(\mem<11> ), .Y(n363) );
  OAI21X1 U581 ( .A(n953), .B(n78), .C(n365), .Y(n623) );
  OAI21X1 U582 ( .A(n33), .B(n940), .C(\mem<10> ), .Y(n365) );
  OAI21X1 U585 ( .A(n951), .B(n78), .C(n366), .Y(n624) );
  OAI21X1 U586 ( .A(n31), .B(n940), .C(\mem<9> ), .Y(n366) );
  OAI21X1 U589 ( .A(n949), .B(n78), .C(n367), .Y(n625) );
  OAI21X1 U590 ( .A(n29), .B(n940), .C(\mem<8> ), .Y(n367) );
  OAI21X1 U593 ( .A(n948), .B(n941), .C(n368), .Y(n626) );
  OAI21X1 U594 ( .A(n27), .B(n940), .C(\mem<7> ), .Y(n368) );
  OAI21X1 U597 ( .A(n947), .B(n941), .C(n370), .Y(n627) );
  OAI21X1 U598 ( .A(n25), .B(n940), .C(\mem<6> ), .Y(n370) );
  OAI21X1 U601 ( .A(n946), .B(n941), .C(n371), .Y(n628) );
  OAI21X1 U602 ( .A(n23), .B(n940), .C(\mem<5> ), .Y(n371) );
  OAI21X1 U605 ( .A(n945), .B(n941), .C(n372), .Y(n629) );
  OAI21X1 U606 ( .A(n21), .B(n940), .C(\mem<4> ), .Y(n372) );
  OAI21X1 U610 ( .A(n944), .B(n941), .C(n373), .Y(n630) );
  OAI21X1 U611 ( .A(n19), .B(n940), .C(\mem<3> ), .Y(n373) );
  OAI21X1 U614 ( .A(n943), .B(n941), .C(n375), .Y(n631) );
  OAI21X1 U615 ( .A(n17), .B(n940), .C(\mem<2> ), .Y(n375) );
  OAI21X1 U618 ( .A(n942), .B(n941), .C(n376), .Y(n632) );
  OAI21X1 U619 ( .A(n15), .B(n940), .C(\mem<1> ), .Y(n376) );
  OAI21X1 U623 ( .A(n939), .B(n941), .C(n377), .Y(n633) );
  OAI21X1 U624 ( .A(n13), .B(n940), .C(\mem<0> ), .Y(n377) );
  BUFX4 U2 ( .A(n641), .Y(n991) );
  BUFX4 U3 ( .A(n223), .Y(n974) );
  BUFX4 U4 ( .A(n205), .Y(n972) );
  BUFX4 U10 ( .A(n187), .Y(n970) );
  BUFX4 U11 ( .A(n169), .Y(n968) );
  BUFX4 U12 ( .A(n150), .Y(n966) );
  BUFX4 U13 ( .A(n133), .Y(n964) );
  BUFX4 U14 ( .A(n78), .Y(n941) );
  INVX2 U15 ( .A(n636), .Y(n637) );
  INVX2 U16 ( .A(n369), .Y(n374) );
  INVX2 U17 ( .A(n360), .Y(n362) );
  INVX2 U18 ( .A(n353), .Y(n354) );
  INVX2 U19 ( .A(n317), .Y(n333) );
  INVX2 U20 ( .A(n296), .Y(n298) );
  INVX2 U21 ( .A(n260), .Y(n262) );
  BUFX4 U22 ( .A(n241), .Y(n976) );
  AND2X1 U23 ( .A(data_in), .B(n4), .Y(n90) );
  AND2X1 U24 ( .A(N25), .B(n999), .Y(n168) );
  AND2X1 U25 ( .A(N25), .B(N24), .Y(n91) );
  AND2X1 U26 ( .A(N23), .B(n997), .Y(n92) );
  INVX1 U27 ( .A(write), .Y(n39) );
  BUFX2 U28 ( .A(n638), .Y(n989) );
  BUFX2 U29 ( .A(n635), .Y(n987) );
  BUFX2 U30 ( .A(n351), .Y(n983) );
  BUFX2 U31 ( .A(n315), .Y(n981) );
  BUFX2 U32 ( .A(n280), .Y(n979) );
  BUFX2 U33 ( .A(n244), .Y(n977) );
  BUFX2 U34 ( .A(n130), .Y(n961) );
  BUFX2 U35 ( .A(n112), .Y(n959) );
  BUFX2 U36 ( .A(n93), .Y(n955) );
  BUFX2 U37 ( .A(n87), .Y(n953) );
  BUFX2 U38 ( .A(n84), .Y(n951) );
  BUFX2 U39 ( .A(n81), .Y(n949) );
  INVX1 U40 ( .A(n48), .Y(n940) );
  INVX1 U41 ( .A(n63), .Y(n963) );
  INVX1 U42 ( .A(n68), .Y(n969) );
  INVX1 U43 ( .A(n69), .Y(n971) );
  INVX1 U44 ( .A(n50), .Y(n942) );
  INVX1 U45 ( .A(n56), .Y(n946) );
  INVX1 U46 ( .A(n74), .Y(n985) );
  INVX1 U47 ( .A(n75), .Y(n986) );
  BUFX2 U48 ( .A(n81), .Y(n950) );
  BUFX2 U81 ( .A(n84), .Y(n952) );
  INVX1 U82 ( .A(n66), .Y(n967) );
  INVX1 U115 ( .A(n72), .Y(n975) );
  INVX1 U116 ( .A(n65), .Y(n965) );
  INVX1 U149 ( .A(n71), .Y(n973) );
  INVX1 U150 ( .A(n53), .Y(n944) );
  INVX1 U183 ( .A(n59), .Y(n948) );
  INVX1 U184 ( .A(n51), .Y(n943) );
  INVX1 U217 ( .A(n57), .Y(n947) );
  BUFX2 U218 ( .A(n87), .Y(n954) );
  BUFX2 U251 ( .A(n112), .Y(n960) );
  BUFX2 U252 ( .A(n130), .Y(n962) );
  INVX1 U285 ( .A(n47), .Y(n939) );
  INVX1 U286 ( .A(n54), .Y(n945) );
  INVX1 U319 ( .A(n60), .Y(n957) );
  INVX1 U320 ( .A(n62), .Y(n958) );
  BUFX2 U353 ( .A(n244), .Y(n978) );
  BUFX2 U354 ( .A(n280), .Y(n980) );
  BUFX2 U387 ( .A(n315), .Y(n982) );
  BUFX2 U388 ( .A(n351), .Y(n984) );
  BUFX2 U421 ( .A(n635), .Y(n988) );
  BUFX2 U422 ( .A(n638), .Y(n990) );
  BUFX2 U455 ( .A(n93), .Y(n956) );
  INVX1 U456 ( .A(n996), .Y(n995) );
  INVX1 U457 ( .A(n998), .Y(n997) );
  INVX2 U490 ( .A(N22), .Y(n998) );
  OR2X2 U491 ( .A(n926), .B(n993), .Y(n1) );
  INVX1 U524 ( .A(n1), .Y(n2) );
  OR2X2 U525 ( .A(n39), .B(rst), .Y(n3) );
  INVX1 U558 ( .A(n3), .Y(n4) );
  AND2X2 U559 ( .A(n9), .B(n7), .Y(n5) );
  AND2X2 U560 ( .A(n690), .B(n914), .Y(n6) );
  INVX1 U563 ( .A(n6), .Y(n7) );
  AND2X2 U564 ( .A(n691), .B(n921), .Y(n8) );
  INVX1 U567 ( .A(n8), .Y(n9) );
  INVX4 U568 ( .A(N18), .Y(n992) );
  MUX2X1 U571 ( .B(\mem<75> ), .A(\mem<74> ), .S(n923), .Y(n829) );
  MUX2X1 U572 ( .B(\mem<87> ), .A(\mem<86> ), .S(n923), .Y(n817) );
  MUX2X1 U575 ( .B(n829), .A(n828), .S(n915), .Y(n827) );
  MUX2X1 U576 ( .B(\mem<21> ), .A(\mem<20> ), .S(n922), .Y(n879) );
  MUX2X1 U579 ( .B(\mem<65> ), .A(\mem<64> ), .S(n923), .Y(n834) );
  MUX2X1 U580 ( .B(\mem<85> ), .A(\mem<84> ), .S(n923), .Y(n816) );
  MUX2X1 U583 ( .B(\mem<69> ), .A(\mem<68> ), .S(n923), .Y(n831) );
  INVX1 U584 ( .A(N28), .Y(n1000) );
  MUX2X1 U587 ( .B(n821), .A(n836), .S(n998), .Y(n840) );
  INVX1 U588 ( .A(n998), .Y(n907) );
  INVX4 U591 ( .A(n992), .Y(n937) );
  OR2X2 U592 ( .A(n992), .B(n993), .Y(n10) );
  INVX1 U595 ( .A(n10), .Y(n11) );
  INVX4 U596 ( .A(n994), .Y(n993) );
  AND2X1 U599 ( .A(n47), .B(n4), .Y(n12) );
  INVX1 U600 ( .A(n12), .Y(n13) );
  AND2X1 U603 ( .A(n50), .B(n4), .Y(n14) );
  INVX1 U604 ( .A(n14), .Y(n15) );
  AND2X1 U607 ( .A(n51), .B(n4), .Y(n16) );
  INVX1 U608 ( .A(n16), .Y(n17) );
  AND2X1 U609 ( .A(n53), .B(n4), .Y(n18) );
  INVX1 U612 ( .A(n18), .Y(n19) );
  AND2X1 U613 ( .A(n54), .B(n4), .Y(n20) );
  INVX1 U616 ( .A(n20), .Y(n21) );
  AND2X1 U617 ( .A(n56), .B(n4), .Y(n22) );
  INVX1 U620 ( .A(n22), .Y(n23) );
  AND2X1 U621 ( .A(n57), .B(n4), .Y(n24) );
  INVX1 U622 ( .A(n24), .Y(n25) );
  AND2X1 U625 ( .A(n59), .B(n4), .Y(n26) );
  INVX1 U626 ( .A(n26), .Y(n27) );
  AND2X1 U627 ( .A(n80), .B(n4), .Y(n28) );
  INVX1 U628 ( .A(n28), .Y(n29) );
  AND2X1 U629 ( .A(n83), .B(n4), .Y(n30) );
  INVX1 U630 ( .A(n30), .Y(n31) );
  AND2X1 U631 ( .A(n86), .B(n4), .Y(n32) );
  INVX1 U632 ( .A(n32), .Y(n33) );
  AND2X1 U633 ( .A(n89), .B(n4), .Y(n34) );
  INVX1 U634 ( .A(n34), .Y(n35) );
  AND2X1 U635 ( .A(n60), .B(n4), .Y(n36) );
  INVX1 U636 ( .A(n36), .Y(n37) );
  AND2X1 U637 ( .A(n62), .B(n4), .Y(n38) );
  INVX1 U638 ( .A(n38), .Y(n40) );
  AND2X1 U639 ( .A(n95), .B(n4), .Y(n41) );
  INVX1 U640 ( .A(n41), .Y(n43) );
  AND2X1 U641 ( .A(n114), .B(n4), .Y(n44) );
  INVX1 U642 ( .A(n44), .Y(n45) );
  AND2X1 U643 ( .A(n647), .B(n2), .Y(n47) );
  AND2X1 U644 ( .A(n649), .B(n643), .Y(n48) );
  AND2X1 U645 ( .A(n647), .B(n11), .Y(n50) );
  AND2X1 U646 ( .A(n647), .B(n358), .Y(n51) );
  AND2X1 U647 ( .A(n647), .B(n356), .Y(n53) );
  AND2X1 U648 ( .A(n651), .B(n2), .Y(n54) );
  AND2X1 U649 ( .A(n651), .B(n11), .Y(n56) );
  AND2X1 U650 ( .A(n651), .B(n358), .Y(n57) );
  AND2X1 U651 ( .A(n651), .B(n356), .Y(n59) );
  AND2X1 U652 ( .A(n2), .B(n355), .Y(n60) );
  AND2X1 U653 ( .A(n11), .B(n355), .Y(n62) );
  AND2X1 U654 ( .A(n649), .B(n645), .Y(n63) );
  AND2X1 U655 ( .A(n649), .B(n111), .Y(n65) );
  AND2X1 U656 ( .A(n649), .B(n92), .Y(n66) );
  AND2X1 U657 ( .A(n653), .B(n643), .Y(n68) );
  AND2X1 U658 ( .A(n653), .B(n645), .Y(n69) );
  AND2X1 U659 ( .A(n653), .B(n111), .Y(n71) );
  AND2X1 U660 ( .A(n653), .B(n92), .Y(n72) );
  AND2X1 U661 ( .A(n643), .B(n91), .Y(n74) );
  AND2X1 U662 ( .A(n645), .B(n91), .Y(n75) );
  AND2X1 U663 ( .A(n48), .B(n90), .Y(n77) );
  INVX1 U664 ( .A(n77), .Y(n78) );
  AND2X1 U665 ( .A(n364), .B(n2), .Y(n80) );
  INVX1 U666 ( .A(n80), .Y(n81) );
  AND2X1 U667 ( .A(n364), .B(n11), .Y(n83) );
  INVX1 U668 ( .A(n83), .Y(n84) );
  AND2X1 U669 ( .A(n364), .B(n358), .Y(n86) );
  INVX1 U670 ( .A(n86), .Y(n87) );
  AND2X1 U671 ( .A(n364), .B(n356), .Y(n89) );
  INVX1 U672 ( .A(n89), .Y(n93) );
  AND2X1 U673 ( .A(n358), .B(n355), .Y(n95) );
  INVX1 U674 ( .A(n95), .Y(n112) );
  AND2X1 U675 ( .A(n355), .B(n356), .Y(n114) );
  INVX1 U676 ( .A(n114), .Y(n130) );
  AND2X1 U677 ( .A(n63), .B(n90), .Y(n131) );
  INVX1 U678 ( .A(n131), .Y(n133) );
  AND2X1 U679 ( .A(n65), .B(n90), .Y(n149) );
  INVX1 U680 ( .A(n149), .Y(n150) );
  AND2X1 U681 ( .A(n66), .B(n90), .Y(n152) );
  INVX1 U682 ( .A(n152), .Y(n169) );
  AND2X1 U683 ( .A(n68), .B(n90), .Y(n171) );
  INVX1 U684 ( .A(n171), .Y(n187) );
  AND2X1 U685 ( .A(n69), .B(n90), .Y(n189) );
  INVX1 U686 ( .A(n189), .Y(n205) );
  AND2X1 U687 ( .A(n71), .B(n90), .Y(n207) );
  INVX1 U688 ( .A(n207), .Y(n223) );
  AND2X1 U689 ( .A(n72), .B(n90), .Y(n225) );
  INVX1 U690 ( .A(n225), .Y(n241) );
  AND2X1 U691 ( .A(n168), .B(n643), .Y(n242) );
  INVX1 U692 ( .A(n242), .Y(n244) );
  AND2X1 U693 ( .A(n242), .B(n90), .Y(n260) );
  AND2X1 U694 ( .A(n168), .B(n645), .Y(n278) );
  INVX1 U695 ( .A(n278), .Y(n280) );
  AND2X1 U696 ( .A(n278), .B(n90), .Y(n296) );
  AND2X1 U697 ( .A(n168), .B(n111), .Y(n314) );
  INVX1 U698 ( .A(n314), .Y(n315) );
  AND2X1 U699 ( .A(n314), .B(n90), .Y(n317) );
  AND2X1 U700 ( .A(n168), .B(n92), .Y(n335) );
  INVX1 U701 ( .A(n335), .Y(n351) );
  AND2X1 U702 ( .A(n335), .B(n90), .Y(n353) );
  AND2X1 U703 ( .A(n74), .B(n90), .Y(n360) );
  AND2X1 U704 ( .A(n75), .B(n90), .Y(n369) );
  AND2X1 U705 ( .A(n111), .B(n91), .Y(n634) );
  INVX1 U706 ( .A(n634), .Y(n635) );
  AND2X1 U707 ( .A(n634), .B(n90), .Y(n636) );
  INVX1 U708 ( .A(n639), .Y(n638) );
  AND2X1 U709 ( .A(n91), .B(n92), .Y(n639) );
  AND2X1 U710 ( .A(n90), .B(n639), .Y(n640) );
  INVX1 U711 ( .A(n640), .Y(n641) );
  OR2X1 U712 ( .A(n997), .B(N23), .Y(n642) );
  INVX1 U713 ( .A(n642), .Y(n643) );
  OR2X1 U714 ( .A(n998), .B(N23), .Y(n644) );
  INVX1 U715 ( .A(n644), .Y(n645) );
  OR2X2 U716 ( .A(n995), .B(N21), .Y(n646) );
  INVX1 U717 ( .A(n646), .Y(n647) );
  OR2X1 U718 ( .A(N24), .B(N25), .Y(n648) );
  INVX1 U719 ( .A(n648), .Y(n649) );
  OR2X2 U720 ( .A(n996), .B(N21), .Y(n650) );
  INVX1 U721 ( .A(n650), .Y(n651) );
  OR2X1 U722 ( .A(n999), .B(N25), .Y(n652) );
  INVX1 U723 ( .A(n652), .Y(n653) );
  MUX2X1 U724 ( .B(n839), .A(n902), .S(n999), .Y(n905) );
  INVX1 U725 ( .A(N24), .Y(n999) );
  MUX2X1 U726 ( .B(n822), .A(n823), .S(n909), .Y(n821) );
  INVX1 U727 ( .A(n908), .Y(n909) );
  INVX1 U728 ( .A(N21), .Y(n908) );
  INVX1 U729 ( .A(N19), .Y(n994) );
  MUX2X1 U730 ( .B(n655), .A(n656), .S(n921), .Y(n654) );
  MUX2X1 U731 ( .B(n658), .A(n659), .S(n921), .Y(n657) );
  MUX2X1 U732 ( .B(n661), .A(n662), .S(n921), .Y(n660) );
  MUX2X1 U733 ( .B(n664), .A(n665), .S(n921), .Y(n663) );
  MUX2X1 U734 ( .B(n667), .A(n668), .S(n910), .Y(n666) );
  MUX2X1 U735 ( .B(n670), .A(n671), .S(n921), .Y(n669) );
  MUX2X1 U736 ( .B(n673), .A(n674), .S(n921), .Y(n672) );
  MUX2X1 U737 ( .B(n676), .A(n677), .S(n921), .Y(n675) );
  MUX2X1 U738 ( .B(n679), .A(n680), .S(n921), .Y(n678) );
  MUX2X1 U739 ( .B(n682), .A(n683), .S(n910), .Y(n681) );
  MUX2X1 U740 ( .B(n685), .A(n686), .S(n921), .Y(n684) );
  MUX2X1 U741 ( .B(n688), .A(n689), .S(n921), .Y(n687) );
  MUX2X1 U742 ( .B(n693), .A(n694), .S(n921), .Y(n692) );
  MUX2X1 U743 ( .B(n696), .A(n697), .S(n910), .Y(n695) );
  MUX2X1 U744 ( .B(n699), .A(n700), .S(n920), .Y(n698) );
  MUX2X1 U745 ( .B(n702), .A(n703), .S(n920), .Y(n701) );
  MUX2X1 U746 ( .B(n705), .A(n706), .S(n920), .Y(n704) );
  MUX2X1 U747 ( .B(n708), .A(n709), .S(n920), .Y(n707) );
  MUX2X1 U748 ( .B(n711), .A(n712), .S(n910), .Y(n710) );
  MUX2X1 U749 ( .B(n714), .A(n715), .S(N23), .Y(n713) );
  MUX2X1 U750 ( .B(n717), .A(n718), .S(n920), .Y(n716) );
  MUX2X1 U751 ( .B(n720), .A(n721), .S(n920), .Y(n719) );
  MUX2X1 U752 ( .B(n723), .A(n724), .S(n920), .Y(n722) );
  MUX2X1 U753 ( .B(n726), .A(n727), .S(n920), .Y(n725) );
  MUX2X1 U754 ( .B(n729), .A(n730), .S(n910), .Y(n728) );
  MUX2X1 U755 ( .B(n732), .A(n733), .S(n920), .Y(n731) );
  MUX2X1 U756 ( .B(n735), .A(n736), .S(n920), .Y(n734) );
  MUX2X1 U757 ( .B(n738), .A(n739), .S(n920), .Y(n737) );
  MUX2X1 U758 ( .B(n741), .A(n742), .S(n920), .Y(n740) );
  MUX2X1 U759 ( .B(n744), .A(n745), .S(n910), .Y(n743) );
  MUX2X1 U760 ( .B(n747), .A(n748), .S(n919), .Y(n746) );
  MUX2X1 U761 ( .B(n750), .A(n751), .S(n919), .Y(n749) );
  MUX2X1 U762 ( .B(n753), .A(n754), .S(n919), .Y(n752) );
  MUX2X1 U763 ( .B(n756), .A(n757), .S(n919), .Y(n755) );
  MUX2X1 U764 ( .B(n759), .A(n760), .S(n910), .Y(n758) );
  MUX2X1 U765 ( .B(n762), .A(n763), .S(n919), .Y(n761) );
  MUX2X1 U766 ( .B(n765), .A(n766), .S(n919), .Y(n764) );
  MUX2X1 U767 ( .B(n768), .A(n769), .S(n919), .Y(n767) );
  MUX2X1 U768 ( .B(n771), .A(n772), .S(n919), .Y(n770) );
  MUX2X1 U769 ( .B(n774), .A(n775), .S(n910), .Y(n773) );
  MUX2X1 U770 ( .B(n777), .A(n778), .S(N23), .Y(n776) );
  MUX2X1 U771 ( .B(n780), .A(n781), .S(n919), .Y(n779) );
  MUX2X1 U772 ( .B(n783), .A(n784), .S(n919), .Y(n782) );
  MUX2X1 U773 ( .B(n786), .A(n787), .S(n919), .Y(n785) );
  MUX2X1 U774 ( .B(n789), .A(n790), .S(n919), .Y(n788) );
  MUX2X1 U775 ( .B(n792), .A(n793), .S(n910), .Y(n791) );
  MUX2X1 U776 ( .B(n795), .A(n796), .S(n918), .Y(n794) );
  MUX2X1 U777 ( .B(n798), .A(n799), .S(n918), .Y(n797) );
  MUX2X1 U778 ( .B(n801), .A(n802), .S(n918), .Y(n800) );
  MUX2X1 U779 ( .B(n804), .A(n805), .S(n918), .Y(n803) );
  MUX2X1 U780 ( .B(n807), .A(n808), .S(n910), .Y(n806) );
  MUX2X1 U781 ( .B(n810), .A(n811), .S(n918), .Y(n809) );
  MUX2X1 U782 ( .B(n813), .A(n814), .S(n918), .Y(n812) );
  MUX2X1 U783 ( .B(n816), .A(n817), .S(n918), .Y(n815) );
  MUX2X1 U784 ( .B(n819), .A(n820), .S(n918), .Y(n818) );
  MUX2X1 U785 ( .B(n825), .A(n826), .S(n918), .Y(n824) );
  MUX2X1 U786 ( .B(n831), .A(n832), .S(n918), .Y(n830) );
  MUX2X1 U787 ( .B(n834), .A(n835), .S(n918), .Y(n833) );
  MUX2X1 U788 ( .B(n837), .A(n838), .S(n910), .Y(n836) );
  MUX2X1 U789 ( .B(n840), .A(n841), .S(N23), .Y(n839) );
  MUX2X1 U790 ( .B(n843), .A(n844), .S(n917), .Y(n842) );
  MUX2X1 U791 ( .B(n846), .A(n847), .S(n917), .Y(n845) );
  MUX2X1 U792 ( .B(n849), .A(n850), .S(n917), .Y(n848) );
  MUX2X1 U793 ( .B(n852), .A(n853), .S(n917), .Y(n851) );
  MUX2X1 U794 ( .B(n855), .A(n856), .S(n909), .Y(n854) );
  MUX2X1 U795 ( .B(n858), .A(n859), .S(n917), .Y(n857) );
  MUX2X1 U796 ( .B(n861), .A(n862), .S(n917), .Y(n860) );
  MUX2X1 U797 ( .B(n864), .A(n865), .S(n917), .Y(n863) );
  MUX2X1 U798 ( .B(n867), .A(n868), .S(n917), .Y(n866) );
  MUX2X1 U799 ( .B(n870), .A(n871), .S(n909), .Y(n869) );
  MUX2X1 U800 ( .B(n873), .A(n874), .S(n917), .Y(n872) );
  MUX2X1 U801 ( .B(n876), .A(n877), .S(n917), .Y(n875) );
  MUX2X1 U802 ( .B(n879), .A(n880), .S(n917), .Y(n878) );
  MUX2X1 U803 ( .B(n882), .A(n883), .S(n917), .Y(n881) );
  MUX2X1 U804 ( .B(n885), .A(n886), .S(n909), .Y(n884) );
  MUX2X1 U805 ( .B(n888), .A(n889), .S(n916), .Y(n887) );
  MUX2X1 U806 ( .B(n891), .A(n892), .S(n916), .Y(n890) );
  MUX2X1 U807 ( .B(n894), .A(n895), .S(n916), .Y(n893) );
  MUX2X1 U808 ( .B(n897), .A(n898), .S(n916), .Y(n896) );
  MUX2X1 U809 ( .B(n900), .A(n901), .S(n909), .Y(n899) );
  MUX2X1 U810 ( .B(n903), .A(n904), .S(N23), .Y(n902) );
  MUX2X1 U811 ( .B(n905), .A(n906), .S(N25), .Y(N28) );
  MUX2X1 U812 ( .B(\mem<254> ), .A(\mem<255> ), .S(n926), .Y(n656) );
  MUX2X1 U813 ( .B(\mem<252> ), .A(\mem<253> ), .S(n926), .Y(n655) );
  MUX2X1 U814 ( .B(\mem<250> ), .A(\mem<251> ), .S(n926), .Y(n659) );
  MUX2X1 U815 ( .B(\mem<248> ), .A(\mem<249> ), .S(n926), .Y(n658) );
  MUX2X1 U816 ( .B(n657), .A(n654), .S(n913), .Y(n668) );
  MUX2X1 U817 ( .B(\mem<246> ), .A(\mem<247> ), .S(n926), .Y(n662) );
  MUX2X1 U818 ( .B(\mem<244> ), .A(\mem<245> ), .S(n926), .Y(n661) );
  MUX2X1 U819 ( .B(\mem<242> ), .A(\mem<243> ), .S(n926), .Y(n665) );
  MUX2X1 U820 ( .B(\mem<240> ), .A(\mem<241> ), .S(n926), .Y(n664) );
  MUX2X1 U821 ( .B(n663), .A(n660), .S(n913), .Y(n667) );
  MUX2X1 U822 ( .B(\mem<238> ), .A(\mem<239> ), .S(n927), .Y(n671) );
  MUX2X1 U823 ( .B(\mem<236> ), .A(\mem<237> ), .S(n927), .Y(n670) );
  MUX2X1 U824 ( .B(\mem<234> ), .A(\mem<235> ), .S(n927), .Y(n674) );
  MUX2X1 U825 ( .B(\mem<232> ), .A(\mem<233> ), .S(n927), .Y(n673) );
  MUX2X1 U826 ( .B(n672), .A(n669), .S(n913), .Y(n683) );
  MUX2X1 U827 ( .B(\mem<230> ), .A(\mem<231> ), .S(n927), .Y(n677) );
  MUX2X1 U828 ( .B(\mem<228> ), .A(\mem<229> ), .S(n927), .Y(n676) );
  MUX2X1 U829 ( .B(\mem<226> ), .A(\mem<227> ), .S(n927), .Y(n680) );
  MUX2X1 U830 ( .B(\mem<224> ), .A(\mem<225> ), .S(n927), .Y(n679) );
  MUX2X1 U831 ( .B(n678), .A(n675), .S(n913), .Y(n682) );
  MUX2X1 U832 ( .B(n681), .A(n666), .S(n907), .Y(n715) );
  MUX2X1 U833 ( .B(\mem<222> ), .A(\mem<223> ), .S(n927), .Y(n686) );
  MUX2X1 U834 ( .B(\mem<220> ), .A(\mem<221> ), .S(n927), .Y(n685) );
  MUX2X1 U835 ( .B(\mem<218> ), .A(\mem<219> ), .S(n927), .Y(n689) );
  MUX2X1 U836 ( .B(\mem<216> ), .A(\mem<217> ), .S(n927), .Y(n688) );
  MUX2X1 U837 ( .B(n687), .A(n684), .S(n913), .Y(n697) );
  MUX2X1 U838 ( .B(\mem<214> ), .A(\mem<215> ), .S(n928), .Y(n691) );
  MUX2X1 U839 ( .B(\mem<212> ), .A(\mem<213> ), .S(n928), .Y(n690) );
  MUX2X1 U840 ( .B(\mem<210> ), .A(\mem<211> ), .S(n928), .Y(n694) );
  MUX2X1 U841 ( .B(\mem<208> ), .A(\mem<209> ), .S(n928), .Y(n693) );
  MUX2X1 U842 ( .B(n692), .A(n5), .S(n913), .Y(n696) );
  MUX2X1 U843 ( .B(\mem<206> ), .A(\mem<207> ), .S(n928), .Y(n700) );
  MUX2X1 U844 ( .B(\mem<204> ), .A(\mem<205> ), .S(n928), .Y(n699) );
  MUX2X1 U845 ( .B(\mem<202> ), .A(\mem<203> ), .S(n928), .Y(n703) );
  MUX2X1 U846 ( .B(\mem<200> ), .A(\mem<201> ), .S(n928), .Y(n702) );
  MUX2X1 U847 ( .B(n701), .A(n698), .S(n913), .Y(n712) );
  MUX2X1 U848 ( .B(\mem<198> ), .A(\mem<199> ), .S(n928), .Y(n706) );
  MUX2X1 U849 ( .B(\mem<196> ), .A(\mem<197> ), .S(n928), .Y(n705) );
  MUX2X1 U850 ( .B(\mem<194> ), .A(\mem<195> ), .S(n928), .Y(n709) );
  MUX2X1 U851 ( .B(\mem<192> ), .A(\mem<193> ), .S(n928), .Y(n708) );
  MUX2X1 U852 ( .B(n707), .A(n704), .S(n913), .Y(n711) );
  MUX2X1 U853 ( .B(n710), .A(n695), .S(n907), .Y(n714) );
  MUX2X1 U854 ( .B(\mem<190> ), .A(\mem<191> ), .S(n929), .Y(n718) );
  MUX2X1 U855 ( .B(\mem<188> ), .A(\mem<189> ), .S(n929), .Y(n717) );
  MUX2X1 U856 ( .B(\mem<186> ), .A(\mem<187> ), .S(n929), .Y(n721) );
  MUX2X1 U857 ( .B(\mem<184> ), .A(\mem<185> ), .S(n929), .Y(n720) );
  MUX2X1 U858 ( .B(n719), .A(n716), .S(n913), .Y(n730) );
  MUX2X1 U859 ( .B(\mem<182> ), .A(\mem<183> ), .S(n929), .Y(n724) );
  MUX2X1 U860 ( .B(\mem<180> ), .A(\mem<181> ), .S(n929), .Y(n723) );
  MUX2X1 U861 ( .B(\mem<178> ), .A(\mem<179> ), .S(n929), .Y(n727) );
  MUX2X1 U862 ( .B(\mem<176> ), .A(\mem<177> ), .S(n929), .Y(n726) );
  MUX2X1 U863 ( .B(n725), .A(n722), .S(n913), .Y(n729) );
  MUX2X1 U864 ( .B(\mem<174> ), .A(\mem<175> ), .S(n929), .Y(n733) );
  MUX2X1 U865 ( .B(\mem<172> ), .A(\mem<173> ), .S(n929), .Y(n732) );
  MUX2X1 U866 ( .B(\mem<170> ), .A(\mem<171> ), .S(n929), .Y(n736) );
  MUX2X1 U867 ( .B(\mem<168> ), .A(\mem<169> ), .S(n929), .Y(n735) );
  MUX2X1 U868 ( .B(n734), .A(n731), .S(n913), .Y(n745) );
  MUX2X1 U869 ( .B(\mem<166> ), .A(\mem<167> ), .S(n930), .Y(n739) );
  MUX2X1 U870 ( .B(\mem<164> ), .A(\mem<165> ), .S(n930), .Y(n738) );
  MUX2X1 U871 ( .B(\mem<162> ), .A(\mem<163> ), .S(n930), .Y(n742) );
  MUX2X1 U872 ( .B(\mem<160> ), .A(\mem<161> ), .S(n930), .Y(n741) );
  MUX2X1 U873 ( .B(n740), .A(n737), .S(n913), .Y(n744) );
  MUX2X1 U874 ( .B(n743), .A(n728), .S(n907), .Y(n778) );
  MUX2X1 U875 ( .B(\mem<158> ), .A(\mem<159> ), .S(n930), .Y(n748) );
  MUX2X1 U876 ( .B(\mem<156> ), .A(\mem<157> ), .S(n930), .Y(n747) );
  MUX2X1 U877 ( .B(\mem<154> ), .A(\mem<155> ), .S(n930), .Y(n751) );
  MUX2X1 U878 ( .B(\mem<152> ), .A(\mem<153> ), .S(n930), .Y(n750) );
  MUX2X1 U879 ( .B(n749), .A(n746), .S(n912), .Y(n760) );
  MUX2X1 U880 ( .B(\mem<150> ), .A(\mem<151> ), .S(n930), .Y(n754) );
  MUX2X1 U881 ( .B(\mem<148> ), .A(\mem<149> ), .S(n930), .Y(n753) );
  MUX2X1 U882 ( .B(\mem<146> ), .A(\mem<147> ), .S(n930), .Y(n757) );
  MUX2X1 U883 ( .B(\mem<144> ), .A(\mem<145> ), .S(n930), .Y(n756) );
  MUX2X1 U884 ( .B(n755), .A(n752), .S(n912), .Y(n759) );
  MUX2X1 U885 ( .B(\mem<142> ), .A(\mem<143> ), .S(n931), .Y(n763) );
  MUX2X1 U886 ( .B(\mem<140> ), .A(\mem<141> ), .S(n931), .Y(n762) );
  MUX2X1 U887 ( .B(\mem<138> ), .A(\mem<139> ), .S(n931), .Y(n766) );
  MUX2X1 U888 ( .B(\mem<136> ), .A(\mem<137> ), .S(n931), .Y(n765) );
  MUX2X1 U889 ( .B(n764), .A(n761), .S(n912), .Y(n775) );
  MUX2X1 U890 ( .B(\mem<134> ), .A(\mem<135> ), .S(n931), .Y(n769) );
  MUX2X1 U891 ( .B(\mem<132> ), .A(\mem<133> ), .S(n931), .Y(n768) );
  MUX2X1 U892 ( .B(\mem<130> ), .A(\mem<131> ), .S(n931), .Y(n772) );
  MUX2X1 U893 ( .B(\mem<128> ), .A(\mem<129> ), .S(n931), .Y(n771) );
  MUX2X1 U894 ( .B(n770), .A(n767), .S(n912), .Y(n774) );
  MUX2X1 U895 ( .B(n773), .A(n758), .S(n907), .Y(n777) );
  MUX2X1 U896 ( .B(n776), .A(n713), .S(N24), .Y(n906) );
  MUX2X1 U897 ( .B(\mem<126> ), .A(\mem<127> ), .S(n931), .Y(n781) );
  MUX2X1 U898 ( .B(\mem<124> ), .A(\mem<125> ), .S(n931), .Y(n780) );
  MUX2X1 U899 ( .B(\mem<122> ), .A(\mem<123> ), .S(n931), .Y(n784) );
  MUX2X1 U900 ( .B(\mem<120> ), .A(\mem<121> ), .S(n931), .Y(n783) );
  MUX2X1 U901 ( .B(n782), .A(n779), .S(n912), .Y(n793) );
  MUX2X1 U902 ( .B(\mem<118> ), .A(\mem<119> ), .S(n932), .Y(n787) );
  MUX2X1 U903 ( .B(\mem<116> ), .A(\mem<117> ), .S(n934), .Y(n786) );
  MUX2X1 U904 ( .B(\mem<114> ), .A(\mem<115> ), .S(n932), .Y(n790) );
  MUX2X1 U905 ( .B(\mem<112> ), .A(\mem<113> ), .S(n934), .Y(n789) );
  MUX2X1 U906 ( .B(n788), .A(n785), .S(n912), .Y(n792) );
  MUX2X1 U907 ( .B(\mem<110> ), .A(\mem<111> ), .S(n933), .Y(n796) );
  MUX2X1 U908 ( .B(\mem<108> ), .A(\mem<109> ), .S(n932), .Y(n795) );
  MUX2X1 U909 ( .B(\mem<106> ), .A(\mem<107> ), .S(n933), .Y(n799) );
  MUX2X1 U910 ( .B(\mem<104> ), .A(\mem<105> ), .S(n932), .Y(n798) );
  MUX2X1 U911 ( .B(n797), .A(n794), .S(n912), .Y(n808) );
  MUX2X1 U912 ( .B(\mem<102> ), .A(\mem<103> ), .S(n933), .Y(n802) );
  MUX2X1 U913 ( .B(\mem<100> ), .A(\mem<101> ), .S(n934), .Y(n801) );
  MUX2X1 U914 ( .B(\mem<98> ), .A(\mem<99> ), .S(n933), .Y(n805) );
  MUX2X1 U915 ( .B(\mem<96> ), .A(\mem<97> ), .S(n933), .Y(n804) );
  MUX2X1 U916 ( .B(n803), .A(n800), .S(n912), .Y(n807) );
  MUX2X1 U917 ( .B(n806), .A(n791), .S(n907), .Y(n841) );
  MUX2X1 U918 ( .B(\mem<94> ), .A(\mem<95> ), .S(n933), .Y(n811) );
  MUX2X1 U919 ( .B(\mem<92> ), .A(\mem<93> ), .S(n932), .Y(n810) );
  MUX2X1 U920 ( .B(\mem<90> ), .A(\mem<91> ), .S(n932), .Y(n814) );
  MUX2X1 U921 ( .B(\mem<88> ), .A(\mem<89> ), .S(n932), .Y(n813) );
  MUX2X1 U922 ( .B(n812), .A(n809), .S(n912), .Y(n823) );
  MUX2X1 U923 ( .B(\mem<82> ), .A(\mem<83> ), .S(n933), .Y(n820) );
  MUX2X1 U924 ( .B(\mem<80> ), .A(\mem<81> ), .S(n934), .Y(n819) );
  MUX2X1 U925 ( .B(n818), .A(n815), .S(n912), .Y(n822) );
  MUX2X1 U926 ( .B(\mem<78> ), .A(\mem<79> ), .S(n933), .Y(n826) );
  MUX2X1 U927 ( .B(\mem<76> ), .A(\mem<77> ), .S(n934), .Y(n825) );
  MUX2X1 U928 ( .B(\mem<72> ), .A(\mem<73> ), .S(n933), .Y(n828) );
  MUX2X1 U929 ( .B(n827), .A(n824), .S(n912), .Y(n838) );
  MUX2X1 U930 ( .B(\mem<70> ), .A(\mem<71> ), .S(n934), .Y(n832) );
  MUX2X1 U931 ( .B(\mem<66> ), .A(\mem<67> ), .S(n932), .Y(n835) );
  MUX2X1 U932 ( .B(n833), .A(n830), .S(n912), .Y(n837) );
  MUX2X1 U933 ( .B(\mem<62> ), .A(\mem<63> ), .S(n933), .Y(n844) );
  MUX2X1 U934 ( .B(\mem<60> ), .A(\mem<61> ), .S(n932), .Y(n843) );
  MUX2X1 U935 ( .B(\mem<58> ), .A(\mem<59> ), .S(n932), .Y(n847) );
  MUX2X1 U936 ( .B(\mem<56> ), .A(\mem<57> ), .S(n933), .Y(n846) );
  MUX2X1 U937 ( .B(n845), .A(n842), .S(n911), .Y(n856) );
  MUX2X1 U938 ( .B(\mem<54> ), .A(\mem<55> ), .S(n933), .Y(n850) );
  MUX2X1 U939 ( .B(\mem<52> ), .A(\mem<53> ), .S(n934), .Y(n849) );
  MUX2X1 U940 ( .B(\mem<50> ), .A(\mem<51> ), .S(n932), .Y(n853) );
  MUX2X1 U941 ( .B(\mem<48> ), .A(\mem<49> ), .S(n934), .Y(n852) );
  MUX2X1 U942 ( .B(n851), .A(n848), .S(n911), .Y(n855) );
  MUX2X1 U943 ( .B(\mem<46> ), .A(\mem<47> ), .S(n935), .Y(n859) );
  MUX2X1 U944 ( .B(\mem<44> ), .A(\mem<45> ), .S(n935), .Y(n858) );
  MUX2X1 U945 ( .B(\mem<42> ), .A(\mem<43> ), .S(n935), .Y(n862) );
  MUX2X1 U946 ( .B(\mem<40> ), .A(\mem<41> ), .S(n935), .Y(n861) );
  MUX2X1 U947 ( .B(n860), .A(n857), .S(n911), .Y(n871) );
  MUX2X1 U948 ( .B(\mem<38> ), .A(\mem<39> ), .S(n935), .Y(n865) );
  MUX2X1 U949 ( .B(\mem<36> ), .A(\mem<37> ), .S(n935), .Y(n864) );
  MUX2X1 U950 ( .B(\mem<34> ), .A(\mem<35> ), .S(n935), .Y(n868) );
  MUX2X1 U951 ( .B(\mem<32> ), .A(\mem<33> ), .S(n935), .Y(n867) );
  MUX2X1 U952 ( .B(n866), .A(n863), .S(n911), .Y(n870) );
  MUX2X1 U953 ( .B(n869), .A(n854), .S(n907), .Y(n904) );
  MUX2X1 U954 ( .B(\mem<30> ), .A(\mem<31> ), .S(n935), .Y(n874) );
  MUX2X1 U955 ( .B(\mem<28> ), .A(\mem<29> ), .S(n935), .Y(n873) );
  MUX2X1 U956 ( .B(\mem<26> ), .A(\mem<27> ), .S(n935), .Y(n877) );
  MUX2X1 U957 ( .B(\mem<24> ), .A(\mem<25> ), .S(n935), .Y(n876) );
  MUX2X1 U958 ( .B(n875), .A(n872), .S(n911), .Y(n886) );
  MUX2X1 U959 ( .B(\mem<22> ), .A(\mem<23> ), .S(n936), .Y(n880) );
  MUX2X1 U960 ( .B(\mem<18> ), .A(\mem<19> ), .S(n936), .Y(n883) );
  MUX2X1 U961 ( .B(\mem<16> ), .A(\mem<17> ), .S(n936), .Y(n882) );
  MUX2X1 U962 ( .B(n881), .A(n878), .S(n911), .Y(n885) );
  MUX2X1 U963 ( .B(\mem<14> ), .A(\mem<15> ), .S(n936), .Y(n889) );
  MUX2X1 U964 ( .B(\mem<12> ), .A(\mem<13> ), .S(n936), .Y(n888) );
  MUX2X1 U965 ( .B(\mem<10> ), .A(\mem<11> ), .S(n936), .Y(n892) );
  MUX2X1 U966 ( .B(\mem<8> ), .A(\mem<9> ), .S(n936), .Y(n891) );
  MUX2X1 U967 ( .B(n890), .A(n887), .S(n911), .Y(n901) );
  MUX2X1 U968 ( .B(\mem<6> ), .A(\mem<7> ), .S(n936), .Y(n895) );
  MUX2X1 U969 ( .B(\mem<4> ), .A(\mem<5> ), .S(n936), .Y(n894) );
  MUX2X1 U970 ( .B(\mem<2> ), .A(\mem<3> ), .S(n936), .Y(n898) );
  MUX2X1 U971 ( .B(\mem<0> ), .A(\mem<1> ), .S(n936), .Y(n897) );
  MUX2X1 U972 ( .B(n896), .A(n893), .S(n911), .Y(n900) );
  MUX2X1 U973 ( .B(n899), .A(n884), .S(n907), .Y(n903) );
  INVX8 U974 ( .A(n908), .Y(n910) );
  INVX8 U975 ( .A(n996), .Y(n911) );
  INVX8 U976 ( .A(n996), .Y(n912) );
  INVX8 U977 ( .A(n996), .Y(n913) );
  INVX8 U978 ( .A(n993), .Y(n914) );
  INVX8 U979 ( .A(n993), .Y(n915) );
  INVX8 U980 ( .A(n915), .Y(n916) );
  INVX8 U981 ( .A(n915), .Y(n917) );
  INVX8 U982 ( .A(n915), .Y(n918) );
  INVX8 U983 ( .A(n914), .Y(n919) );
  INVX8 U984 ( .A(n914), .Y(n920) );
  INVX8 U985 ( .A(n914), .Y(n921) );
  INVX8 U986 ( .A(n937), .Y(n922) );
  INVX8 U987 ( .A(n938), .Y(n923) );
  INVX8 U988 ( .A(n938), .Y(n924) );
  INVX8 U989 ( .A(n938), .Y(n925) );
  INVX8 U990 ( .A(n925), .Y(n926) );
  INVX8 U991 ( .A(n925), .Y(n927) );
  INVX8 U992 ( .A(n925), .Y(n928) );
  INVX8 U993 ( .A(n924), .Y(n929) );
  INVX8 U994 ( .A(n924), .Y(n930) );
  INVX8 U995 ( .A(n924), .Y(n931) );
  INVX8 U996 ( .A(n923), .Y(n932) );
  INVX8 U997 ( .A(n923), .Y(n933) );
  INVX8 U998 ( .A(n923), .Y(n934) );
  INVX8 U999 ( .A(n922), .Y(n935) );
  INVX8 U1000 ( .A(n922), .Y(n936) );
  INVX8 U1001 ( .A(n992), .Y(n938) );
  INVX8 U1002 ( .A(N20), .Y(n996) );
  NOR3X1 U1003 ( .A(write), .B(rst), .C(n1000), .Y(data_out) );
endmodule


module memc_Size16_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2400), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2401), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2402), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2403), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2404), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2405), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2406), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2407), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2408), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2409), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2410), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2411), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2412), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2413), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2414), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2415), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2416), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2417), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2418), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2419), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2420), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2421), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2422), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2423), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2424), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2425), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2426), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2427), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2428), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2429), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2430), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2431), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2432), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2433), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2434), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2435), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2436), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2437), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2438), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2439), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2440), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2441), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2442), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2443), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2444), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2445), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2446), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2447), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2448), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2449), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2450), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2451), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2452), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2453), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2454), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2455), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2456), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2457), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2458), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2459), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2460), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2461), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2462), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2463), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2464), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2465), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2466), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2467), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2468), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2469), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2470), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2471), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2472), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2473), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2474), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2475), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2476), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2477), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2478), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2479), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2480), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2481), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2482), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2483), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2484), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2485), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2486), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2487), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2488), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2489), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2490), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2491), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2492), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2493), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2494), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2495), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2496), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2497), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2498), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2499), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2500), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2501), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2502), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2503), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2504), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2505), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2506), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2507), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2508), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2509), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2510), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2511), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2512), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2513), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2514), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2515), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2516), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2517), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2518), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2519), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2520), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2521), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2522), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2523), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2524), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2525), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2526), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2527), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2528), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2529), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2530), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2531), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2532), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2533), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2534), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2535), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2536), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2537), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2538), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2539), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2540), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2541), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2542), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2543), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2544), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2545), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2546), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2547), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2548), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2549), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2550), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2551), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2552), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2553), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2554), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2555), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2556), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2557), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2558), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2559), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2560), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2561), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2562), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2563), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2564), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2565), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2566), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2567), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2568), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2569), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2570), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2571), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2572), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2573), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2574), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2575), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2576), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2577), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2578), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2579), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2580), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2581), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2582), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2583), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2584), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2585), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2586), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2587), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2588), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2589), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2590), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2591), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2592), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2593), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2594), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2595), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2596), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2597), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2598), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2599), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2600), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2601), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2602), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2603), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2604), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2605), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2606), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2607), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2608), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2609), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2610), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2611), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2612), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2613), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2614), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2615), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2616), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2617), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2618), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2619), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2620), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2621), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2622), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2623), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2624), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2625), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2626), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2627), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2628), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2629), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2630), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2631), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2632), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2633), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2634), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2635), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2636), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2637), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2638), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2639), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2640), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2641), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2642), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2643), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2644), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2645), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2646), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2647), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2648), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2649), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2650), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2651), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2652), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2653), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2654), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2655), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2656), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2657), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2658), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2659), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2660), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2661), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2662), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2663), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2664), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2665), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2666), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2667), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2668), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2669), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2670), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2671), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2672), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2673), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2674), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2675), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2676), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2677), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2678), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2679), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2680), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2681), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2682), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2683), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2684), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2685), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2686), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2687), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2688), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2689), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2690), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2691), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2692), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2693), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2694), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2695), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2696), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2697), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2698), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2699), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2700), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2701), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2702), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2703), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2704), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2705), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2706), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2707), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2708), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2709), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2710), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2711), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2712), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2713), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2714), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2715), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2716), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2717), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2718), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2719), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2720), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2721), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2722), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2723), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2724), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2725), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2726), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2727), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2728), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2729), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2730), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2731), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2732), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2733), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2734), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2735), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2736), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2737), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2738), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2739), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2740), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2741), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2742), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2743), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2744), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2745), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2746), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2747), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2748), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2749), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2750), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2751), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2752), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2753), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2754), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2755), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2756), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2757), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2758), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2759), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2760), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2761), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2762), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2763), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2764), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2765), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2766), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2767), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2768), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2769), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2770), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2771), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2772), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2773), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2774), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2775), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2776), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2777), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2778), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2779), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2780), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2781), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2782), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2783), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2784), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2785), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2786), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2787), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2788), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2789), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2790), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2791), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2792), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2793), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2794), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2795), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2796), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2797), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2798), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2799), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2800), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2801), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2802), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2803), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2804), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2805), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2806), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2807), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2808), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2809), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2810), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2811), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2812), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2813), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2814), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2815), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2816), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2817), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2818), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2819), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2820), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2821), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2822), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2823), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2824), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2825), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2826), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2827), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2828), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2829), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2830), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2831), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2832), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2833), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2834), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2835), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2836), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2837), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2838), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2839), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2840), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2841), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2842), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2843), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2844), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2845), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2846), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2847), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2848), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2849), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2850), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2851), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2852), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2853), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2854), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2855), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2856), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2857), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2858), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2859), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2860), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2861), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2862), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2863), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2864), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2865), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2866), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2867), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2868), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2869), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2870), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2871), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2872), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2873), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2874), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2875), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2876), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2877), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2878), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2879), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2880), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2881), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2882), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2883), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2884), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2885), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2886), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2887), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2888), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2889), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2890), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2891), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2892), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2893), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2894), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2895), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2896), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2897), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2898), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2899), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2900), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2901), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2902), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2903), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2904), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2905), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2906), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2907), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2908), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2909), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2910), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2911), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2912) );
  INVX1 U2 ( .A(n111), .Y(n1) );
  INVX1 U3 ( .A(n113), .Y(n2) );
  INVX1 U4 ( .A(n113), .Y(n3) );
  INVX4 U5 ( .A(n58), .Y(n59) );
  INVX4 U6 ( .A(n18), .Y(n19) );
  INVX4 U7 ( .A(n16), .Y(n17) );
  INVX4 U8 ( .A(n12), .Y(n13) );
  INVX4 U9 ( .A(n10), .Y(n11) );
  INVX4 U10 ( .A(n4), .Y(n5) );
  INVX4 U11 ( .A(n89), .Y(n90) );
  INVX4 U12 ( .A(n24), .Y(n25) );
  INVX4 U13 ( .A(n53), .Y(n54) );
  INVX4 U14 ( .A(n8), .Y(n9) );
  INVX4 U15 ( .A(n60), .Y(n61) );
  INVX4 U16 ( .A(n26), .Y(n27) );
  INVX1 U17 ( .A(n2224), .Y(n2228) );
  INVX1 U18 ( .A(n2384), .Y(n2221) );
  INVX1 U19 ( .A(n2382), .Y(n2222) );
  INVX2 U20 ( .A(n2224), .Y(n2230) );
  INVX1 U21 ( .A(n2224), .Y(n2229) );
  INVX1 U22 ( .A(n2224), .Y(n2225) );
  INVX1 U23 ( .A(n2382), .Y(n2223) );
  INVX2 U24 ( .A(n2224), .Y(n2227) );
  INVX2 U25 ( .A(n2224), .Y(n2226) );
  INVX1 U26 ( .A(n2384), .Y(n2220) );
  INVX1 U27 ( .A(n2210), .Y(N26) );
  INVX1 U28 ( .A(n2212), .Y(N24) );
  INVX2 U29 ( .A(n2231), .Y(n2232) );
  INVX1 U30 ( .A(n2231), .Y(n2234) );
  INVX2 U31 ( .A(n2231), .Y(n2235) );
  INVX2 U32 ( .A(n2231), .Y(n2236) );
  INVX2 U33 ( .A(n2231), .Y(n2237) );
  INVX2 U34 ( .A(n2231), .Y(n2238) );
  INVX2 U35 ( .A(n2231), .Y(n2239) );
  INVX2 U36 ( .A(n2231), .Y(n2240) );
  INVX2 U37 ( .A(n2231), .Y(n2241) );
  INVX1 U38 ( .A(n2204), .Y(N32) );
  INVX1 U39 ( .A(n2205), .Y(N31) );
  INVX1 U40 ( .A(n2206), .Y(N30) );
  INVX1 U41 ( .A(n2207), .Y(N29) );
  INVX1 U42 ( .A(n2208), .Y(N28) );
  INVX1 U43 ( .A(n2209), .Y(N27) );
  INVX1 U44 ( .A(n2211), .Y(N25) );
  INVX1 U45 ( .A(n2214), .Y(N22) );
  INVX1 U46 ( .A(n2215), .Y(N21) );
  INVX1 U47 ( .A(n2217), .Y(N19) );
  INVX1 U48 ( .A(n2218), .Y(N18) );
  INVX1 U49 ( .A(n2219), .Y(N17) );
  INVX1 U50 ( .A(n2213), .Y(N23) );
  INVX1 U51 ( .A(n2216), .Y(N20) );
  BUFX2 U52 ( .A(n1667), .Y(n2275) );
  BUFX2 U53 ( .A(n1669), .Y(n2277) );
  BUFX2 U54 ( .A(n1671), .Y(n2279) );
  BUFX2 U55 ( .A(n1673), .Y(n2281) );
  BUFX2 U56 ( .A(n1675), .Y(n2283) );
  BUFX2 U57 ( .A(n1677), .Y(n2285) );
  BUFX2 U58 ( .A(n1679), .Y(n2288) );
  BUFX2 U59 ( .A(n1681), .Y(n2290) );
  BUFX2 U60 ( .A(n1683), .Y(n2292) );
  BUFX2 U61 ( .A(n1685), .Y(n2295) );
  BUFX2 U62 ( .A(n1687), .Y(n2297) );
  BUFX2 U63 ( .A(n1689), .Y(n2300) );
  BUFX2 U64 ( .A(n1691), .Y(n2303) );
  BUFX2 U65 ( .A(n1693), .Y(n2305) );
  BUFX2 U66 ( .A(n1695), .Y(n2308) );
  BUFX2 U67 ( .A(n1697), .Y(n2310) );
  BUFX2 U68 ( .A(n1699), .Y(n2312) );
  BUFX2 U69 ( .A(n1701), .Y(n2314) );
  BUFX2 U70 ( .A(n1703), .Y(n2316) );
  BUFX2 U71 ( .A(n1705), .Y(n2318) );
  BUFX2 U72 ( .A(n1707), .Y(n2320) );
  BUFX2 U73 ( .A(n1709), .Y(n2323) );
  BUFX2 U74 ( .A(n1711), .Y(n2325) );
  BUFX2 U75 ( .A(n1713), .Y(n2327) );
  BUFX2 U76 ( .A(n1715), .Y(n2329) );
  BUFX2 U77 ( .A(n1717), .Y(n2331) );
  BUFX2 U78 ( .A(n1719), .Y(n2333) );
  BUFX2 U79 ( .A(n1721), .Y(n2335) );
  INVX1 U80 ( .A(n2378), .Y(n2242) );
  INVX2 U81 ( .A(n2379), .Y(n2224) );
  INVX2 U82 ( .A(n2376), .Y(n2272) );
  INVX4 U83 ( .A(n2272), .Y(n2273) );
  INVX1 U84 ( .A(n2384), .Y(n2383) );
  INVX1 U85 ( .A(N14), .Y(n2384) );
  INVX1 U86 ( .A(n2382), .Y(n2381) );
  INVX1 U87 ( .A(N13), .Y(n2382) );
  BUFX2 U88 ( .A(n1669), .Y(n2278) );
  BUFX2 U89 ( .A(n1691), .Y(n2304) );
  BUFX2 U90 ( .A(n1693), .Y(n2306) );
  BUFX2 U91 ( .A(n1671), .Y(n2280) );
  BUFX2 U92 ( .A(n1673), .Y(n2282) );
  BUFX2 U93 ( .A(n1695), .Y(n2309) );
  BUFX2 U94 ( .A(n1697), .Y(n2311) );
  BUFX2 U95 ( .A(n1699), .Y(n2313) );
  BUFX2 U96 ( .A(n1701), .Y(n2315) );
  BUFX2 U97 ( .A(n1703), .Y(n2317) );
  BUFX2 U98 ( .A(n1705), .Y(n2319) );
  BUFX2 U99 ( .A(n1707), .Y(n2321) );
  BUFX2 U100 ( .A(n1709), .Y(n2324) );
  BUFX2 U101 ( .A(n1711), .Y(n2326) );
  BUFX2 U102 ( .A(n1713), .Y(n2328) );
  BUFX2 U103 ( .A(n1715), .Y(n2330) );
  BUFX2 U104 ( .A(n1717), .Y(n2332) );
  BUFX2 U105 ( .A(n1719), .Y(n2334) );
  BUFX2 U106 ( .A(n1721), .Y(n2336) );
  INVX1 U107 ( .A(n1664), .Y(n2322) );
  INVX1 U108 ( .A(n1665), .Y(n2337) );
  BUFX2 U109 ( .A(n1685), .Y(n2296) );
  BUFX2 U110 ( .A(n1687), .Y(n2298) );
  BUFX2 U111 ( .A(n1689), .Y(n2301) );
  INVX1 U112 ( .A(rst), .Y(n2375) );
  BUFX2 U113 ( .A(n1667), .Y(n2276) );
  BUFX2 U114 ( .A(n1675), .Y(n2284) );
  BUFX2 U115 ( .A(n1677), .Y(n2286) );
  BUFX2 U116 ( .A(n1679), .Y(n2289) );
  BUFX2 U117 ( .A(n1681), .Y(n2291) );
  BUFX2 U118 ( .A(n1683), .Y(n2293) );
  INVX1 U119 ( .A(n1663), .Y(n2307) );
  AND2X2 U120 ( .A(n2340), .B(n1674), .Y(n4) );
  AND2X2 U121 ( .A(n2340), .B(n1676), .Y(n6) );
  INVX1 U122 ( .A(n6), .Y(n7) );
  AND2X2 U123 ( .A(n2339), .B(n1678), .Y(n8) );
  AND2X2 U124 ( .A(n2340), .B(n1661), .Y(n10) );
  AND2X2 U125 ( .A(n2340), .B(n1680), .Y(n12) );
  AND2X2 U126 ( .A(n2339), .B(n1682), .Y(n14) );
  INVX1 U127 ( .A(n14), .Y(n15) );
  AND2X2 U128 ( .A(n2340), .B(n1666), .Y(n16) );
  AND2X2 U129 ( .A(n2340), .B(n1684), .Y(n18) );
  AND2X2 U130 ( .A(n2339), .B(n1686), .Y(n20) );
  INVX1 U131 ( .A(n20), .Y(n21) );
  AND2X2 U132 ( .A(n2338), .B(n1688), .Y(n22) );
  INVX1 U133 ( .A(n22), .Y(n23) );
  AND2X2 U134 ( .A(n2339), .B(n1664), .Y(n24) );
  AND2X2 U135 ( .A(n2338), .B(n1665), .Y(n26) );
  OR2X2 U136 ( .A(n1723), .B(n180), .Y(n28) );
  INVX1 U137 ( .A(n28), .Y(\data_out<0> ) );
  AND2X2 U138 ( .A(n2375), .B(n1723), .Y(n30) );
  AND2X2 U139 ( .A(\mem<30><0> ), .B(n54), .Y(n31) );
  INVX1 U140 ( .A(n31), .Y(n32) );
  AND2X2 U141 ( .A(\mem<29><0> ), .B(n56), .Y(n33) );
  INVX1 U142 ( .A(n33), .Y(n34) );
  AND2X2 U143 ( .A(\mem<28><0> ), .B(n59), .Y(n35) );
  INVX1 U144 ( .A(n35), .Y(n36) );
  AND2X2 U145 ( .A(\data_in<0> ), .B(n2340), .Y(n37) );
  AND2X2 U146 ( .A(\data_in<1> ), .B(n2340), .Y(n38) );
  AND2X2 U147 ( .A(\data_in<2> ), .B(n2340), .Y(n39) );
  AND2X2 U148 ( .A(\data_in<3> ), .B(n2340), .Y(n40) );
  AND2X2 U149 ( .A(\data_in<4> ), .B(n2340), .Y(n41) );
  AND2X2 U150 ( .A(\data_in<5> ), .B(n2340), .Y(n42) );
  AND2X2 U151 ( .A(\data_in<6> ), .B(n2340), .Y(n43) );
  AND2X2 U152 ( .A(\data_in<7> ), .B(n2340), .Y(n44) );
  AND2X2 U153 ( .A(\data_in<8> ), .B(n2340), .Y(n45) );
  AND2X2 U154 ( .A(\data_in<9> ), .B(n2340), .Y(n46) );
  AND2X2 U155 ( .A(\data_in<10> ), .B(n2340), .Y(n47) );
  AND2X2 U156 ( .A(\data_in<11> ), .B(n2339), .Y(n48) );
  AND2X2 U157 ( .A(\data_in<12> ), .B(n2339), .Y(n49) );
  AND2X2 U158 ( .A(\data_in<13> ), .B(n2339), .Y(n50) );
  AND2X2 U159 ( .A(\data_in<14> ), .B(n2339), .Y(n51) );
  AND2X2 U160 ( .A(\data_in<15> ), .B(n2339), .Y(n52) );
  AND2X2 U161 ( .A(n2339), .B(n1668), .Y(n53) );
  AND2X2 U162 ( .A(n2339), .B(n1670), .Y(n55) );
  INVX1 U163 ( .A(n55), .Y(n56) );
  INVX1 U164 ( .A(n55), .Y(n57) );
  AND2X2 U165 ( .A(n2340), .B(n1672), .Y(n58) );
  AND2X2 U166 ( .A(n2338), .B(n1690), .Y(n60) );
  AND2X2 U167 ( .A(n2338), .B(n1692), .Y(n62) );
  INVX1 U168 ( .A(n62), .Y(n63) );
  INVX1 U169 ( .A(n62), .Y(n64) );
  AND2X2 U170 ( .A(n2338), .B(n1663), .Y(n65) );
  INVX1 U171 ( .A(n65), .Y(n66) );
  INVX1 U172 ( .A(n65), .Y(n67) );
  AND2X2 U173 ( .A(n2338), .B(n1694), .Y(n68) );
  INVX1 U174 ( .A(n68), .Y(n69) );
  INVX1 U175 ( .A(n68), .Y(n70) );
  AND2X2 U176 ( .A(n2338), .B(n1696), .Y(n71) );
  INVX1 U177 ( .A(n71), .Y(n72) );
  INVX1 U178 ( .A(n71), .Y(n73) );
  AND2X2 U179 ( .A(n2338), .B(n1698), .Y(n74) );
  INVX1 U180 ( .A(n74), .Y(n75) );
  INVX1 U181 ( .A(n74), .Y(n76) );
  AND2X2 U182 ( .A(n2338), .B(n1700), .Y(n77) );
  INVX1 U183 ( .A(n77), .Y(n78) );
  INVX1 U184 ( .A(n77), .Y(n79) );
  AND2X2 U185 ( .A(n2338), .B(n1702), .Y(n80) );
  INVX1 U186 ( .A(n80), .Y(n81) );
  INVX1 U187 ( .A(n80), .Y(n82) );
  AND2X2 U188 ( .A(n2338), .B(n1704), .Y(n83) );
  INVX1 U189 ( .A(n83), .Y(n84) );
  INVX1 U190 ( .A(n83), .Y(n85) );
  AND2X2 U191 ( .A(n2338), .B(n1706), .Y(n86) );
  INVX1 U192 ( .A(n86), .Y(n87) );
  INVX1 U193 ( .A(n86), .Y(n88) );
  AND2X2 U194 ( .A(n2339), .B(n1708), .Y(n89) );
  AND2X2 U195 ( .A(n2339), .B(n1710), .Y(n91) );
  INVX1 U196 ( .A(n91), .Y(n92) );
  INVX1 U197 ( .A(n91), .Y(n93) );
  AND2X2 U198 ( .A(n2339), .B(n1712), .Y(n94) );
  INVX1 U199 ( .A(n94), .Y(n95) );
  INVX1 U200 ( .A(n94), .Y(n96) );
  AND2X2 U201 ( .A(n2339), .B(n1714), .Y(n97) );
  INVX1 U202 ( .A(n97), .Y(n98) );
  INVX1 U203 ( .A(n97), .Y(n99) );
  AND2X2 U204 ( .A(n2339), .B(n1716), .Y(n100) );
  INVX1 U205 ( .A(n100), .Y(n101) );
  INVX1 U206 ( .A(n100), .Y(n102) );
  AND2X2 U207 ( .A(n2339), .B(n1718), .Y(n103) );
  INVX1 U208 ( .A(n103), .Y(n104) );
  INVX1 U209 ( .A(n103), .Y(n105) );
  AND2X2 U210 ( .A(n2339), .B(n1720), .Y(n106) );
  INVX1 U211 ( .A(n106), .Y(n107) );
  INVX1 U212 ( .A(n106), .Y(n108) );
  INVX1 U213 ( .A(n113), .Y(n109) );
  INVX1 U214 ( .A(n111), .Y(n110) );
  OR2X2 U215 ( .A(write), .B(rst), .Y(n111) );
  INVX1 U216 ( .A(n111), .Y(n112) );
  OR2X2 U217 ( .A(write), .B(rst), .Y(n113) );
  INVX1 U218 ( .A(n113), .Y(n114) );
  INVX4 U219 ( .A(n2342), .Y(n2338) );
  AND2X2 U220 ( .A(\mem<23><0> ), .B(n13), .Y(n115) );
  INVX1 U221 ( .A(n115), .Y(n116) );
  AND2X2 U222 ( .A(\mem<23><1> ), .B(n13), .Y(n117) );
  INVX1 U223 ( .A(n117), .Y(n118) );
  AND2X2 U224 ( .A(\mem<23><2> ), .B(n13), .Y(n119) );
  INVX1 U225 ( .A(n119), .Y(n120) );
  AND2X2 U226 ( .A(\mem<23><3> ), .B(n13), .Y(n121) );
  INVX1 U227 ( .A(n121), .Y(n122) );
  AND2X2 U228 ( .A(\mem<23><4> ), .B(n13), .Y(n123) );
  INVX1 U229 ( .A(n123), .Y(n124) );
  AND2X2 U230 ( .A(\mem<23><5> ), .B(n13), .Y(n125) );
  INVX1 U231 ( .A(n125), .Y(n126) );
  AND2X2 U232 ( .A(\mem<23><6> ), .B(n13), .Y(n127) );
  INVX1 U233 ( .A(n127), .Y(n128) );
  AND2X2 U234 ( .A(\mem<23><7> ), .B(n13), .Y(n129) );
  INVX1 U235 ( .A(n129), .Y(n130) );
  AND2X2 U236 ( .A(\mem<22><0> ), .B(n2294), .Y(n131) );
  INVX1 U237 ( .A(n131), .Y(n132) );
  AND2X2 U238 ( .A(\mem<22><1> ), .B(n2294), .Y(n133) );
  INVX1 U239 ( .A(n133), .Y(n134) );
  AND2X2 U240 ( .A(\mem<22><2> ), .B(n2294), .Y(n135) );
  INVX1 U241 ( .A(n135), .Y(n136) );
  AND2X2 U242 ( .A(\mem<22><3> ), .B(n2294), .Y(n137) );
  INVX1 U243 ( .A(n137), .Y(n138) );
  AND2X2 U244 ( .A(\mem<22><4> ), .B(n2294), .Y(n139) );
  INVX1 U245 ( .A(n139), .Y(n140) );
  AND2X2 U246 ( .A(\mem<22><5> ), .B(n2294), .Y(n141) );
  INVX1 U247 ( .A(n141), .Y(n142) );
  AND2X2 U248 ( .A(\mem<22><6> ), .B(n2294), .Y(n143) );
  INVX1 U249 ( .A(n143), .Y(n144) );
  AND2X2 U250 ( .A(\mem<22><7> ), .B(n2294), .Y(n145) );
  INVX1 U251 ( .A(n145), .Y(n146) );
  AND2X2 U252 ( .A(\mem<21><0> ), .B(n19), .Y(n147) );
  INVX1 U253 ( .A(n147), .Y(n148) );
  AND2X2 U254 ( .A(\mem<21><1> ), .B(n19), .Y(n149) );
  INVX1 U255 ( .A(n149), .Y(n150) );
  AND2X2 U256 ( .A(\mem<21><2> ), .B(n19), .Y(n151) );
  INVX1 U257 ( .A(n151), .Y(n152) );
  AND2X2 U258 ( .A(\mem<21><3> ), .B(n19), .Y(n153) );
  INVX1 U259 ( .A(n153), .Y(n154) );
  AND2X2 U260 ( .A(\mem<21><4> ), .B(n19), .Y(n155) );
  INVX1 U261 ( .A(n155), .Y(n156) );
  AND2X2 U262 ( .A(\mem<21><5> ), .B(n19), .Y(n157) );
  INVX1 U263 ( .A(n157), .Y(n158) );
  AND2X2 U264 ( .A(\mem<21><6> ), .B(n19), .Y(n159) );
  INVX1 U265 ( .A(n159), .Y(n160) );
  AND2X2 U266 ( .A(\mem<21><7> ), .B(n19), .Y(n161) );
  INVX1 U267 ( .A(n161), .Y(n162) );
  AND2X2 U268 ( .A(\mem<20><0> ), .B(n2299), .Y(n163) );
  INVX1 U269 ( .A(n163), .Y(n164) );
  AND2X2 U270 ( .A(\mem<20><1> ), .B(n2299), .Y(n165) );
  INVX1 U271 ( .A(n165), .Y(n166) );
  AND2X2 U272 ( .A(\mem<20><2> ), .B(n2299), .Y(n167) );
  INVX1 U273 ( .A(n167), .Y(n168) );
  AND2X2 U274 ( .A(\mem<20><3> ), .B(n2299), .Y(n169) );
  INVX1 U275 ( .A(n169), .Y(n170) );
  AND2X2 U276 ( .A(\mem<20><4> ), .B(n2299), .Y(n171) );
  INVX1 U277 ( .A(n171), .Y(n172) );
  AND2X2 U278 ( .A(\mem<20><5> ), .B(n2299), .Y(n173) );
  INVX1 U279 ( .A(n173), .Y(n174) );
  AND2X2 U280 ( .A(\mem<20><6> ), .B(n2299), .Y(n175) );
  INVX1 U281 ( .A(n175), .Y(n176) );
  AND2X2 U282 ( .A(\mem<20><7> ), .B(n2299), .Y(n177) );
  INVX1 U283 ( .A(n177), .Y(n178) );
  AND2X1 U284 ( .A(n2375), .B(N32), .Y(n179) );
  INVX1 U285 ( .A(n179), .Y(n180) );
  INVX1 U286 ( .A(n2377), .Y(n2376) );
  INVX1 U287 ( .A(n2380), .Y(n2379) );
  AND2X1 U288 ( .A(n2379), .B(n2233), .Y(n181) );
  AND2X1 U289 ( .A(n2912), .B(n2383), .Y(n182) );
  AND2X2 U290 ( .A(\mem<31><0> ), .B(n17), .Y(n183) );
  INVX1 U291 ( .A(n183), .Y(n184) );
  AND2X2 U292 ( .A(\mem<31><1> ), .B(n17), .Y(n185) );
  INVX1 U293 ( .A(n185), .Y(n186) );
  AND2X2 U294 ( .A(\mem<31><2> ), .B(n17), .Y(n187) );
  INVX1 U295 ( .A(n187), .Y(n188) );
  AND2X2 U296 ( .A(\mem<31><3> ), .B(n17), .Y(n189) );
  INVX1 U297 ( .A(n189), .Y(n190) );
  AND2X2 U298 ( .A(\mem<31><4> ), .B(n17), .Y(n191) );
  INVX1 U299 ( .A(n191), .Y(n192) );
  AND2X2 U300 ( .A(\mem<31><5> ), .B(n17), .Y(n193) );
  INVX1 U301 ( .A(n193), .Y(n194) );
  AND2X2 U302 ( .A(\mem<31><6> ), .B(n17), .Y(n195) );
  INVX1 U303 ( .A(n195), .Y(n196) );
  AND2X2 U304 ( .A(\mem<31><7> ), .B(n17), .Y(n197) );
  INVX1 U305 ( .A(n197), .Y(n198) );
  AND2X2 U306 ( .A(\mem<31><8> ), .B(n17), .Y(n199) );
  INVX1 U307 ( .A(n199), .Y(n200) );
  AND2X2 U308 ( .A(\mem<31><9> ), .B(n17), .Y(n201) );
  INVX1 U309 ( .A(n201), .Y(n202) );
  AND2X2 U310 ( .A(\mem<31><10> ), .B(n17), .Y(n203) );
  INVX1 U311 ( .A(n203), .Y(n204) );
  AND2X2 U312 ( .A(\mem<31><11> ), .B(n17), .Y(n205) );
  INVX1 U313 ( .A(n205), .Y(n206) );
  AND2X2 U314 ( .A(\mem<31><12> ), .B(n17), .Y(n207) );
  INVX1 U315 ( .A(n207), .Y(n208) );
  AND2X2 U316 ( .A(\mem<31><13> ), .B(n17), .Y(n209) );
  INVX1 U317 ( .A(n209), .Y(n210) );
  AND2X2 U318 ( .A(\mem<31><14> ), .B(n17), .Y(n211) );
  INVX1 U319 ( .A(n211), .Y(n212) );
  AND2X2 U320 ( .A(\mem<31><15> ), .B(n17), .Y(n213) );
  INVX1 U321 ( .A(n213), .Y(n215) );
  AND2X2 U322 ( .A(\mem<30><1> ), .B(n54), .Y(n216) );
  INVX1 U323 ( .A(n216), .Y(n217) );
  AND2X2 U324 ( .A(\mem<30><2> ), .B(n54), .Y(n218) );
  INVX1 U325 ( .A(n218), .Y(n219) );
  AND2X2 U326 ( .A(\mem<30><3> ), .B(n54), .Y(n220) );
  INVX1 U327 ( .A(n220), .Y(n221) );
  AND2X2 U328 ( .A(\mem<30><4> ), .B(n54), .Y(n222) );
  INVX1 U329 ( .A(n222), .Y(n223) );
  AND2X2 U330 ( .A(\mem<30><5> ), .B(n54), .Y(n224) );
  INVX1 U331 ( .A(n224), .Y(n225) );
  AND2X2 U332 ( .A(\mem<30><6> ), .B(n54), .Y(n226) );
  INVX1 U333 ( .A(n226), .Y(n227) );
  AND2X2 U334 ( .A(\mem<30><7> ), .B(n54), .Y(n228) );
  INVX1 U335 ( .A(n228), .Y(n229) );
  AND2X2 U336 ( .A(\mem<30><8> ), .B(n54), .Y(n230) );
  INVX1 U337 ( .A(n230), .Y(n231) );
  AND2X2 U338 ( .A(\mem<30><9> ), .B(n54), .Y(n232) );
  INVX1 U339 ( .A(n232), .Y(n233) );
  AND2X2 U340 ( .A(\mem<30><10> ), .B(n54), .Y(n234) );
  INVX1 U341 ( .A(n234), .Y(n235) );
  AND2X2 U342 ( .A(\mem<30><11> ), .B(n54), .Y(n236) );
  INVX1 U343 ( .A(n236), .Y(n237) );
  AND2X2 U344 ( .A(\mem<30><12> ), .B(n54), .Y(n238) );
  INVX1 U345 ( .A(n238), .Y(n239) );
  AND2X2 U346 ( .A(\mem<30><13> ), .B(n54), .Y(n240) );
  INVX1 U347 ( .A(n240), .Y(n241) );
  AND2X2 U348 ( .A(\mem<30><14> ), .B(n54), .Y(n242) );
  INVX1 U349 ( .A(n242), .Y(n243) );
  AND2X2 U350 ( .A(\mem<30><15> ), .B(n54), .Y(n244) );
  INVX1 U351 ( .A(n244), .Y(n245) );
  AND2X2 U352 ( .A(\mem<29><1> ), .B(n56), .Y(n246) );
  INVX1 U353 ( .A(n246), .Y(n247) );
  AND2X2 U354 ( .A(\mem<29><2> ), .B(n56), .Y(n248) );
  INVX1 U355 ( .A(n248), .Y(n249) );
  AND2X2 U356 ( .A(\mem<29><3> ), .B(n56), .Y(n250) );
  INVX1 U357 ( .A(n250), .Y(n251) );
  AND2X2 U358 ( .A(\mem<29><4> ), .B(n56), .Y(n252) );
  INVX1 U359 ( .A(n252), .Y(n253) );
  AND2X2 U360 ( .A(\mem<29><5> ), .B(n56), .Y(n254) );
  INVX1 U361 ( .A(n254), .Y(n255) );
  AND2X2 U362 ( .A(\mem<29><6> ), .B(n56), .Y(n256) );
  INVX1 U363 ( .A(n256), .Y(n257) );
  AND2X2 U364 ( .A(\mem<29><7> ), .B(n56), .Y(n258) );
  INVX1 U365 ( .A(n258), .Y(n259) );
  AND2X2 U366 ( .A(\mem<29><8> ), .B(n57), .Y(n260) );
  INVX1 U367 ( .A(n260), .Y(n261) );
  AND2X2 U368 ( .A(\mem<29><9> ), .B(n57), .Y(n262) );
  INVX1 U369 ( .A(n262), .Y(n263) );
  AND2X2 U370 ( .A(\mem<29><10> ), .B(n57), .Y(n264) );
  INVX1 U371 ( .A(n264), .Y(n265) );
  AND2X2 U372 ( .A(\mem<29><11> ), .B(n57), .Y(n266) );
  INVX1 U373 ( .A(n266), .Y(n267) );
  AND2X2 U374 ( .A(\mem<29><12> ), .B(n57), .Y(n268) );
  INVX1 U375 ( .A(n268), .Y(n269) );
  AND2X2 U376 ( .A(\mem<29><13> ), .B(n57), .Y(n270) );
  INVX1 U377 ( .A(n270), .Y(n271) );
  AND2X2 U378 ( .A(\mem<29><14> ), .B(n57), .Y(n272) );
  INVX1 U379 ( .A(n272), .Y(n273) );
  AND2X2 U380 ( .A(\mem<29><15> ), .B(n57), .Y(n274) );
  INVX1 U381 ( .A(n274), .Y(n275) );
  AND2X2 U382 ( .A(\mem<28><1> ), .B(n59), .Y(n276) );
  INVX1 U383 ( .A(n276), .Y(n277) );
  AND2X2 U384 ( .A(\mem<28><2> ), .B(n59), .Y(n278) );
  INVX1 U385 ( .A(n278), .Y(n279) );
  AND2X2 U386 ( .A(\mem<28><3> ), .B(n59), .Y(n280) );
  INVX1 U387 ( .A(n280), .Y(n281) );
  AND2X2 U388 ( .A(\mem<28><4> ), .B(n59), .Y(n282) );
  INVX1 U389 ( .A(n282), .Y(n283) );
  AND2X2 U390 ( .A(\mem<28><5> ), .B(n59), .Y(n284) );
  INVX1 U391 ( .A(n284), .Y(n285) );
  AND2X2 U392 ( .A(\mem<28><6> ), .B(n59), .Y(n286) );
  INVX1 U393 ( .A(n286), .Y(n287) );
  AND2X2 U394 ( .A(\mem<28><7> ), .B(n59), .Y(n288) );
  INVX1 U395 ( .A(n288), .Y(n289) );
  AND2X2 U396 ( .A(\mem<28><8> ), .B(n59), .Y(n290) );
  INVX1 U397 ( .A(n290), .Y(n291) );
  AND2X2 U398 ( .A(\mem<28><9> ), .B(n59), .Y(n292) );
  INVX1 U399 ( .A(n292), .Y(n293) );
  AND2X2 U400 ( .A(\mem<28><10> ), .B(n59), .Y(n294) );
  INVX1 U401 ( .A(n294), .Y(n295) );
  AND2X2 U402 ( .A(\mem<28><11> ), .B(n59), .Y(n296) );
  INVX1 U403 ( .A(n296), .Y(n297) );
  AND2X2 U404 ( .A(\mem<28><12> ), .B(n59), .Y(n298) );
  INVX1 U405 ( .A(n298), .Y(n299) );
  AND2X2 U406 ( .A(\mem<28><13> ), .B(n59), .Y(n300) );
  INVX1 U407 ( .A(n300), .Y(n301) );
  AND2X2 U408 ( .A(\mem<28><14> ), .B(n59), .Y(n302) );
  INVX1 U409 ( .A(n302), .Y(n303) );
  AND2X2 U410 ( .A(\mem<28><15> ), .B(n59), .Y(n304) );
  INVX1 U411 ( .A(n304), .Y(n305) );
  AND2X2 U412 ( .A(\mem<27><0> ), .B(n5), .Y(n306) );
  INVX1 U413 ( .A(n306), .Y(n307) );
  AND2X2 U414 ( .A(\mem<27><1> ), .B(n5), .Y(n308) );
  INVX1 U415 ( .A(n308), .Y(n309) );
  AND2X2 U416 ( .A(\mem<27><2> ), .B(n5), .Y(n310) );
  INVX1 U417 ( .A(n310), .Y(n311) );
  AND2X2 U418 ( .A(\mem<27><3> ), .B(n5), .Y(n312) );
  INVX1 U419 ( .A(n312), .Y(n313) );
  AND2X2 U420 ( .A(\mem<27><4> ), .B(n5), .Y(n314) );
  INVX1 U421 ( .A(n314), .Y(n315) );
  AND2X2 U422 ( .A(\mem<27><5> ), .B(n5), .Y(n316) );
  INVX1 U423 ( .A(n316), .Y(n317) );
  AND2X2 U424 ( .A(\mem<27><6> ), .B(n5), .Y(n318) );
  INVX1 U425 ( .A(n318), .Y(n319) );
  AND2X2 U426 ( .A(\mem<27><7> ), .B(n5), .Y(n320) );
  INVX1 U427 ( .A(n320), .Y(n321) );
  AND2X2 U428 ( .A(\mem<27><8> ), .B(n5), .Y(n322) );
  INVX1 U429 ( .A(n322), .Y(n323) );
  AND2X2 U430 ( .A(\mem<27><9> ), .B(n5), .Y(n324) );
  INVX1 U431 ( .A(n324), .Y(n325) );
  AND2X2 U432 ( .A(\mem<27><10> ), .B(n5), .Y(n326) );
  INVX1 U433 ( .A(n326), .Y(n327) );
  AND2X2 U434 ( .A(\mem<27><11> ), .B(n5), .Y(n328) );
  INVX1 U435 ( .A(n328), .Y(n329) );
  AND2X2 U436 ( .A(\mem<27><12> ), .B(n5), .Y(n330) );
  INVX1 U437 ( .A(n330), .Y(n331) );
  AND2X2 U438 ( .A(\mem<27><13> ), .B(n5), .Y(n332) );
  INVX1 U439 ( .A(n332), .Y(n333) );
  AND2X2 U440 ( .A(\mem<27><14> ), .B(n5), .Y(n334) );
  INVX1 U441 ( .A(n334), .Y(n335) );
  AND2X2 U442 ( .A(\mem<27><15> ), .B(n5), .Y(n336) );
  INVX1 U443 ( .A(n336), .Y(n337) );
  AND2X2 U444 ( .A(\mem<26><0> ), .B(n2287), .Y(n338) );
  INVX1 U445 ( .A(n338), .Y(n339) );
  AND2X2 U446 ( .A(\mem<26><1> ), .B(n2287), .Y(n340) );
  INVX1 U447 ( .A(n340), .Y(n341) );
  AND2X2 U448 ( .A(\mem<26><2> ), .B(n2287), .Y(n342) );
  INVX1 U449 ( .A(n342), .Y(n343) );
  AND2X2 U450 ( .A(\mem<26><3> ), .B(n2287), .Y(n344) );
  INVX1 U451 ( .A(n344), .Y(n345) );
  AND2X2 U452 ( .A(\mem<26><4> ), .B(n2287), .Y(n346) );
  INVX1 U453 ( .A(n346), .Y(n347) );
  AND2X2 U454 ( .A(\mem<26><5> ), .B(n2287), .Y(n348) );
  INVX1 U455 ( .A(n348), .Y(n349) );
  AND2X2 U456 ( .A(\mem<26><6> ), .B(n2287), .Y(n350) );
  INVX1 U457 ( .A(n350), .Y(n351) );
  AND2X2 U458 ( .A(\mem<26><7> ), .B(n2287), .Y(n352) );
  INVX1 U459 ( .A(n352), .Y(n353) );
  AND2X2 U460 ( .A(\mem<26><8> ), .B(n2287), .Y(n354) );
  INVX1 U461 ( .A(n354), .Y(n355) );
  AND2X2 U462 ( .A(\mem<26><9> ), .B(n2287), .Y(n356) );
  INVX1 U463 ( .A(n356), .Y(n357) );
  AND2X2 U464 ( .A(\mem<26><10> ), .B(n2287), .Y(n358) );
  INVX1 U465 ( .A(n358), .Y(n359) );
  AND2X2 U466 ( .A(\mem<26><11> ), .B(n2287), .Y(n360) );
  INVX1 U467 ( .A(n360), .Y(n361) );
  AND2X2 U468 ( .A(\mem<26><12> ), .B(n2287), .Y(n362) );
  INVX1 U469 ( .A(n362), .Y(n363) );
  AND2X2 U470 ( .A(\mem<26><13> ), .B(n2287), .Y(n364) );
  INVX1 U471 ( .A(n364), .Y(n365) );
  AND2X2 U472 ( .A(\mem<26><14> ), .B(n2287), .Y(n366) );
  INVX1 U473 ( .A(n366), .Y(n367) );
  AND2X2 U474 ( .A(\mem<26><15> ), .B(n2287), .Y(n368) );
  INVX1 U475 ( .A(n368), .Y(n369) );
  AND2X2 U476 ( .A(\mem<25><0> ), .B(n9), .Y(n370) );
  INVX1 U477 ( .A(n370), .Y(n371) );
  AND2X2 U478 ( .A(\mem<25><1> ), .B(n9), .Y(n372) );
  INVX1 U479 ( .A(n372), .Y(n373) );
  AND2X2 U480 ( .A(\mem<25><2> ), .B(n9), .Y(n374) );
  INVX1 U481 ( .A(n374), .Y(n375) );
  AND2X2 U482 ( .A(\mem<25><3> ), .B(n9), .Y(n376) );
  INVX1 U483 ( .A(n376), .Y(n377) );
  AND2X2 U484 ( .A(\mem<25><4> ), .B(n9), .Y(n378) );
  INVX1 U485 ( .A(n378), .Y(n379) );
  AND2X2 U486 ( .A(\mem<25><5> ), .B(n9), .Y(n380) );
  INVX1 U487 ( .A(n380), .Y(n381) );
  AND2X2 U488 ( .A(\mem<25><6> ), .B(n9), .Y(n382) );
  INVX1 U489 ( .A(n382), .Y(n383) );
  AND2X2 U490 ( .A(\mem<25><7> ), .B(n9), .Y(n384) );
  INVX1 U491 ( .A(n384), .Y(n385) );
  AND2X2 U492 ( .A(\mem<25><8> ), .B(n9), .Y(n386) );
  INVX1 U493 ( .A(n386), .Y(n387) );
  AND2X2 U494 ( .A(\mem<25><9> ), .B(n9), .Y(n388) );
  INVX1 U495 ( .A(n388), .Y(n389) );
  AND2X2 U496 ( .A(\mem<25><10> ), .B(n9), .Y(n390) );
  INVX1 U497 ( .A(n390), .Y(n391) );
  AND2X2 U498 ( .A(\mem<25><11> ), .B(n9), .Y(n392) );
  INVX1 U499 ( .A(n392), .Y(n393) );
  AND2X2 U500 ( .A(\mem<25><12> ), .B(n9), .Y(n394) );
  INVX1 U501 ( .A(n394), .Y(n395) );
  AND2X2 U502 ( .A(\mem<25><13> ), .B(n9), .Y(n396) );
  INVX1 U503 ( .A(n396), .Y(n397) );
  AND2X2 U504 ( .A(\mem<25><14> ), .B(n9), .Y(n398) );
  INVX1 U505 ( .A(n398), .Y(n399) );
  AND2X2 U506 ( .A(\mem<25><15> ), .B(n9), .Y(n400) );
  INVX1 U507 ( .A(n400), .Y(n401) );
  AND2X2 U508 ( .A(\mem<24><0> ), .B(n11), .Y(n402) );
  INVX1 U509 ( .A(n402), .Y(n403) );
  AND2X2 U510 ( .A(\mem<24><1> ), .B(n11), .Y(n404) );
  INVX1 U511 ( .A(n404), .Y(n405) );
  AND2X2 U512 ( .A(\mem<24><2> ), .B(n11), .Y(n406) );
  INVX1 U513 ( .A(n406), .Y(n407) );
  AND2X2 U514 ( .A(\mem<24><3> ), .B(n11), .Y(n408) );
  INVX1 U515 ( .A(n408), .Y(n409) );
  AND2X2 U516 ( .A(\mem<24><4> ), .B(n11), .Y(n410) );
  INVX1 U517 ( .A(n410), .Y(n411) );
  AND2X2 U518 ( .A(\mem<24><5> ), .B(n11), .Y(n412) );
  INVX1 U519 ( .A(n412), .Y(n413) );
  AND2X2 U520 ( .A(\mem<24><6> ), .B(n11), .Y(n414) );
  INVX1 U521 ( .A(n414), .Y(n415) );
  AND2X2 U522 ( .A(\mem<24><7> ), .B(n11), .Y(n416) );
  INVX1 U523 ( .A(n416), .Y(n417) );
  AND2X2 U524 ( .A(\mem<24><8> ), .B(n11), .Y(n418) );
  INVX1 U525 ( .A(n418), .Y(n419) );
  AND2X2 U526 ( .A(\mem<24><9> ), .B(n11), .Y(n420) );
  INVX1 U527 ( .A(n420), .Y(n421) );
  AND2X2 U528 ( .A(\mem<24><10> ), .B(n11), .Y(n422) );
  INVX1 U529 ( .A(n422), .Y(n423) );
  AND2X2 U530 ( .A(\mem<24><11> ), .B(n11), .Y(n424) );
  INVX1 U531 ( .A(n424), .Y(n425) );
  AND2X2 U532 ( .A(\mem<24><12> ), .B(n11), .Y(n426) );
  INVX1 U533 ( .A(n426), .Y(n427) );
  AND2X2 U534 ( .A(\mem<24><13> ), .B(n11), .Y(n428) );
  INVX1 U535 ( .A(n428), .Y(n429) );
  AND2X2 U536 ( .A(\mem<24><14> ), .B(n11), .Y(n430) );
  INVX1 U537 ( .A(n430), .Y(n431) );
  AND2X2 U538 ( .A(\mem<24><15> ), .B(n11), .Y(n432) );
  INVX1 U539 ( .A(n432), .Y(n433) );
  AND2X2 U540 ( .A(\mem<23><8> ), .B(n13), .Y(n434) );
  INVX1 U541 ( .A(n434), .Y(n435) );
  AND2X2 U542 ( .A(\mem<23><9> ), .B(n13), .Y(n436) );
  INVX1 U543 ( .A(n436), .Y(n437) );
  AND2X2 U544 ( .A(\mem<23><10> ), .B(n13), .Y(n438) );
  INVX1 U545 ( .A(n438), .Y(n439) );
  AND2X2 U546 ( .A(\mem<23><11> ), .B(n13), .Y(n440) );
  INVX1 U547 ( .A(n440), .Y(n441) );
  AND2X2 U548 ( .A(\mem<23><12> ), .B(n13), .Y(n442) );
  INVX1 U549 ( .A(n442), .Y(n443) );
  AND2X2 U550 ( .A(\mem<23><13> ), .B(n13), .Y(n444) );
  INVX1 U551 ( .A(n444), .Y(n445) );
  AND2X2 U552 ( .A(\mem<23><14> ), .B(n13), .Y(n446) );
  INVX1 U553 ( .A(n446), .Y(n447) );
  AND2X2 U554 ( .A(\mem<23><15> ), .B(n13), .Y(n448) );
  INVX1 U555 ( .A(n448), .Y(n449) );
  AND2X2 U556 ( .A(\mem<22><8> ), .B(n2294), .Y(n450) );
  INVX1 U557 ( .A(n450), .Y(n451) );
  AND2X2 U558 ( .A(\mem<22><9> ), .B(n2294), .Y(n452) );
  INVX1 U559 ( .A(n452), .Y(n453) );
  AND2X2 U560 ( .A(\mem<22><10> ), .B(n2294), .Y(n454) );
  INVX1 U561 ( .A(n454), .Y(n455) );
  AND2X2 U562 ( .A(\mem<22><11> ), .B(n2294), .Y(n456) );
  INVX1 U563 ( .A(n456), .Y(n457) );
  AND2X2 U564 ( .A(\mem<22><12> ), .B(n2294), .Y(n458) );
  INVX1 U565 ( .A(n458), .Y(n459) );
  AND2X2 U566 ( .A(\mem<22><13> ), .B(n2294), .Y(n460) );
  INVX1 U567 ( .A(n460), .Y(n461) );
  AND2X2 U568 ( .A(\mem<22><14> ), .B(n2294), .Y(n462) );
  INVX1 U569 ( .A(n462), .Y(n463) );
  AND2X2 U570 ( .A(\mem<22><15> ), .B(n2294), .Y(n464) );
  INVX1 U571 ( .A(n464), .Y(n465) );
  AND2X2 U572 ( .A(\mem<21><8> ), .B(n19), .Y(n466) );
  INVX1 U573 ( .A(n466), .Y(n467) );
  AND2X2 U574 ( .A(\mem<21><9> ), .B(n19), .Y(n468) );
  INVX1 U575 ( .A(n468), .Y(n469) );
  AND2X2 U576 ( .A(\mem<21><10> ), .B(n19), .Y(n470) );
  INVX1 U577 ( .A(n470), .Y(n471) );
  AND2X2 U578 ( .A(\mem<21><11> ), .B(n19), .Y(n472) );
  INVX1 U579 ( .A(n472), .Y(n473) );
  AND2X2 U580 ( .A(\mem<21><12> ), .B(n19), .Y(n474) );
  INVX1 U581 ( .A(n474), .Y(n475) );
  AND2X2 U582 ( .A(\mem<21><13> ), .B(n19), .Y(n476) );
  INVX1 U583 ( .A(n476), .Y(n477) );
  AND2X2 U584 ( .A(\mem<21><14> ), .B(n19), .Y(n478) );
  INVX1 U585 ( .A(n478), .Y(n479) );
  AND2X2 U586 ( .A(\mem<21><15> ), .B(n19), .Y(n480) );
  INVX1 U587 ( .A(n480), .Y(n481) );
  AND2X2 U588 ( .A(\mem<20><8> ), .B(n2299), .Y(n482) );
  INVX1 U589 ( .A(n482), .Y(n483) );
  AND2X2 U590 ( .A(\mem<20><9> ), .B(n2299), .Y(n484) );
  INVX1 U591 ( .A(n484), .Y(n485) );
  AND2X2 U592 ( .A(\mem<20><10> ), .B(n2299), .Y(n486) );
  INVX1 U593 ( .A(n486), .Y(n487) );
  AND2X2 U594 ( .A(\mem<20><11> ), .B(n2299), .Y(n488) );
  INVX1 U595 ( .A(n488), .Y(n489) );
  AND2X2 U596 ( .A(\mem<20><12> ), .B(n2299), .Y(n490) );
  INVX1 U597 ( .A(n490), .Y(n491) );
  AND2X2 U598 ( .A(\mem<20><13> ), .B(n2299), .Y(n492) );
  INVX1 U599 ( .A(n492), .Y(n493) );
  AND2X2 U600 ( .A(\mem<20><14> ), .B(n2299), .Y(n494) );
  INVX1 U601 ( .A(n494), .Y(n495) );
  AND2X2 U602 ( .A(\mem<20><15> ), .B(n2299), .Y(n496) );
  INVX1 U603 ( .A(n496), .Y(n497) );
  AND2X2 U604 ( .A(\mem<19><0> ), .B(n2302), .Y(n498) );
  INVX1 U605 ( .A(n498), .Y(n499) );
  AND2X2 U606 ( .A(\mem<19><1> ), .B(n2302), .Y(n500) );
  INVX1 U607 ( .A(n500), .Y(n501) );
  AND2X2 U608 ( .A(\mem<19><2> ), .B(n2302), .Y(n502) );
  INVX1 U609 ( .A(n502), .Y(n503) );
  AND2X2 U610 ( .A(\mem<19><3> ), .B(n2302), .Y(n504) );
  INVX1 U611 ( .A(n504), .Y(n505) );
  AND2X2 U612 ( .A(\mem<19><4> ), .B(n2302), .Y(n506) );
  INVX1 U613 ( .A(n506), .Y(n507) );
  AND2X2 U614 ( .A(\mem<19><5> ), .B(n2302), .Y(n508) );
  INVX1 U615 ( .A(n508), .Y(n509) );
  AND2X2 U616 ( .A(\mem<19><6> ), .B(n2302), .Y(n510) );
  INVX1 U617 ( .A(n510), .Y(n511) );
  AND2X2 U618 ( .A(\mem<19><7> ), .B(n2302), .Y(n512) );
  INVX1 U619 ( .A(n512), .Y(n513) );
  AND2X2 U620 ( .A(\mem<19><8> ), .B(n2302), .Y(n514) );
  INVX1 U621 ( .A(n514), .Y(n515) );
  AND2X2 U622 ( .A(\mem<19><9> ), .B(n2302), .Y(n516) );
  INVX1 U623 ( .A(n516), .Y(n517) );
  AND2X2 U624 ( .A(\mem<19><10> ), .B(n2302), .Y(n518) );
  INVX1 U625 ( .A(n518), .Y(n519) );
  AND2X2 U626 ( .A(\mem<19><11> ), .B(n2302), .Y(n520) );
  INVX1 U627 ( .A(n520), .Y(n521) );
  AND2X2 U628 ( .A(\mem<19><12> ), .B(n2302), .Y(n522) );
  INVX1 U629 ( .A(n522), .Y(n523) );
  AND2X2 U630 ( .A(\mem<19><13> ), .B(n2302), .Y(n524) );
  INVX1 U631 ( .A(n524), .Y(n525) );
  AND2X2 U632 ( .A(\mem<19><14> ), .B(n2302), .Y(n526) );
  INVX1 U633 ( .A(n526), .Y(n527) );
  AND2X2 U634 ( .A(\mem<19><15> ), .B(n2302), .Y(n528) );
  INVX1 U635 ( .A(n528), .Y(n529) );
  AND2X2 U636 ( .A(\mem<18><0> ), .B(n61), .Y(n530) );
  INVX1 U637 ( .A(n530), .Y(n531) );
  AND2X2 U638 ( .A(\mem<18><1> ), .B(n61), .Y(n532) );
  INVX1 U639 ( .A(n532), .Y(n533) );
  AND2X2 U640 ( .A(\mem<18><2> ), .B(n61), .Y(n534) );
  INVX1 U641 ( .A(n534), .Y(n535) );
  AND2X2 U642 ( .A(\mem<18><3> ), .B(n61), .Y(n536) );
  INVX1 U643 ( .A(n536), .Y(n537) );
  AND2X2 U644 ( .A(\mem<18><4> ), .B(n61), .Y(n538) );
  INVX1 U645 ( .A(n538), .Y(n539) );
  AND2X2 U646 ( .A(\mem<18><5> ), .B(n61), .Y(n540) );
  INVX1 U647 ( .A(n540), .Y(n541) );
  AND2X2 U648 ( .A(\mem<18><6> ), .B(n61), .Y(n542) );
  INVX1 U649 ( .A(n542), .Y(n543) );
  AND2X2 U650 ( .A(\mem<18><7> ), .B(n61), .Y(n544) );
  INVX1 U651 ( .A(n544), .Y(n545) );
  AND2X2 U652 ( .A(\mem<18><8> ), .B(n61), .Y(n546) );
  INVX1 U653 ( .A(n546), .Y(n547) );
  AND2X2 U654 ( .A(\mem<18><9> ), .B(n61), .Y(n548) );
  INVX1 U655 ( .A(n548), .Y(n549) );
  AND2X2 U656 ( .A(\mem<18><10> ), .B(n61), .Y(n550) );
  INVX1 U657 ( .A(n550), .Y(n551) );
  AND2X2 U658 ( .A(\mem<18><11> ), .B(n61), .Y(n552) );
  INVX1 U659 ( .A(n552), .Y(n553) );
  AND2X2 U660 ( .A(\mem<18><12> ), .B(n61), .Y(n554) );
  INVX1 U661 ( .A(n554), .Y(n555) );
  AND2X2 U662 ( .A(\mem<18><13> ), .B(n61), .Y(n556) );
  INVX1 U663 ( .A(n556), .Y(n557) );
  AND2X2 U664 ( .A(\mem<18><14> ), .B(n61), .Y(n558) );
  INVX1 U665 ( .A(n558), .Y(n559) );
  AND2X2 U666 ( .A(\mem<18><15> ), .B(n61), .Y(n560) );
  INVX1 U667 ( .A(n560), .Y(n561) );
  AND2X2 U668 ( .A(\mem<17><0> ), .B(n64), .Y(n562) );
  INVX1 U669 ( .A(n562), .Y(n563) );
  AND2X2 U670 ( .A(\mem<17><1> ), .B(n64), .Y(n564) );
  INVX1 U671 ( .A(n564), .Y(n565) );
  AND2X2 U672 ( .A(\mem<17><2> ), .B(n64), .Y(n566) );
  INVX1 U673 ( .A(n566), .Y(n567) );
  AND2X2 U674 ( .A(\mem<17><3> ), .B(n64), .Y(n568) );
  INVX1 U675 ( .A(n568), .Y(n569) );
  AND2X2 U676 ( .A(\mem<17><4> ), .B(n64), .Y(n570) );
  INVX1 U677 ( .A(n570), .Y(n571) );
  AND2X2 U678 ( .A(\mem<17><5> ), .B(n64), .Y(n572) );
  INVX1 U679 ( .A(n572), .Y(n573) );
  AND2X2 U680 ( .A(\mem<17><6> ), .B(n64), .Y(n574) );
  INVX1 U681 ( .A(n574), .Y(n575) );
  AND2X2 U682 ( .A(\mem<17><7> ), .B(n64), .Y(n576) );
  INVX1 U683 ( .A(n576), .Y(n577) );
  AND2X2 U684 ( .A(\mem<17><8> ), .B(n63), .Y(n578) );
  INVX1 U685 ( .A(n578), .Y(n579) );
  AND2X2 U686 ( .A(\mem<17><9> ), .B(n63), .Y(n580) );
  INVX1 U687 ( .A(n580), .Y(n581) );
  AND2X2 U688 ( .A(\mem<17><10> ), .B(n63), .Y(n582) );
  INVX1 U689 ( .A(n582), .Y(n583) );
  AND2X2 U690 ( .A(\mem<17><11> ), .B(n63), .Y(n584) );
  INVX1 U691 ( .A(n584), .Y(n585) );
  AND2X2 U692 ( .A(\mem<17><12> ), .B(n63), .Y(n586) );
  INVX1 U693 ( .A(n586), .Y(n587) );
  AND2X2 U694 ( .A(\mem<17><13> ), .B(n63), .Y(n588) );
  INVX1 U695 ( .A(n588), .Y(n589) );
  AND2X2 U696 ( .A(\mem<17><14> ), .B(n63), .Y(n590) );
  INVX1 U697 ( .A(n590), .Y(n591) );
  AND2X2 U698 ( .A(\mem<17><15> ), .B(n63), .Y(n592) );
  INVX1 U699 ( .A(n592), .Y(n593) );
  AND2X2 U700 ( .A(\mem<16><0> ), .B(n66), .Y(n594) );
  INVX1 U701 ( .A(n594), .Y(n595) );
  AND2X2 U702 ( .A(\mem<16><1> ), .B(n66), .Y(n596) );
  INVX1 U703 ( .A(n596), .Y(n597) );
  AND2X2 U704 ( .A(\mem<16><2> ), .B(n66), .Y(n598) );
  INVX1 U705 ( .A(n598), .Y(n599) );
  AND2X2 U706 ( .A(\mem<16><3> ), .B(n66), .Y(n600) );
  INVX1 U707 ( .A(n600), .Y(n601) );
  AND2X2 U708 ( .A(\mem<16><4> ), .B(n66), .Y(n602) );
  INVX1 U709 ( .A(n602), .Y(n603) );
  AND2X2 U710 ( .A(\mem<16><5> ), .B(n66), .Y(n604) );
  INVX1 U711 ( .A(n604), .Y(n605) );
  AND2X2 U712 ( .A(\mem<16><6> ), .B(n66), .Y(n606) );
  INVX1 U713 ( .A(n606), .Y(n607) );
  AND2X2 U714 ( .A(\mem<16><7> ), .B(n66), .Y(n608) );
  INVX1 U715 ( .A(n608), .Y(n609) );
  AND2X2 U716 ( .A(\mem<16><8> ), .B(n67), .Y(n610) );
  INVX1 U717 ( .A(n610), .Y(n611) );
  AND2X2 U718 ( .A(\mem<16><9> ), .B(n67), .Y(n612) );
  INVX1 U719 ( .A(n612), .Y(n613) );
  AND2X2 U720 ( .A(\mem<16><10> ), .B(n67), .Y(n614) );
  INVX1 U721 ( .A(n614), .Y(n615) );
  AND2X2 U722 ( .A(\mem<16><11> ), .B(n67), .Y(n616) );
  INVX1 U723 ( .A(n616), .Y(n617) );
  AND2X2 U724 ( .A(\mem<16><12> ), .B(n67), .Y(n618) );
  INVX1 U725 ( .A(n618), .Y(n619) );
  AND2X2 U726 ( .A(\mem<16><13> ), .B(n67), .Y(n620) );
  INVX1 U727 ( .A(n620), .Y(n621) );
  AND2X2 U728 ( .A(\mem<16><14> ), .B(n67), .Y(n622) );
  INVX1 U729 ( .A(n622), .Y(n623) );
  AND2X2 U730 ( .A(\mem<16><15> ), .B(n67), .Y(n624) );
  INVX1 U731 ( .A(n624), .Y(n625) );
  AND2X2 U732 ( .A(\mem<15><0> ), .B(n70), .Y(n626) );
  INVX1 U733 ( .A(n626), .Y(n627) );
  AND2X2 U734 ( .A(\mem<15><1> ), .B(n70), .Y(n628) );
  INVX1 U735 ( .A(n628), .Y(n629) );
  AND2X2 U736 ( .A(\mem<15><2> ), .B(n70), .Y(n630) );
  INVX1 U737 ( .A(n630), .Y(n631) );
  AND2X2 U738 ( .A(\mem<15><3> ), .B(n70), .Y(n632) );
  INVX1 U739 ( .A(n632), .Y(n633) );
  AND2X2 U740 ( .A(\mem<15><4> ), .B(n70), .Y(n634) );
  INVX1 U741 ( .A(n634), .Y(n635) );
  AND2X2 U742 ( .A(\mem<15><5> ), .B(n70), .Y(n636) );
  INVX1 U743 ( .A(n636), .Y(n637) );
  AND2X2 U744 ( .A(\mem<15><6> ), .B(n70), .Y(n638) );
  INVX1 U745 ( .A(n638), .Y(n639) );
  AND2X2 U746 ( .A(\mem<15><7> ), .B(n70), .Y(n640) );
  INVX1 U747 ( .A(n640), .Y(n641) );
  AND2X2 U748 ( .A(\mem<15><8> ), .B(n69), .Y(n642) );
  INVX1 U749 ( .A(n642), .Y(n643) );
  AND2X2 U750 ( .A(\mem<15><9> ), .B(n69), .Y(n644) );
  INVX1 U751 ( .A(n644), .Y(n645) );
  AND2X2 U752 ( .A(\mem<15><10> ), .B(n69), .Y(n646) );
  INVX1 U753 ( .A(n646), .Y(n647) );
  AND2X2 U754 ( .A(\mem<15><11> ), .B(n69), .Y(n648) );
  INVX1 U755 ( .A(n648), .Y(n649) );
  AND2X2 U756 ( .A(\mem<15><12> ), .B(n69), .Y(n650) );
  INVX1 U757 ( .A(n650), .Y(n1163) );
  AND2X2 U758 ( .A(\mem<15><13> ), .B(n69), .Y(n1164) );
  INVX1 U759 ( .A(n1164), .Y(n1165) );
  AND2X2 U760 ( .A(\mem<15><14> ), .B(n69), .Y(n1166) );
  INVX1 U761 ( .A(n1166), .Y(n1167) );
  AND2X2 U762 ( .A(\mem<15><15> ), .B(n69), .Y(n1168) );
  INVX1 U763 ( .A(n1168), .Y(n1169) );
  AND2X2 U764 ( .A(\mem<14><0> ), .B(n73), .Y(n1170) );
  INVX1 U765 ( .A(n1170), .Y(n1171) );
  AND2X2 U766 ( .A(\mem<14><1> ), .B(n73), .Y(n1172) );
  INVX1 U767 ( .A(n1172), .Y(n1173) );
  AND2X2 U768 ( .A(\mem<14><2> ), .B(n73), .Y(n1174) );
  INVX1 U769 ( .A(n1174), .Y(n1175) );
  AND2X2 U770 ( .A(\mem<14><3> ), .B(n73), .Y(n1176) );
  INVX1 U771 ( .A(n1176), .Y(n1177) );
  AND2X2 U772 ( .A(\mem<14><4> ), .B(n73), .Y(n1178) );
  INVX1 U773 ( .A(n1178), .Y(n1179) );
  AND2X2 U774 ( .A(\mem<14><5> ), .B(n73), .Y(n1180) );
  INVX1 U775 ( .A(n1180), .Y(n1181) );
  AND2X2 U776 ( .A(\mem<14><6> ), .B(n73), .Y(n1182) );
  INVX1 U777 ( .A(n1182), .Y(n1183) );
  AND2X2 U778 ( .A(\mem<14><7> ), .B(n73), .Y(n1184) );
  INVX1 U779 ( .A(n1184), .Y(n1185) );
  AND2X2 U780 ( .A(\mem<14><8> ), .B(n72), .Y(n1186) );
  INVX1 U781 ( .A(n1186), .Y(n1187) );
  AND2X2 U782 ( .A(\mem<14><9> ), .B(n72), .Y(n1188) );
  INVX1 U783 ( .A(n1188), .Y(n1189) );
  AND2X2 U784 ( .A(\mem<14><10> ), .B(n72), .Y(n1190) );
  INVX1 U785 ( .A(n1190), .Y(n1191) );
  AND2X2 U786 ( .A(\mem<14><11> ), .B(n72), .Y(n1192) );
  INVX1 U787 ( .A(n1192), .Y(n1193) );
  AND2X2 U788 ( .A(\mem<14><12> ), .B(n72), .Y(n1194) );
  INVX1 U789 ( .A(n1194), .Y(n1195) );
  AND2X2 U790 ( .A(\mem<14><13> ), .B(n72), .Y(n1196) );
  INVX1 U791 ( .A(n1196), .Y(n1197) );
  AND2X2 U792 ( .A(\mem<14><14> ), .B(n72), .Y(n1198) );
  INVX1 U793 ( .A(n1198), .Y(n1199) );
  AND2X2 U794 ( .A(\mem<14><15> ), .B(n72), .Y(n1200) );
  INVX1 U795 ( .A(n1200), .Y(n1201) );
  AND2X2 U796 ( .A(\mem<13><0> ), .B(n76), .Y(n1202) );
  INVX1 U797 ( .A(n1202), .Y(n1203) );
  AND2X2 U798 ( .A(\mem<13><1> ), .B(n76), .Y(n1204) );
  INVX1 U799 ( .A(n1204), .Y(n1205) );
  AND2X2 U800 ( .A(\mem<13><2> ), .B(n76), .Y(n1206) );
  INVX1 U801 ( .A(n1206), .Y(n1207) );
  AND2X2 U802 ( .A(\mem<13><3> ), .B(n76), .Y(n1208) );
  INVX1 U803 ( .A(n1208), .Y(n1209) );
  AND2X2 U804 ( .A(\mem<13><4> ), .B(n76), .Y(n1210) );
  INVX1 U805 ( .A(n1210), .Y(n1211) );
  AND2X2 U806 ( .A(\mem<13><5> ), .B(n76), .Y(n1212) );
  INVX1 U807 ( .A(n1212), .Y(n1213) );
  AND2X2 U808 ( .A(\mem<13><6> ), .B(n76), .Y(n1214) );
  INVX1 U809 ( .A(n1214), .Y(n1215) );
  AND2X2 U810 ( .A(\mem<13><7> ), .B(n76), .Y(n1216) );
  INVX1 U811 ( .A(n1216), .Y(n1217) );
  AND2X2 U812 ( .A(\mem<13><8> ), .B(n75), .Y(n1218) );
  INVX1 U813 ( .A(n1218), .Y(n1219) );
  AND2X2 U814 ( .A(\mem<13><9> ), .B(n75), .Y(n1220) );
  INVX1 U815 ( .A(n1220), .Y(n1221) );
  AND2X2 U816 ( .A(\mem<13><10> ), .B(n75), .Y(n1222) );
  INVX1 U817 ( .A(n1222), .Y(n1223) );
  AND2X2 U818 ( .A(\mem<13><11> ), .B(n75), .Y(n1224) );
  INVX1 U819 ( .A(n1224), .Y(n1225) );
  AND2X2 U820 ( .A(\mem<13><12> ), .B(n75), .Y(n1226) );
  INVX1 U821 ( .A(n1226), .Y(n1227) );
  AND2X2 U822 ( .A(\mem<13><13> ), .B(n75), .Y(n1228) );
  INVX1 U823 ( .A(n1228), .Y(n1229) );
  AND2X2 U824 ( .A(\mem<13><14> ), .B(n75), .Y(n1230) );
  INVX1 U825 ( .A(n1230), .Y(n1231) );
  AND2X2 U826 ( .A(\mem<13><15> ), .B(n75), .Y(n1232) );
  INVX1 U827 ( .A(n1232), .Y(n1233) );
  AND2X2 U828 ( .A(\mem<12><0> ), .B(n79), .Y(n1234) );
  INVX1 U829 ( .A(n1234), .Y(n1235) );
  AND2X2 U830 ( .A(\mem<12><1> ), .B(n79), .Y(n1236) );
  INVX1 U831 ( .A(n1236), .Y(n1237) );
  AND2X2 U832 ( .A(\mem<12><2> ), .B(n79), .Y(n1238) );
  INVX1 U833 ( .A(n1238), .Y(n1239) );
  AND2X2 U834 ( .A(\mem<12><3> ), .B(n79), .Y(n1240) );
  INVX1 U835 ( .A(n1240), .Y(n1241) );
  AND2X2 U836 ( .A(\mem<12><4> ), .B(n79), .Y(n1242) );
  INVX1 U837 ( .A(n1242), .Y(n1243) );
  AND2X2 U838 ( .A(\mem<12><5> ), .B(n79), .Y(n1244) );
  INVX1 U839 ( .A(n1244), .Y(n1245) );
  AND2X2 U840 ( .A(\mem<12><6> ), .B(n79), .Y(n1246) );
  INVX1 U841 ( .A(n1246), .Y(n1247) );
  AND2X2 U842 ( .A(\mem<12><7> ), .B(n79), .Y(n1248) );
  INVX1 U843 ( .A(n1248), .Y(n1249) );
  AND2X2 U844 ( .A(\mem<12><8> ), .B(n78), .Y(n1250) );
  INVX1 U845 ( .A(n1250), .Y(n1251) );
  AND2X2 U846 ( .A(\mem<12><9> ), .B(n78), .Y(n1252) );
  INVX1 U847 ( .A(n1252), .Y(n1253) );
  AND2X2 U848 ( .A(\mem<12><10> ), .B(n78), .Y(n1254) );
  INVX1 U849 ( .A(n1254), .Y(n1255) );
  AND2X2 U850 ( .A(\mem<12><11> ), .B(n78), .Y(n1256) );
  INVX1 U851 ( .A(n1256), .Y(n1257) );
  AND2X2 U852 ( .A(\mem<12><12> ), .B(n78), .Y(n1258) );
  INVX1 U853 ( .A(n1258), .Y(n1259) );
  AND2X2 U854 ( .A(\mem<12><13> ), .B(n78), .Y(n1260) );
  INVX1 U855 ( .A(n1260), .Y(n1261) );
  AND2X2 U856 ( .A(\mem<12><14> ), .B(n78), .Y(n1262) );
  INVX1 U857 ( .A(n1262), .Y(n1263) );
  AND2X2 U858 ( .A(\mem<12><15> ), .B(n78), .Y(n1264) );
  INVX1 U859 ( .A(n1264), .Y(n1265) );
  AND2X2 U860 ( .A(\mem<11><0> ), .B(n82), .Y(n1266) );
  INVX1 U861 ( .A(n1266), .Y(n1267) );
  AND2X2 U862 ( .A(\mem<11><1> ), .B(n82), .Y(n1268) );
  INVX1 U863 ( .A(n1268), .Y(n1269) );
  AND2X2 U864 ( .A(\mem<11><2> ), .B(n82), .Y(n1270) );
  INVX1 U865 ( .A(n1270), .Y(n1271) );
  AND2X2 U866 ( .A(\mem<11><3> ), .B(n82), .Y(n1272) );
  INVX1 U867 ( .A(n1272), .Y(n1273) );
  AND2X2 U868 ( .A(\mem<11><4> ), .B(n82), .Y(n1274) );
  INVX1 U869 ( .A(n1274), .Y(n1275) );
  AND2X2 U870 ( .A(\mem<11><5> ), .B(n82), .Y(n1276) );
  INVX1 U871 ( .A(n1276), .Y(n1277) );
  AND2X2 U872 ( .A(\mem<11><6> ), .B(n82), .Y(n1278) );
  INVX1 U873 ( .A(n1278), .Y(n1279) );
  AND2X2 U874 ( .A(\mem<11><7> ), .B(n82), .Y(n1280) );
  INVX1 U875 ( .A(n1280), .Y(n1281) );
  AND2X2 U876 ( .A(\mem<11><8> ), .B(n81), .Y(n1282) );
  INVX1 U877 ( .A(n1282), .Y(n1283) );
  AND2X2 U878 ( .A(\mem<11><9> ), .B(n81), .Y(n1284) );
  INVX1 U879 ( .A(n1284), .Y(n1285) );
  AND2X2 U880 ( .A(\mem<11><10> ), .B(n81), .Y(n1286) );
  INVX1 U881 ( .A(n1286), .Y(n1287) );
  AND2X2 U882 ( .A(\mem<11><11> ), .B(n81), .Y(n1288) );
  INVX1 U883 ( .A(n1288), .Y(n1289) );
  AND2X2 U884 ( .A(\mem<11><12> ), .B(n81), .Y(n1290) );
  INVX1 U885 ( .A(n1290), .Y(n1291) );
  AND2X2 U886 ( .A(\mem<11><13> ), .B(n81), .Y(n1292) );
  INVX1 U887 ( .A(n1292), .Y(n1293) );
  AND2X2 U888 ( .A(\mem<11><14> ), .B(n81), .Y(n1294) );
  INVX1 U889 ( .A(n1294), .Y(n1295) );
  AND2X2 U890 ( .A(\mem<11><15> ), .B(n81), .Y(n1296) );
  INVX1 U891 ( .A(n1296), .Y(n1297) );
  AND2X2 U892 ( .A(\mem<10><0> ), .B(n85), .Y(n1298) );
  INVX1 U893 ( .A(n1298), .Y(n1299) );
  AND2X2 U894 ( .A(\mem<10><1> ), .B(n85), .Y(n1300) );
  INVX1 U895 ( .A(n1300), .Y(n1301) );
  AND2X2 U896 ( .A(\mem<10><2> ), .B(n85), .Y(n1302) );
  INVX1 U897 ( .A(n1302), .Y(n1303) );
  AND2X2 U898 ( .A(\mem<10><3> ), .B(n85), .Y(n1304) );
  INVX1 U899 ( .A(n1304), .Y(n1305) );
  AND2X2 U900 ( .A(\mem<10><4> ), .B(n85), .Y(n1306) );
  INVX1 U901 ( .A(n1306), .Y(n1307) );
  AND2X2 U902 ( .A(\mem<10><5> ), .B(n85), .Y(n1308) );
  INVX1 U903 ( .A(n1308), .Y(n1309) );
  AND2X2 U904 ( .A(\mem<10><6> ), .B(n85), .Y(n1310) );
  INVX1 U905 ( .A(n1310), .Y(n1311) );
  AND2X2 U906 ( .A(\mem<10><7> ), .B(n85), .Y(n1312) );
  INVX1 U907 ( .A(n1312), .Y(n1313) );
  AND2X2 U908 ( .A(\mem<10><8> ), .B(n84), .Y(n1314) );
  INVX1 U909 ( .A(n1314), .Y(n1315) );
  AND2X2 U910 ( .A(\mem<10><9> ), .B(n84), .Y(n1316) );
  INVX1 U911 ( .A(n1316), .Y(n1317) );
  AND2X2 U912 ( .A(\mem<10><10> ), .B(n84), .Y(n1318) );
  INVX1 U913 ( .A(n1318), .Y(n1319) );
  AND2X2 U914 ( .A(\mem<10><11> ), .B(n84), .Y(n1320) );
  INVX1 U915 ( .A(n1320), .Y(n1321) );
  AND2X2 U916 ( .A(\mem<10><12> ), .B(n84), .Y(n1322) );
  INVX1 U917 ( .A(n1322), .Y(n1323) );
  AND2X2 U918 ( .A(\mem<10><13> ), .B(n84), .Y(n1324) );
  INVX1 U919 ( .A(n1324), .Y(n1325) );
  AND2X2 U920 ( .A(\mem<10><14> ), .B(n84), .Y(n1326) );
  INVX1 U921 ( .A(n1326), .Y(n1327) );
  AND2X2 U922 ( .A(\mem<10><15> ), .B(n84), .Y(n1328) );
  INVX1 U923 ( .A(n1328), .Y(n1329) );
  AND2X2 U924 ( .A(\mem<9><0> ), .B(n88), .Y(n1330) );
  INVX1 U925 ( .A(n1330), .Y(n1331) );
  AND2X2 U926 ( .A(\mem<9><1> ), .B(n88), .Y(n1332) );
  INVX1 U927 ( .A(n1332), .Y(n1333) );
  AND2X2 U928 ( .A(\mem<9><2> ), .B(n88), .Y(n1334) );
  INVX1 U929 ( .A(n1334), .Y(n1335) );
  AND2X2 U930 ( .A(\mem<9><3> ), .B(n88), .Y(n1336) );
  INVX1 U931 ( .A(n1336), .Y(n1337) );
  AND2X2 U932 ( .A(\mem<9><4> ), .B(n88), .Y(n1338) );
  INVX1 U933 ( .A(n1338), .Y(n1339) );
  AND2X2 U934 ( .A(\mem<9><5> ), .B(n88), .Y(n1340) );
  INVX1 U935 ( .A(n1340), .Y(n1341) );
  AND2X2 U936 ( .A(\mem<9><6> ), .B(n88), .Y(n1342) );
  INVX1 U937 ( .A(n1342), .Y(n1343) );
  AND2X2 U938 ( .A(\mem<9><7> ), .B(n88), .Y(n1344) );
  INVX1 U939 ( .A(n1344), .Y(n1345) );
  AND2X2 U940 ( .A(\mem<9><8> ), .B(n87), .Y(n1346) );
  INVX1 U941 ( .A(n1346), .Y(n1347) );
  AND2X2 U942 ( .A(\mem<9><9> ), .B(n87), .Y(n1348) );
  INVX1 U943 ( .A(n1348), .Y(n1349) );
  AND2X2 U944 ( .A(\mem<9><10> ), .B(n87), .Y(n1350) );
  INVX1 U945 ( .A(n1350), .Y(n1351) );
  AND2X2 U946 ( .A(\mem<9><11> ), .B(n87), .Y(n1352) );
  INVX1 U947 ( .A(n1352), .Y(n1353) );
  AND2X2 U948 ( .A(\mem<9><12> ), .B(n87), .Y(n1354) );
  INVX1 U949 ( .A(n1354), .Y(n1355) );
  AND2X2 U950 ( .A(\mem<9><13> ), .B(n87), .Y(n1356) );
  INVX1 U951 ( .A(n1356), .Y(n1357) );
  AND2X2 U952 ( .A(\mem<9><14> ), .B(n87), .Y(n1358) );
  INVX1 U953 ( .A(n1358), .Y(n1359) );
  AND2X2 U954 ( .A(\mem<9><15> ), .B(n87), .Y(n1360) );
  INVX1 U955 ( .A(n1360), .Y(n1361) );
  AND2X2 U956 ( .A(\mem<8><0> ), .B(n25), .Y(n1362) );
  INVX1 U957 ( .A(n1362), .Y(n1363) );
  AND2X2 U958 ( .A(\mem<8><1> ), .B(n25), .Y(n1364) );
  INVX1 U959 ( .A(n1364), .Y(n1365) );
  AND2X2 U960 ( .A(\mem<8><2> ), .B(n25), .Y(n1366) );
  INVX1 U961 ( .A(n1366), .Y(n1367) );
  AND2X2 U962 ( .A(\mem<8><3> ), .B(n25), .Y(n1368) );
  INVX1 U963 ( .A(n1368), .Y(n1369) );
  AND2X2 U964 ( .A(\mem<8><4> ), .B(n25), .Y(n1370) );
  INVX1 U965 ( .A(n1370), .Y(n1371) );
  AND2X2 U966 ( .A(\mem<8><5> ), .B(n25), .Y(n1372) );
  INVX1 U967 ( .A(n1372), .Y(n1373) );
  AND2X2 U968 ( .A(\mem<8><6> ), .B(n25), .Y(n1374) );
  INVX1 U969 ( .A(n1374), .Y(n1375) );
  AND2X2 U970 ( .A(\mem<8><7> ), .B(n25), .Y(n1376) );
  INVX1 U971 ( .A(n1376), .Y(n1377) );
  AND2X2 U972 ( .A(\mem<8><8> ), .B(n25), .Y(n1378) );
  INVX1 U973 ( .A(n1378), .Y(n1379) );
  AND2X2 U974 ( .A(\mem<8><9> ), .B(n25), .Y(n1380) );
  INVX1 U975 ( .A(n1380), .Y(n1381) );
  AND2X2 U976 ( .A(\mem<8><10> ), .B(n25), .Y(n1382) );
  INVX1 U977 ( .A(n1382), .Y(n1383) );
  AND2X2 U978 ( .A(\mem<8><11> ), .B(n25), .Y(n1384) );
  INVX1 U979 ( .A(n1384), .Y(n1385) );
  AND2X2 U980 ( .A(\mem<8><12> ), .B(n25), .Y(n1386) );
  INVX1 U981 ( .A(n1386), .Y(n1387) );
  AND2X2 U982 ( .A(\mem<8><13> ), .B(n25), .Y(n1388) );
  INVX1 U983 ( .A(n1388), .Y(n1389) );
  AND2X2 U984 ( .A(\mem<8><14> ), .B(n25), .Y(n1390) );
  INVX1 U985 ( .A(n1390), .Y(n1391) );
  AND2X2 U986 ( .A(\mem<8><15> ), .B(n25), .Y(n1392) );
  INVX1 U987 ( .A(n1392), .Y(n1393) );
  AND2X2 U988 ( .A(\mem<7><0> ), .B(n90), .Y(n1394) );
  INVX1 U989 ( .A(n1394), .Y(n1395) );
  AND2X2 U990 ( .A(\mem<7><1> ), .B(n90), .Y(n1396) );
  INVX1 U991 ( .A(n1396), .Y(n1397) );
  AND2X2 U992 ( .A(\mem<7><2> ), .B(n90), .Y(n1398) );
  INVX1 U993 ( .A(n1398), .Y(n1399) );
  AND2X2 U994 ( .A(\mem<7><3> ), .B(n90), .Y(n1400) );
  INVX1 U995 ( .A(n1400), .Y(n1401) );
  AND2X2 U996 ( .A(\mem<7><4> ), .B(n90), .Y(n1402) );
  INVX1 U997 ( .A(n1402), .Y(n1403) );
  AND2X2 U998 ( .A(\mem<7><5> ), .B(n90), .Y(n1404) );
  INVX1 U999 ( .A(n1404), .Y(n1405) );
  AND2X2 U1000 ( .A(\mem<7><6> ), .B(n90), .Y(n1406) );
  INVX1 U1001 ( .A(n1406), .Y(n1407) );
  AND2X2 U1002 ( .A(\mem<7><7> ), .B(n90), .Y(n1408) );
  INVX1 U1003 ( .A(n1408), .Y(n1409) );
  AND2X2 U1004 ( .A(\mem<7><8> ), .B(n90), .Y(n1410) );
  INVX1 U1005 ( .A(n1410), .Y(n1411) );
  AND2X2 U1006 ( .A(\mem<7><9> ), .B(n90), .Y(n1412) );
  INVX1 U1007 ( .A(n1412), .Y(n1413) );
  AND2X2 U1008 ( .A(\mem<7><10> ), .B(n90), .Y(n1414) );
  INVX1 U1009 ( .A(n1414), .Y(n1415) );
  AND2X2 U1010 ( .A(\mem<7><11> ), .B(n90), .Y(n1416) );
  INVX1 U1011 ( .A(n1416), .Y(n1417) );
  AND2X2 U1012 ( .A(\mem<7><12> ), .B(n90), .Y(n1418) );
  INVX1 U1013 ( .A(n1418), .Y(n1419) );
  AND2X2 U1014 ( .A(\mem<7><13> ), .B(n90), .Y(n1420) );
  INVX1 U1015 ( .A(n1420), .Y(n1421) );
  AND2X2 U1016 ( .A(\mem<7><14> ), .B(n90), .Y(n1422) );
  INVX1 U1017 ( .A(n1422), .Y(n1423) );
  AND2X2 U1018 ( .A(\mem<7><15> ), .B(n90), .Y(n1424) );
  INVX1 U1019 ( .A(n1424), .Y(n1425) );
  AND2X2 U1020 ( .A(\mem<6><0> ), .B(n93), .Y(n1426) );
  INVX1 U1021 ( .A(n1426), .Y(n1427) );
  AND2X2 U1022 ( .A(\mem<6><1> ), .B(n93), .Y(n1428) );
  INVX1 U1023 ( .A(n1428), .Y(n1429) );
  AND2X2 U1024 ( .A(\mem<6><2> ), .B(n93), .Y(n1430) );
  INVX1 U1025 ( .A(n1430), .Y(n1431) );
  AND2X2 U1026 ( .A(\mem<6><3> ), .B(n93), .Y(n1432) );
  INVX1 U1027 ( .A(n1432), .Y(n1433) );
  AND2X2 U1028 ( .A(\mem<6><4> ), .B(n93), .Y(n1434) );
  INVX1 U1029 ( .A(n1434), .Y(n1435) );
  AND2X2 U1030 ( .A(\mem<6><5> ), .B(n93), .Y(n1436) );
  INVX1 U1031 ( .A(n1436), .Y(n1437) );
  AND2X2 U1032 ( .A(\mem<6><6> ), .B(n93), .Y(n1438) );
  INVX1 U1033 ( .A(n1438), .Y(n1439) );
  AND2X2 U1034 ( .A(\mem<6><7> ), .B(n93), .Y(n1440) );
  INVX1 U1035 ( .A(n1440), .Y(n1441) );
  AND2X2 U1036 ( .A(\mem<6><8> ), .B(n92), .Y(n1442) );
  INVX1 U1037 ( .A(n1442), .Y(n1443) );
  AND2X2 U1038 ( .A(\mem<6><9> ), .B(n92), .Y(n1444) );
  INVX1 U1039 ( .A(n1444), .Y(n1445) );
  AND2X2 U1040 ( .A(\mem<6><10> ), .B(n92), .Y(n1446) );
  INVX1 U1041 ( .A(n1446), .Y(n1447) );
  AND2X2 U1042 ( .A(\mem<6><11> ), .B(n92), .Y(n1448) );
  INVX1 U1043 ( .A(n1448), .Y(n1449) );
  AND2X2 U1044 ( .A(\mem<6><12> ), .B(n92), .Y(n1450) );
  INVX1 U1045 ( .A(n1450), .Y(n1451) );
  AND2X2 U1046 ( .A(\mem<6><13> ), .B(n92), .Y(n1452) );
  INVX1 U1047 ( .A(n1452), .Y(n1453) );
  AND2X2 U1048 ( .A(\mem<6><14> ), .B(n92), .Y(n1454) );
  INVX1 U1049 ( .A(n1454), .Y(n1455) );
  AND2X2 U1050 ( .A(\mem<6><15> ), .B(n92), .Y(n1456) );
  INVX1 U1051 ( .A(n1456), .Y(n1457) );
  AND2X2 U1052 ( .A(\mem<5><0> ), .B(n96), .Y(n1458) );
  INVX1 U1053 ( .A(n1458), .Y(n1459) );
  AND2X2 U1054 ( .A(\mem<5><1> ), .B(n96), .Y(n1460) );
  INVX1 U1055 ( .A(n1460), .Y(n1461) );
  AND2X2 U1056 ( .A(\mem<5><2> ), .B(n96), .Y(n1462) );
  INVX1 U1057 ( .A(n1462), .Y(n1463) );
  AND2X2 U1058 ( .A(\mem<5><3> ), .B(n96), .Y(n1464) );
  INVX1 U1059 ( .A(n1464), .Y(n1465) );
  AND2X2 U1060 ( .A(\mem<5><4> ), .B(n96), .Y(n1466) );
  INVX1 U1061 ( .A(n1466), .Y(n1467) );
  AND2X2 U1062 ( .A(\mem<5><5> ), .B(n96), .Y(n1468) );
  INVX1 U1063 ( .A(n1468), .Y(n1469) );
  AND2X2 U1064 ( .A(\mem<5><6> ), .B(n96), .Y(n1470) );
  INVX1 U1065 ( .A(n1470), .Y(n1471) );
  AND2X2 U1066 ( .A(\mem<5><7> ), .B(n96), .Y(n1472) );
  INVX1 U1067 ( .A(n1472), .Y(n1473) );
  AND2X2 U1068 ( .A(\mem<5><8> ), .B(n95), .Y(n1474) );
  INVX1 U1069 ( .A(n1474), .Y(n1475) );
  AND2X2 U1070 ( .A(\mem<5><9> ), .B(n95), .Y(n1476) );
  INVX1 U1071 ( .A(n1476), .Y(n1477) );
  AND2X2 U1072 ( .A(\mem<5><10> ), .B(n95), .Y(n1478) );
  INVX1 U1073 ( .A(n1478), .Y(n1479) );
  AND2X2 U1074 ( .A(\mem<5><11> ), .B(n95), .Y(n1480) );
  INVX1 U1075 ( .A(n1480), .Y(n1481) );
  AND2X2 U1076 ( .A(\mem<5><12> ), .B(n95), .Y(n1482) );
  INVX1 U1077 ( .A(n1482), .Y(n1483) );
  AND2X2 U1078 ( .A(\mem<5><13> ), .B(n95), .Y(n1484) );
  INVX1 U1079 ( .A(n1484), .Y(n1485) );
  AND2X2 U1080 ( .A(\mem<5><14> ), .B(n95), .Y(n1486) );
  INVX1 U1081 ( .A(n1486), .Y(n1487) );
  AND2X2 U1082 ( .A(\mem<5><15> ), .B(n95), .Y(n1488) );
  INVX1 U1083 ( .A(n1488), .Y(n1489) );
  AND2X2 U1084 ( .A(\mem<4><0> ), .B(n99), .Y(n1490) );
  INVX1 U1085 ( .A(n1490), .Y(n1491) );
  AND2X2 U1086 ( .A(\mem<4><1> ), .B(n99), .Y(n1492) );
  INVX1 U1087 ( .A(n1492), .Y(n1493) );
  AND2X2 U1088 ( .A(\mem<4><2> ), .B(n99), .Y(n1494) );
  INVX1 U1089 ( .A(n1494), .Y(n1495) );
  AND2X2 U1090 ( .A(\mem<4><3> ), .B(n99), .Y(n1496) );
  INVX1 U1091 ( .A(n1496), .Y(n1497) );
  AND2X2 U1092 ( .A(\mem<4><4> ), .B(n99), .Y(n1498) );
  INVX1 U1093 ( .A(n1498), .Y(n1499) );
  AND2X2 U1094 ( .A(\mem<4><5> ), .B(n99), .Y(n1500) );
  INVX1 U1095 ( .A(n1500), .Y(n1501) );
  AND2X2 U1096 ( .A(\mem<4><6> ), .B(n99), .Y(n1502) );
  INVX1 U1097 ( .A(n1502), .Y(n1503) );
  AND2X2 U1098 ( .A(\mem<4><7> ), .B(n99), .Y(n1504) );
  INVX1 U1099 ( .A(n1504), .Y(n1505) );
  AND2X2 U1100 ( .A(\mem<4><8> ), .B(n98), .Y(n1506) );
  INVX1 U1101 ( .A(n1506), .Y(n1507) );
  AND2X2 U1102 ( .A(\mem<4><9> ), .B(n98), .Y(n1508) );
  INVX1 U1103 ( .A(n1508), .Y(n1509) );
  AND2X2 U1104 ( .A(\mem<4><10> ), .B(n98), .Y(n1510) );
  INVX1 U1105 ( .A(n1510), .Y(n1511) );
  AND2X2 U1106 ( .A(\mem<4><11> ), .B(n98), .Y(n1512) );
  INVX1 U1107 ( .A(n1512), .Y(n1513) );
  AND2X2 U1108 ( .A(\mem<4><12> ), .B(n98), .Y(n1514) );
  INVX1 U1109 ( .A(n1514), .Y(n1515) );
  AND2X2 U1110 ( .A(\mem<4><13> ), .B(n98), .Y(n1516) );
  INVX1 U1111 ( .A(n1516), .Y(n1517) );
  AND2X2 U1112 ( .A(\mem<4><14> ), .B(n98), .Y(n1518) );
  INVX1 U1113 ( .A(n1518), .Y(n1519) );
  AND2X2 U1114 ( .A(\mem<4><15> ), .B(n98), .Y(n1520) );
  INVX1 U1115 ( .A(n1520), .Y(n1521) );
  AND2X2 U1116 ( .A(\mem<3><0> ), .B(n102), .Y(n1522) );
  INVX1 U1117 ( .A(n1522), .Y(n1523) );
  AND2X2 U1118 ( .A(\mem<3><1> ), .B(n102), .Y(n1524) );
  INVX1 U1119 ( .A(n1524), .Y(n1525) );
  AND2X2 U1120 ( .A(\mem<3><2> ), .B(n102), .Y(n1526) );
  INVX1 U1121 ( .A(n1526), .Y(n1527) );
  AND2X2 U1122 ( .A(\mem<3><3> ), .B(n102), .Y(n1528) );
  INVX1 U1123 ( .A(n1528), .Y(n1529) );
  AND2X2 U1124 ( .A(\mem<3><4> ), .B(n102), .Y(n1530) );
  INVX1 U1125 ( .A(n1530), .Y(n1531) );
  AND2X2 U1126 ( .A(\mem<3><5> ), .B(n102), .Y(n1532) );
  INVX1 U1127 ( .A(n1532), .Y(n1533) );
  AND2X2 U1128 ( .A(\mem<3><6> ), .B(n102), .Y(n1534) );
  INVX1 U1129 ( .A(n1534), .Y(n1535) );
  AND2X2 U1130 ( .A(\mem<3><7> ), .B(n102), .Y(n1536) );
  INVX1 U1131 ( .A(n1536), .Y(n1537) );
  AND2X2 U1132 ( .A(\mem<3><8> ), .B(n101), .Y(n1538) );
  INVX1 U1133 ( .A(n1538), .Y(n1539) );
  AND2X2 U1134 ( .A(\mem<3><9> ), .B(n101), .Y(n1540) );
  INVX1 U1135 ( .A(n1540), .Y(n1541) );
  AND2X2 U1136 ( .A(\mem<3><10> ), .B(n101), .Y(n1542) );
  INVX1 U1137 ( .A(n1542), .Y(n1543) );
  AND2X2 U1138 ( .A(\mem<3><11> ), .B(n101), .Y(n1544) );
  INVX1 U1139 ( .A(n1544), .Y(n1545) );
  AND2X2 U1140 ( .A(\mem<3><12> ), .B(n101), .Y(n1546) );
  INVX1 U1141 ( .A(n1546), .Y(n1547) );
  AND2X2 U1142 ( .A(\mem<3><13> ), .B(n101), .Y(n1548) );
  INVX1 U1143 ( .A(n1548), .Y(n1549) );
  AND2X2 U1144 ( .A(\mem<3><14> ), .B(n101), .Y(n1550) );
  INVX1 U1145 ( .A(n1550), .Y(n1551) );
  AND2X2 U1146 ( .A(\mem<3><15> ), .B(n101), .Y(n1552) );
  INVX1 U1147 ( .A(n1552), .Y(n1553) );
  AND2X2 U1148 ( .A(\mem<2><0> ), .B(n105), .Y(n1554) );
  INVX1 U1149 ( .A(n1554), .Y(n1555) );
  AND2X2 U1150 ( .A(\mem<2><1> ), .B(n105), .Y(n1556) );
  INVX1 U1151 ( .A(n1556), .Y(n1557) );
  AND2X2 U1152 ( .A(\mem<2><2> ), .B(n105), .Y(n1558) );
  INVX1 U1153 ( .A(n1558), .Y(n1559) );
  AND2X2 U1154 ( .A(\mem<2><3> ), .B(n105), .Y(n1560) );
  INVX1 U1155 ( .A(n1560), .Y(n1561) );
  AND2X2 U1156 ( .A(\mem<2><4> ), .B(n105), .Y(n1562) );
  INVX1 U1157 ( .A(n1562), .Y(n1563) );
  AND2X2 U1158 ( .A(\mem<2><5> ), .B(n105), .Y(n1564) );
  INVX1 U1159 ( .A(n1564), .Y(n1565) );
  AND2X2 U1160 ( .A(\mem<2><6> ), .B(n105), .Y(n1566) );
  INVX1 U1161 ( .A(n1566), .Y(n1567) );
  AND2X2 U1162 ( .A(\mem<2><7> ), .B(n105), .Y(n1568) );
  INVX1 U1163 ( .A(n1568), .Y(n1569) );
  AND2X2 U1164 ( .A(\mem<2><8> ), .B(n104), .Y(n1570) );
  INVX1 U1165 ( .A(n1570), .Y(n1571) );
  AND2X2 U1166 ( .A(\mem<2><9> ), .B(n104), .Y(n1572) );
  INVX1 U1167 ( .A(n1572), .Y(n1573) );
  AND2X2 U1168 ( .A(\mem<2><10> ), .B(n104), .Y(n1574) );
  INVX1 U1169 ( .A(n1574), .Y(n1575) );
  AND2X2 U1170 ( .A(\mem<2><11> ), .B(n104), .Y(n1576) );
  INVX1 U1171 ( .A(n1576), .Y(n1577) );
  AND2X2 U1172 ( .A(\mem<2><12> ), .B(n104), .Y(n1578) );
  INVX1 U1173 ( .A(n1578), .Y(n1579) );
  AND2X2 U1174 ( .A(\mem<2><13> ), .B(n104), .Y(n1580) );
  INVX1 U1175 ( .A(n1580), .Y(n1581) );
  AND2X2 U1177 ( .A(\mem<2><14> ), .B(n104), .Y(n1582) );
  INVX1 U1178 ( .A(n1582), .Y(n1583) );
  AND2X2 U1179 ( .A(\mem<2><15> ), .B(n104), .Y(n1584) );
  INVX1 U1180 ( .A(n1584), .Y(n1585) );
  AND2X2 U1181 ( .A(\mem<1><0> ), .B(n108), .Y(n1586) );
  INVX1 U1182 ( .A(n1586), .Y(n1587) );
  AND2X2 U1183 ( .A(\mem<1><1> ), .B(n108), .Y(n1588) );
  INVX1 U1184 ( .A(n1588), .Y(n1589) );
  AND2X2 U1185 ( .A(\mem<1><2> ), .B(n108), .Y(n1590) );
  INVX1 U1186 ( .A(n1590), .Y(n1591) );
  AND2X2 U1187 ( .A(\mem<1><3> ), .B(n108), .Y(n1592) );
  INVX1 U1188 ( .A(n1592), .Y(n1593) );
  AND2X2 U1189 ( .A(\mem<1><4> ), .B(n108), .Y(n1594) );
  INVX1 U1190 ( .A(n1594), .Y(n1595) );
  AND2X2 U1191 ( .A(\mem<1><5> ), .B(n108), .Y(n1596) );
  INVX1 U1192 ( .A(n1596), .Y(n1597) );
  AND2X2 U1193 ( .A(\mem<1><6> ), .B(n108), .Y(n1598) );
  INVX1 U1194 ( .A(n1598), .Y(n1599) );
  AND2X2 U1195 ( .A(\mem<1><7> ), .B(n108), .Y(n1600) );
  INVX1 U1196 ( .A(n1600), .Y(n1601) );
  AND2X2 U1197 ( .A(\mem<1><8> ), .B(n107), .Y(n1602) );
  INVX1 U1198 ( .A(n1602), .Y(n1603) );
  AND2X2 U1199 ( .A(\mem<1><9> ), .B(n107), .Y(n1604) );
  INVX1 U1200 ( .A(n1604), .Y(n1605) );
  AND2X2 U1201 ( .A(\mem<1><10> ), .B(n107), .Y(n1606) );
  INVX1 U1202 ( .A(n1606), .Y(n1607) );
  AND2X2 U1203 ( .A(\mem<1><11> ), .B(n107), .Y(n1608) );
  INVX1 U1204 ( .A(n1608), .Y(n1609) );
  AND2X2 U1205 ( .A(\mem<1><12> ), .B(n107), .Y(n1610) );
  INVX1 U1206 ( .A(n1610), .Y(n1611) );
  AND2X2 U1207 ( .A(\mem<1><13> ), .B(n107), .Y(n1612) );
  INVX1 U1208 ( .A(n1612), .Y(n1613) );
  AND2X2 U1209 ( .A(\mem<1><14> ), .B(n107), .Y(n1614) );
  INVX1 U1210 ( .A(n1614), .Y(n1615) );
  AND2X2 U1211 ( .A(\mem<1><15> ), .B(n107), .Y(n1616) );
  INVX1 U1212 ( .A(n1616), .Y(n1617) );
  AND2X2 U1213 ( .A(\mem<0><0> ), .B(n27), .Y(n1618) );
  INVX1 U1214 ( .A(n1618), .Y(n1619) );
  AND2X2 U1215 ( .A(\mem<0><1> ), .B(n27), .Y(n1620) );
  INVX1 U1216 ( .A(n1620), .Y(n1621) );
  AND2X2 U1217 ( .A(\mem<0><2> ), .B(n27), .Y(n1622) );
  INVX1 U1218 ( .A(n1622), .Y(n1623) );
  AND2X2 U1219 ( .A(\mem<0><3> ), .B(n27), .Y(n1624) );
  INVX1 U1220 ( .A(n1624), .Y(n1625) );
  AND2X2 U1221 ( .A(\mem<0><4> ), .B(n27), .Y(n1626) );
  INVX1 U1222 ( .A(n1626), .Y(n1627) );
  AND2X2 U1223 ( .A(\mem<0><5> ), .B(n27), .Y(n1628) );
  INVX1 U1224 ( .A(n1628), .Y(n1629) );
  AND2X2 U1225 ( .A(\mem<0><6> ), .B(n27), .Y(n1630) );
  INVX1 U1226 ( .A(n1630), .Y(n1631) );
  AND2X2 U1227 ( .A(\mem<0><7> ), .B(n27), .Y(n1632) );
  INVX1 U1228 ( .A(n1632), .Y(n1633) );
  AND2X2 U1229 ( .A(\mem<0><8> ), .B(n27), .Y(n1634) );
  INVX1 U1230 ( .A(n1634), .Y(n1635) );
  AND2X2 U1231 ( .A(\mem<0><9> ), .B(n27), .Y(n1636) );
  INVX1 U1232 ( .A(n1636), .Y(n1637) );
  AND2X2 U1233 ( .A(\mem<0><10> ), .B(n27), .Y(n1638) );
  INVX1 U1234 ( .A(n1638), .Y(n1639) );
  AND2X2 U1235 ( .A(\mem<0><11> ), .B(n27), .Y(n1640) );
  INVX1 U1236 ( .A(n1640), .Y(n1641) );
  AND2X2 U1237 ( .A(\mem<0><12> ), .B(n27), .Y(n1642) );
  INVX1 U1238 ( .A(n1642), .Y(n1643) );
  AND2X2 U1239 ( .A(\mem<0><13> ), .B(n27), .Y(n1644) );
  INVX1 U1240 ( .A(n1644), .Y(n1645) );
  AND2X2 U1241 ( .A(\mem<0><14> ), .B(n27), .Y(n1646) );
  INVX1 U1242 ( .A(n1646), .Y(n1647) );
  AND2X2 U1243 ( .A(\mem<0><15> ), .B(n27), .Y(n1648) );
  INVX1 U1244 ( .A(n1648), .Y(n1649) );
  BUFX2 U1245 ( .A(n2385), .Y(n1650) );
  INVX1 U1246 ( .A(n1650), .Y(n2393) );
  BUFX2 U1247 ( .A(n2386), .Y(n1651) );
  INVX1 U1248 ( .A(n1651), .Y(n2394) );
  BUFX2 U1249 ( .A(n2387), .Y(n1652) );
  INVX1 U1250 ( .A(n1652), .Y(n2395) );
  BUFX2 U1251 ( .A(n2388), .Y(n1653) );
  INVX1 U1252 ( .A(n1653), .Y(n2396) );
  BUFX2 U1253 ( .A(n2389), .Y(n1654) );
  INVX1 U1254 ( .A(n1654), .Y(n2397) );
  BUFX2 U1255 ( .A(n2390), .Y(n1655) );
  INVX1 U1256 ( .A(n1655), .Y(n2391) );
  BUFX2 U1257 ( .A(n2392), .Y(n1656) );
  INVX1 U1258 ( .A(n1656), .Y(n2398) );
  AND2X1 U1259 ( .A(n2376), .B(n181), .Y(n1657) );
  AND2X1 U1260 ( .A(n2381), .B(n182), .Y(n1658) );
  INVX4 U1261 ( .A(n30), .Y(n2341) );
  INVX1 U1262 ( .A(n30), .Y(n2342) );
  INVX4 U1263 ( .A(n37), .Y(n2344) );
  INVX4 U1264 ( .A(n38), .Y(n2346) );
  INVX4 U1265 ( .A(n39), .Y(n2348) );
  INVX4 U1266 ( .A(n40), .Y(n2350) );
  INVX4 U1267 ( .A(n41), .Y(n2352) );
  INVX4 U1268 ( .A(n42), .Y(n2354) );
  INVX4 U1269 ( .A(n43), .Y(n2356) );
  INVX4 U1270 ( .A(n44), .Y(n2358) );
  INVX4 U1271 ( .A(n45), .Y(n2360) );
  INVX4 U1272 ( .A(n46), .Y(n2362) );
  INVX4 U1273 ( .A(n47), .Y(n2364) );
  INVX4 U1274 ( .A(n48), .Y(n2366) );
  INVX4 U1275 ( .A(n49), .Y(n2368) );
  INVX4 U1276 ( .A(n50), .Y(n2370) );
  INVX4 U1277 ( .A(n51), .Y(n2372) );
  INVX4 U1278 ( .A(n52), .Y(n2374) );
  AND2X1 U1279 ( .A(n2377), .B(n181), .Y(n1659) );
  AND2X1 U1280 ( .A(n2382), .B(n182), .Y(n1660) );
  AND2X1 U1281 ( .A(n1658), .B(n2399), .Y(n1661) );
  INVX1 U1282 ( .A(n1661), .Y(n1662) );
  AND2X1 U1283 ( .A(n2399), .B(n1660), .Y(n1663) );
  AND2X1 U1284 ( .A(n2399), .B(n2391), .Y(n1664) );
  AND2X1 U1285 ( .A(n2399), .B(n2398), .Y(n1665) );
  AND2X1 U1286 ( .A(n1657), .B(n1658), .Y(n1666) );
  INVX1 U1287 ( .A(n1666), .Y(n1667) );
  AND2X1 U1288 ( .A(n1658), .B(n1659), .Y(n1668) );
  INVX1 U1289 ( .A(n1668), .Y(n1669) );
  AND2X1 U1290 ( .A(n1658), .B(n2393), .Y(n1670) );
  INVX1 U1291 ( .A(n1670), .Y(n1671) );
  AND2X1 U1292 ( .A(n1658), .B(n2394), .Y(n1672) );
  INVX1 U1293 ( .A(n1672), .Y(n1673) );
  AND2X1 U1294 ( .A(n1658), .B(n2395), .Y(n1674) );
  INVX1 U1295 ( .A(n1674), .Y(n1675) );
  AND2X1 U1296 ( .A(n1658), .B(n2396), .Y(n1676) );
  INVX1 U1297 ( .A(n1676), .Y(n1677) );
  BUFX2 U1298 ( .A(n7), .Y(n2287) );
  AND2X1 U1299 ( .A(n1658), .B(n2397), .Y(n1678) );
  INVX1 U1300 ( .A(n1678), .Y(n1679) );
  AND2X1 U1301 ( .A(n1657), .B(n1660), .Y(n1680) );
  INVX1 U1302 ( .A(n1680), .Y(n1681) );
  AND2X1 U1303 ( .A(n1659), .B(n1660), .Y(n1682) );
  INVX1 U1304 ( .A(n1682), .Y(n1683) );
  BUFX2 U1305 ( .A(n15), .Y(n2294) );
  AND2X1 U1306 ( .A(n2393), .B(n1660), .Y(n1684) );
  INVX1 U1307 ( .A(n1684), .Y(n1685) );
  AND2X1 U1308 ( .A(n2394), .B(n1660), .Y(n1686) );
  INVX1 U1309 ( .A(n1686), .Y(n1687) );
  BUFX2 U1310 ( .A(n21), .Y(n2299) );
  AND2X1 U1311 ( .A(n2395), .B(n1660), .Y(n1688) );
  INVX1 U1312 ( .A(n1688), .Y(n1689) );
  BUFX2 U1313 ( .A(n23), .Y(n2302) );
  AND2X1 U1314 ( .A(n2396), .B(n1660), .Y(n1690) );
  INVX1 U1315 ( .A(n1690), .Y(n1691) );
  AND2X1 U1316 ( .A(n2397), .B(n1660), .Y(n1692) );
  INVX1 U1317 ( .A(n1692), .Y(n1693) );
  AND2X1 U1318 ( .A(n1657), .B(n2391), .Y(n1694) );
  INVX1 U1319 ( .A(n1694), .Y(n1695) );
  AND2X1 U1320 ( .A(n1659), .B(n2391), .Y(n1696) );
  INVX1 U1321 ( .A(n1696), .Y(n1697) );
  AND2X1 U1322 ( .A(n2393), .B(n2391), .Y(n1698) );
  INVX1 U1323 ( .A(n1698), .Y(n1699) );
  AND2X1 U1324 ( .A(n2394), .B(n2391), .Y(n1700) );
  INVX1 U1325 ( .A(n1700), .Y(n1701) );
  AND2X1 U1326 ( .A(n2395), .B(n2391), .Y(n1702) );
  INVX1 U1327 ( .A(n1702), .Y(n1703) );
  AND2X1 U1328 ( .A(n2396), .B(n2391), .Y(n1704) );
  INVX1 U1329 ( .A(n1704), .Y(n1705) );
  AND2X1 U1330 ( .A(n2397), .B(n2391), .Y(n1706) );
  INVX1 U1331 ( .A(n1706), .Y(n1707) );
  AND2X1 U1332 ( .A(n1657), .B(n2398), .Y(n1708) );
  INVX1 U1333 ( .A(n1708), .Y(n1709) );
  AND2X1 U1334 ( .A(n1659), .B(n2398), .Y(n1710) );
  INVX1 U1335 ( .A(n1710), .Y(n1711) );
  AND2X1 U1336 ( .A(n2393), .B(n2398), .Y(n1712) );
  INVX1 U1337 ( .A(n1712), .Y(n1713) );
  AND2X1 U1338 ( .A(n2394), .B(n2398), .Y(n1714) );
  INVX1 U1339 ( .A(n1714), .Y(n1715) );
  AND2X1 U1340 ( .A(n2395), .B(n2398), .Y(n1716) );
  INVX1 U1341 ( .A(n1716), .Y(n1717) );
  AND2X1 U1342 ( .A(n2396), .B(n2398), .Y(n1718) );
  INVX1 U1343 ( .A(n1718), .Y(n1719) );
  AND2X1 U1344 ( .A(n2397), .B(n2398), .Y(n1720) );
  INVX1 U1345 ( .A(n1720), .Y(n1721) );
  INVX1 U1346 ( .A(write), .Y(n1722) );
  INVX1 U1347 ( .A(n1722), .Y(n1723) );
  INVX1 U1348 ( .A(N12), .Y(n2380) );
  MUX2X1 U1349 ( .B(n1725), .A(n1726), .S(n2232), .Y(n1724) );
  MUX2X1 U1350 ( .B(n1728), .A(n1729), .S(n2232), .Y(n1727) );
  MUX2X1 U1351 ( .B(n1731), .A(n1732), .S(n2232), .Y(n1730) );
  MUX2X1 U1352 ( .B(n1734), .A(n1735), .S(n2232), .Y(n1733) );
  MUX2X1 U1353 ( .B(n1737), .A(n1738), .S(n2223), .Y(n1736) );
  MUX2X1 U1354 ( .B(n1740), .A(n1741), .S(n2232), .Y(n1739) );
  MUX2X1 U1355 ( .B(n1743), .A(n1744), .S(n2232), .Y(n1742) );
  MUX2X1 U1356 ( .B(n1746), .A(n1747), .S(n2232), .Y(n1745) );
  MUX2X1 U1357 ( .B(n1749), .A(n1750), .S(n2232), .Y(n1748) );
  MUX2X1 U1358 ( .B(n1752), .A(n1753), .S(n2223), .Y(n1751) );
  MUX2X1 U1359 ( .B(n1755), .A(n1756), .S(n2233), .Y(n1754) );
  MUX2X1 U1360 ( .B(n1758), .A(n1759), .S(n2233), .Y(n1757) );
  MUX2X1 U1361 ( .B(n1761), .A(n1762), .S(n2233), .Y(n1760) );
  MUX2X1 U1362 ( .B(n1764), .A(n1765), .S(n2233), .Y(n1763) );
  MUX2X1 U1363 ( .B(n1767), .A(n1768), .S(n2223), .Y(n1766) );
  MUX2X1 U1364 ( .B(n1770), .A(n1771), .S(n2233), .Y(n1769) );
  MUX2X1 U1365 ( .B(n1773), .A(n1774), .S(n2233), .Y(n1772) );
  MUX2X1 U1366 ( .B(n1776), .A(n1777), .S(n2233), .Y(n1775) );
  MUX2X1 U1367 ( .B(n1779), .A(n1780), .S(n2233), .Y(n1778) );
  MUX2X1 U1368 ( .B(n1782), .A(n1783), .S(n2223), .Y(n1781) );
  MUX2X1 U1369 ( .B(n1785), .A(n1786), .S(n2233), .Y(n1784) );
  MUX2X1 U1370 ( .B(n1788), .A(n1789), .S(n2233), .Y(n1787) );
  MUX2X1 U1371 ( .B(n1791), .A(n1792), .S(n2233), .Y(n1790) );
  MUX2X1 U1372 ( .B(n1794), .A(n1795), .S(n2233), .Y(n1793) );
  MUX2X1 U1373 ( .B(n1797), .A(n1798), .S(n2223), .Y(n1796) );
  MUX2X1 U1374 ( .B(n1800), .A(n1801), .S(n2233), .Y(n1799) );
  MUX2X1 U1375 ( .B(n1803), .A(n1804), .S(n2233), .Y(n1802) );
  MUX2X1 U1376 ( .B(n1806), .A(n1807), .S(n2233), .Y(n1805) );
  MUX2X1 U1377 ( .B(n1809), .A(n1810), .S(n2233), .Y(n1808) );
  MUX2X1 U1378 ( .B(n1812), .A(n1813), .S(n2223), .Y(n1811) );
  MUX2X1 U1379 ( .B(n1815), .A(n1816), .S(n2233), .Y(n1814) );
  MUX2X1 U1380 ( .B(n1818), .A(n1819), .S(n2233), .Y(n1817) );
  MUX2X1 U1381 ( .B(n1821), .A(n1822), .S(n2233), .Y(n1820) );
  MUX2X1 U1382 ( .B(n1824), .A(n1825), .S(n2233), .Y(n1823) );
  MUX2X1 U1383 ( .B(n1827), .A(n1828), .S(n2223), .Y(n1826) );
  MUX2X1 U1384 ( .B(n1830), .A(n1831), .S(n2233), .Y(n1829) );
  MUX2X1 U1385 ( .B(n1833), .A(n1834), .S(n2233), .Y(n1832) );
  MUX2X1 U1386 ( .B(n1836), .A(n1837), .S(n2233), .Y(n1835) );
  MUX2X1 U1387 ( .B(n1839), .A(n1840), .S(n2233), .Y(n1838) );
  MUX2X1 U1388 ( .B(n1842), .A(n1843), .S(n2223), .Y(n1841) );
  MUX2X1 U1389 ( .B(n1845), .A(n1846), .S(n2234), .Y(n1844) );
  MUX2X1 U1390 ( .B(n1848), .A(n1849), .S(n2234), .Y(n1847) );
  MUX2X1 U1391 ( .B(n1851), .A(n1852), .S(n2234), .Y(n1850) );
  MUX2X1 U1392 ( .B(n1854), .A(n1855), .S(n2234), .Y(n1853) );
  MUX2X1 U1393 ( .B(n1857), .A(n1858), .S(n2223), .Y(n1856) );
  MUX2X1 U1394 ( .B(n1860), .A(n1861), .S(n2234), .Y(n1859) );
  MUX2X1 U1395 ( .B(n1863), .A(n1864), .S(n2234), .Y(n1862) );
  MUX2X1 U1396 ( .B(n1866), .A(n1867), .S(n2234), .Y(n1865) );
  MUX2X1 U1397 ( .B(n1869), .A(n1870), .S(n2234), .Y(n1868) );
  MUX2X1 U1398 ( .B(n1872), .A(n1873), .S(n2223), .Y(n1871) );
  MUX2X1 U1399 ( .B(n1875), .A(n1876), .S(n2234), .Y(n1874) );
  MUX2X1 U1400 ( .B(n1878), .A(n1879), .S(n2234), .Y(n1877) );
  MUX2X1 U1401 ( .B(n1881), .A(n1882), .S(n2234), .Y(n1880) );
  MUX2X1 U1402 ( .B(n1884), .A(n1885), .S(n2234), .Y(n1883) );
  MUX2X1 U1403 ( .B(n1887), .A(n1888), .S(n2223), .Y(n1886) );
  MUX2X1 U1404 ( .B(n1890), .A(n1891), .S(n2235), .Y(n1889) );
  MUX2X1 U1405 ( .B(n1893), .A(n1894), .S(n2235), .Y(n1892) );
  MUX2X1 U1406 ( .B(n1896), .A(n1897), .S(n2235), .Y(n1895) );
  MUX2X1 U1407 ( .B(n1899), .A(n1900), .S(n2235), .Y(n1898) );
  MUX2X1 U1408 ( .B(n1902), .A(n1903), .S(n2223), .Y(n1901) );
  MUX2X1 U1409 ( .B(n1905), .A(n1906), .S(n2235), .Y(n1904) );
  MUX2X1 U1410 ( .B(n1908), .A(n1909), .S(n2235), .Y(n1907) );
  MUX2X1 U1411 ( .B(n1911), .A(n1912), .S(n2235), .Y(n1910) );
  MUX2X1 U1412 ( .B(n1914), .A(n1915), .S(n2235), .Y(n1913) );
  MUX2X1 U1413 ( .B(n1917), .A(n1918), .S(n2222), .Y(n1916) );
  MUX2X1 U1414 ( .B(n1920), .A(n1921), .S(n2235), .Y(n1919) );
  MUX2X1 U1415 ( .B(n1923), .A(n1924), .S(n2235), .Y(n1922) );
  MUX2X1 U1416 ( .B(n1926), .A(n1927), .S(n2235), .Y(n1925) );
  MUX2X1 U1417 ( .B(n1929), .A(n1930), .S(n2235), .Y(n1928) );
  MUX2X1 U1418 ( .B(n1932), .A(n1933), .S(n2222), .Y(n1931) );
  MUX2X1 U1419 ( .B(n1935), .A(n1936), .S(n2236), .Y(n1934) );
  MUX2X1 U1420 ( .B(n1938), .A(n1939), .S(n2236), .Y(n1937) );
  MUX2X1 U1421 ( .B(n1941), .A(n1942), .S(n2236), .Y(n1940) );
  MUX2X1 U1422 ( .B(n1944), .A(n1945), .S(n2236), .Y(n1943) );
  MUX2X1 U1423 ( .B(n1947), .A(n1948), .S(n2222), .Y(n1946) );
  MUX2X1 U1424 ( .B(n1950), .A(n1951), .S(n2236), .Y(n1949) );
  MUX2X1 U1425 ( .B(n1953), .A(n1954), .S(n2236), .Y(n1952) );
  MUX2X1 U1426 ( .B(n1956), .A(n1957), .S(n2236), .Y(n1955) );
  MUX2X1 U1427 ( .B(n1959), .A(n1960), .S(n2236), .Y(n1958) );
  MUX2X1 U1428 ( .B(n1962), .A(n1963), .S(n2222), .Y(n1961) );
  MUX2X1 U1429 ( .B(n1965), .A(n1966), .S(n2236), .Y(n1964) );
  MUX2X1 U1430 ( .B(n1968), .A(n1969), .S(n2236), .Y(n1967) );
  MUX2X1 U1431 ( .B(n1971), .A(n1972), .S(n2236), .Y(n1970) );
  MUX2X1 U1432 ( .B(n1974), .A(n1975), .S(n2236), .Y(n1973) );
  MUX2X1 U1433 ( .B(n1977), .A(n1978), .S(n2222), .Y(n1976) );
  MUX2X1 U1434 ( .B(n1980), .A(n1981), .S(n2237), .Y(n1979) );
  MUX2X1 U1435 ( .B(n1983), .A(n1984), .S(n2237), .Y(n1982) );
  MUX2X1 U1436 ( .B(n1986), .A(n1987), .S(n2237), .Y(n1985) );
  MUX2X1 U1437 ( .B(n1989), .A(n1990), .S(n2237), .Y(n1988) );
  MUX2X1 U1438 ( .B(n1992), .A(n1993), .S(n2222), .Y(n1991) );
  MUX2X1 U1439 ( .B(n1995), .A(n1996), .S(n2237), .Y(n1994) );
  MUX2X1 U1440 ( .B(n1998), .A(n1999), .S(n2237), .Y(n1997) );
  MUX2X1 U1441 ( .B(n2001), .A(n2002), .S(n2237), .Y(n2000) );
  MUX2X1 U1442 ( .B(n2004), .A(n2005), .S(n2237), .Y(n2003) );
  MUX2X1 U1443 ( .B(n2007), .A(n2008), .S(n2222), .Y(n2006) );
  MUX2X1 U1444 ( .B(n2010), .A(n2011), .S(n2237), .Y(n2009) );
  MUX2X1 U1445 ( .B(n2013), .A(n2014), .S(n2237), .Y(n2012) );
  MUX2X1 U1446 ( .B(n2016), .A(n2017), .S(n2237), .Y(n2015) );
  MUX2X1 U1447 ( .B(n2019), .A(n2020), .S(n2237), .Y(n2018) );
  MUX2X1 U1448 ( .B(n2022), .A(n2023), .S(n2222), .Y(n2021) );
  MUX2X1 U1449 ( .B(n2025), .A(n2026), .S(n2238), .Y(n2024) );
  MUX2X1 U1450 ( .B(n2028), .A(n2029), .S(n2238), .Y(n2027) );
  MUX2X1 U1451 ( .B(n2031), .A(n2032), .S(n2238), .Y(n2030) );
  MUX2X1 U1452 ( .B(n2034), .A(n2035), .S(n2238), .Y(n2033) );
  MUX2X1 U1453 ( .B(n2037), .A(n2038), .S(n2222), .Y(n2036) );
  MUX2X1 U1454 ( .B(n2040), .A(n2041), .S(n2238), .Y(n2039) );
  MUX2X1 U1455 ( .B(n2043), .A(n2044), .S(n2238), .Y(n2042) );
  MUX2X1 U1456 ( .B(n2046), .A(n2047), .S(n2238), .Y(n2045) );
  MUX2X1 U1457 ( .B(n2049), .A(n2050), .S(n2238), .Y(n2048) );
  MUX2X1 U1458 ( .B(n2052), .A(n2053), .S(n2222), .Y(n2051) );
  MUX2X1 U1459 ( .B(n2055), .A(n2056), .S(n2238), .Y(n2054) );
  MUX2X1 U1460 ( .B(n2058), .A(n2059), .S(n2238), .Y(n2057) );
  MUX2X1 U1461 ( .B(n2061), .A(n2062), .S(n2238), .Y(n2060) );
  MUX2X1 U1462 ( .B(n2064), .A(n2065), .S(n2238), .Y(n2063) );
  MUX2X1 U1463 ( .B(n2067), .A(n2068), .S(n2222), .Y(n2066) );
  MUX2X1 U1464 ( .B(n2070), .A(n2071), .S(n2239), .Y(n2069) );
  MUX2X1 U1465 ( .B(n2073), .A(n2074), .S(n2239), .Y(n2072) );
  MUX2X1 U1466 ( .B(n2076), .A(n2077), .S(n2239), .Y(n2075) );
  MUX2X1 U1467 ( .B(n2079), .A(n2080), .S(n2239), .Y(n2078) );
  MUX2X1 U1468 ( .B(n2082), .A(n2083), .S(n2222), .Y(n2081) );
  MUX2X1 U1469 ( .B(n2085), .A(n2086), .S(n2239), .Y(n2084) );
  MUX2X1 U1470 ( .B(n2088), .A(n2089), .S(n2239), .Y(n2087) );
  MUX2X1 U1471 ( .B(n2091), .A(n2092), .S(n2239), .Y(n2090) );
  MUX2X1 U1472 ( .B(n2094), .A(n2095), .S(n2239), .Y(n2093) );
  MUX2X1 U1473 ( .B(n2097), .A(n2098), .S(n2381), .Y(n2096) );
  MUX2X1 U1474 ( .B(n2100), .A(n2101), .S(n2239), .Y(n2099) );
  MUX2X1 U1475 ( .B(n2103), .A(n2104), .S(n2239), .Y(n2102) );
  MUX2X1 U1476 ( .B(n2106), .A(n2107), .S(n2239), .Y(n2105) );
  MUX2X1 U1477 ( .B(n2109), .A(n2110), .S(n2239), .Y(n2108) );
  MUX2X1 U1478 ( .B(n2112), .A(n2113), .S(n2381), .Y(n2111) );
  MUX2X1 U1479 ( .B(n2115), .A(n2116), .S(n2240), .Y(n2114) );
  MUX2X1 U1480 ( .B(n2118), .A(n2119), .S(n2240), .Y(n2117) );
  MUX2X1 U1481 ( .B(n2121), .A(n2122), .S(n2240), .Y(n2120) );
  MUX2X1 U1482 ( .B(n2124), .A(n2125), .S(n2240), .Y(n2123) );
  MUX2X1 U1483 ( .B(n2127), .A(n2128), .S(n2222), .Y(n2126) );
  MUX2X1 U1484 ( .B(n2130), .A(n2131), .S(n2240), .Y(n2129) );
  MUX2X1 U1485 ( .B(n2133), .A(n2134), .S(n2240), .Y(n2132) );
  MUX2X1 U1486 ( .B(n2136), .A(n2137), .S(n2240), .Y(n2135) );
  MUX2X1 U1487 ( .B(n2139), .A(n2140), .S(n2240), .Y(n2138) );
  MUX2X1 U1488 ( .B(n2142), .A(n2143), .S(n2222), .Y(n2141) );
  MUX2X1 U1489 ( .B(n2145), .A(n2146), .S(n2240), .Y(n2144) );
  MUX2X1 U1490 ( .B(n2148), .A(n2149), .S(n2240), .Y(n2147) );
  MUX2X1 U1491 ( .B(n2151), .A(n2152), .S(n2240), .Y(n2150) );
  MUX2X1 U1492 ( .B(n2154), .A(n2155), .S(n2240), .Y(n2153) );
  MUX2X1 U1493 ( .B(n2157), .A(n2158), .S(n2222), .Y(n2156) );
  MUX2X1 U1494 ( .B(n2160), .A(n2161), .S(n2241), .Y(n2159) );
  MUX2X1 U1495 ( .B(n2163), .A(n2164), .S(n2241), .Y(n2162) );
  MUX2X1 U1496 ( .B(n2166), .A(n2167), .S(n2241), .Y(n2165) );
  MUX2X1 U1497 ( .B(n2169), .A(n2170), .S(n2241), .Y(n2168) );
  MUX2X1 U1498 ( .B(n2172), .A(n2173), .S(n2222), .Y(n2171) );
  MUX2X1 U1499 ( .B(n2175), .A(n2176), .S(n2241), .Y(n2174) );
  MUX2X1 U1500 ( .B(n2178), .A(n2179), .S(n2241), .Y(n2177) );
  MUX2X1 U1501 ( .B(n2181), .A(n2182), .S(n2241), .Y(n2180) );
  MUX2X1 U1502 ( .B(n2184), .A(n2185), .S(n2241), .Y(n2183) );
  MUX2X1 U1503 ( .B(n2187), .A(n2188), .S(n2222), .Y(n2186) );
  MUX2X1 U1504 ( .B(n2190), .A(n2191), .S(n2241), .Y(n2189) );
  MUX2X1 U1505 ( .B(n2193), .A(n2194), .S(n2241), .Y(n2192) );
  MUX2X1 U1506 ( .B(n2196), .A(n2197), .S(n2241), .Y(n2195) );
  MUX2X1 U1507 ( .B(n2199), .A(n2200), .S(n2241), .Y(n2198) );
  MUX2X1 U1508 ( .B(n2202), .A(n2203), .S(n2222), .Y(n2201) );
  MUX2X1 U1509 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n2250), .Y(n1726) );
  MUX2X1 U1510 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n2250), .Y(n1725) );
  MUX2X1 U1511 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n2250), .Y(n1729) );
  MUX2X1 U1512 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n2250), .Y(n1728) );
  MUX2X1 U1513 ( .B(n1727), .A(n1724), .S(n2230), .Y(n1738) );
  MUX2X1 U1514 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n2251), .Y(n1732) );
  MUX2X1 U1515 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n2251), .Y(n1731) );
  MUX2X1 U1516 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n2251), .Y(n1735) );
  MUX2X1 U1517 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n2251), .Y(n1734) );
  MUX2X1 U1518 ( .B(n1733), .A(n1730), .S(n2230), .Y(n1737) );
  MUX2X1 U1519 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n2251), .Y(n1741) );
  MUX2X1 U1520 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n2251), .Y(n1740) );
  MUX2X1 U1521 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n2251), .Y(n1744) );
  MUX2X1 U1522 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n2251), .Y(n1743) );
  MUX2X1 U1523 ( .B(n1742), .A(n1739), .S(n2230), .Y(n1753) );
  MUX2X1 U1524 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n2251), .Y(n1747) );
  MUX2X1 U1525 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n2251), .Y(n1746) );
  MUX2X1 U1526 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n2251), .Y(n1750) );
  MUX2X1 U1527 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n2251), .Y(n1749) );
  MUX2X1 U1528 ( .B(n1748), .A(n1745), .S(n2230), .Y(n1752) );
  MUX2X1 U1529 ( .B(n1751), .A(n1736), .S(n2221), .Y(n2204) );
  MUX2X1 U1530 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n2252), .Y(n1756) );
  MUX2X1 U1531 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n2252), .Y(n1755) );
  MUX2X1 U1532 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n2252), .Y(n1759) );
  MUX2X1 U1533 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n2252), .Y(n1758) );
  MUX2X1 U1534 ( .B(n1757), .A(n1754), .S(n2230), .Y(n1768) );
  MUX2X1 U1535 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n2252), .Y(n1762) );
  MUX2X1 U1536 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n2252), .Y(n1761) );
  MUX2X1 U1537 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n2252), .Y(n1765) );
  MUX2X1 U1538 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n2252), .Y(n1764) );
  MUX2X1 U1539 ( .B(n1763), .A(n1760), .S(n2230), .Y(n1767) );
  MUX2X1 U1540 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n2252), .Y(n1771) );
  MUX2X1 U1541 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n2252), .Y(n1770) );
  MUX2X1 U1542 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n2252), .Y(n1774) );
  MUX2X1 U1543 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n2252), .Y(n1773) );
  MUX2X1 U1544 ( .B(n1772), .A(n1769), .S(n2230), .Y(n1783) );
  MUX2X1 U1545 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n2253), .Y(n1777) );
  MUX2X1 U1546 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n2253), .Y(n1776) );
  MUX2X1 U1547 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n2253), .Y(n1780) );
  MUX2X1 U1548 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n2253), .Y(n1779) );
  MUX2X1 U1549 ( .B(n1778), .A(n1775), .S(n2230), .Y(n1782) );
  MUX2X1 U1550 ( .B(n1781), .A(n1766), .S(n2221), .Y(n2205) );
  MUX2X1 U1551 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n2253), .Y(n1786) );
  MUX2X1 U1552 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n2253), .Y(n1785) );
  MUX2X1 U1553 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n2253), .Y(n1789) );
  MUX2X1 U1554 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n2253), .Y(n1788) );
  MUX2X1 U1555 ( .B(n1787), .A(n1784), .S(n2230), .Y(n1798) );
  MUX2X1 U1556 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n2253), .Y(n1792) );
  MUX2X1 U1557 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n2253), .Y(n1791) );
  MUX2X1 U1558 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n2253), .Y(n1795) );
  MUX2X1 U1559 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n2253), .Y(n1794) );
  MUX2X1 U1560 ( .B(n1793), .A(n1790), .S(n2230), .Y(n1797) );
  MUX2X1 U1561 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n2254), .Y(n1801) );
  MUX2X1 U1562 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n2254), .Y(n1800) );
  MUX2X1 U1563 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n2254), .Y(n1804) );
  MUX2X1 U1564 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n2254), .Y(n1803) );
  MUX2X1 U1565 ( .B(n1802), .A(n1799), .S(n2230), .Y(n1813) );
  MUX2X1 U1566 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n2254), .Y(n1807) );
  MUX2X1 U1567 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n2254), .Y(n1806) );
  MUX2X1 U1568 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n2254), .Y(n1810) );
  MUX2X1 U1569 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n2254), .Y(n1809) );
  MUX2X1 U1570 ( .B(n1808), .A(n1805), .S(n2230), .Y(n1812) );
  MUX2X1 U1571 ( .B(n1811), .A(n1796), .S(n2221), .Y(n2206) );
  MUX2X1 U1572 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n2254), .Y(n1816) );
  MUX2X1 U1573 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n2254), .Y(n1815) );
  MUX2X1 U1574 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n2254), .Y(n1819) );
  MUX2X1 U1575 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n2254), .Y(n1818) );
  MUX2X1 U1576 ( .B(n1817), .A(n1814), .S(n2229), .Y(n1828) );
  MUX2X1 U1577 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n2255), .Y(n1822) );
  MUX2X1 U1578 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n2255), .Y(n1821) );
  MUX2X1 U1579 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n2255), .Y(n1825) );
  MUX2X1 U1580 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n2255), .Y(n1824) );
  MUX2X1 U1581 ( .B(n1823), .A(n1820), .S(n2229), .Y(n1827) );
  MUX2X1 U1582 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n2255), .Y(n1831) );
  MUX2X1 U1583 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n2255), .Y(n1830) );
  MUX2X1 U1584 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n2255), .Y(n1834) );
  MUX2X1 U1585 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n2255), .Y(n1833) );
  MUX2X1 U1586 ( .B(n1832), .A(n1829), .S(n2229), .Y(n1843) );
  MUX2X1 U1587 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n2255), .Y(n1837) );
  MUX2X1 U1588 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n2255), .Y(n1836) );
  MUX2X1 U1589 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n2255), .Y(n1840) );
  MUX2X1 U1590 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n2255), .Y(n1839) );
  MUX2X1 U1591 ( .B(n1838), .A(n1835), .S(n2229), .Y(n1842) );
  MUX2X1 U1592 ( .B(n1841), .A(n1826), .S(n2221), .Y(n2207) );
  MUX2X1 U1593 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n2256), .Y(n1846) );
  MUX2X1 U1594 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n2256), .Y(n1845) );
  MUX2X1 U1595 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n2256), .Y(n1849) );
  MUX2X1 U1596 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n2256), .Y(n1848) );
  MUX2X1 U1597 ( .B(n1847), .A(n1844), .S(n2229), .Y(n1858) );
  MUX2X1 U1598 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n2256), .Y(n1852) );
  MUX2X1 U1599 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n2256), .Y(n1851) );
  MUX2X1 U1600 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n2256), .Y(n1855) );
  MUX2X1 U1601 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n2256), .Y(n1854) );
  MUX2X1 U1602 ( .B(n1853), .A(n1850), .S(n2229), .Y(n1857) );
  MUX2X1 U1603 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n2256), .Y(n1861) );
  MUX2X1 U1604 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n2256), .Y(n1860) );
  MUX2X1 U1605 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n2256), .Y(n1864) );
  MUX2X1 U1606 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n2256), .Y(n1863) );
  MUX2X1 U1607 ( .B(n1862), .A(n1859), .S(n2229), .Y(n1873) );
  MUX2X1 U1608 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n2257), .Y(n1867) );
  MUX2X1 U1609 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n2257), .Y(n1866) );
  MUX2X1 U1610 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n2257), .Y(n1870) );
  MUX2X1 U1611 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n2257), .Y(n1869) );
  MUX2X1 U1612 ( .B(n1868), .A(n1865), .S(n2229), .Y(n1872) );
  MUX2X1 U1613 ( .B(n1871), .A(n1856), .S(n2221), .Y(n2208) );
  MUX2X1 U1614 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n2257), .Y(n1876) );
  MUX2X1 U1615 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n2257), .Y(n1875) );
  MUX2X1 U1616 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n2257), .Y(n1879) );
  MUX2X1 U1617 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n2257), .Y(n1878) );
  MUX2X1 U1618 ( .B(n1877), .A(n1874), .S(n2229), .Y(n1888) );
  MUX2X1 U1619 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n2257), .Y(n1882) );
  MUX2X1 U1620 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n2257), .Y(n1881) );
  MUX2X1 U1621 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n2257), .Y(n1885) );
  MUX2X1 U1622 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n2257), .Y(n1884) );
  MUX2X1 U1623 ( .B(n1883), .A(n1880), .S(n2229), .Y(n1887) );
  MUX2X1 U1624 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n2258), .Y(n1891) );
  MUX2X1 U1625 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n2258), .Y(n1890) );
  MUX2X1 U1626 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n2258), .Y(n1894) );
  MUX2X1 U1627 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n2258), .Y(n1893) );
  MUX2X1 U1628 ( .B(n1892), .A(n1889), .S(n2229), .Y(n1903) );
  MUX2X1 U1629 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n2258), .Y(n1897) );
  MUX2X1 U1630 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n2258), .Y(n1896) );
  MUX2X1 U1631 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n2258), .Y(n1900) );
  MUX2X1 U1632 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n2258), .Y(n1899) );
  MUX2X1 U1633 ( .B(n1898), .A(n1895), .S(n2229), .Y(n1902) );
  MUX2X1 U1634 ( .B(n1901), .A(n1886), .S(n2221), .Y(n2209) );
  MUX2X1 U1635 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n2258), .Y(n1906) );
  MUX2X1 U1636 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n2258), .Y(n1905) );
  MUX2X1 U1637 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n2258), .Y(n1909) );
  MUX2X1 U1638 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n2258), .Y(n1908) );
  MUX2X1 U1639 ( .B(n1907), .A(n1904), .S(n2228), .Y(n1918) );
  MUX2X1 U1640 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n2259), .Y(n1912) );
  MUX2X1 U1641 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n2259), .Y(n1911) );
  MUX2X1 U1642 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n2259), .Y(n1915) );
  MUX2X1 U1643 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n2259), .Y(n1914) );
  MUX2X1 U1644 ( .B(n1913), .A(n1910), .S(n2228), .Y(n1917) );
  MUX2X1 U1645 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n2259), .Y(n1921) );
  MUX2X1 U1646 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n2259), .Y(n1920) );
  MUX2X1 U1647 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n2259), .Y(n1924) );
  MUX2X1 U1648 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n2259), .Y(n1923) );
  MUX2X1 U1649 ( .B(n1922), .A(n1919), .S(n2228), .Y(n1933) );
  MUX2X1 U1650 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n2259), .Y(n1927) );
  MUX2X1 U1651 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n2259), .Y(n1926) );
  MUX2X1 U1652 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n2259), .Y(n1930) );
  MUX2X1 U1653 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n2259), .Y(n1929) );
  MUX2X1 U1654 ( .B(n1928), .A(n1925), .S(n2228), .Y(n1932) );
  MUX2X1 U1655 ( .B(n1931), .A(n1916), .S(n2221), .Y(n2210) );
  MUX2X1 U1656 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n2260), .Y(n1936) );
  MUX2X1 U1657 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n2260), .Y(n1935) );
  MUX2X1 U1658 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n2260), .Y(n1939) );
  MUX2X1 U1659 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n2260), .Y(n1938) );
  MUX2X1 U1660 ( .B(n1937), .A(n1934), .S(n2228), .Y(n1948) );
  MUX2X1 U1661 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n2260), .Y(n1942) );
  MUX2X1 U1662 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n2260), .Y(n1941) );
  MUX2X1 U1663 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n2260), .Y(n1945) );
  MUX2X1 U1664 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n2260), .Y(n1944) );
  MUX2X1 U1665 ( .B(n1943), .A(n1940), .S(n2228), .Y(n1947) );
  MUX2X1 U1666 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n2260), .Y(n1951) );
  MUX2X1 U1667 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n2260), .Y(n1950) );
  MUX2X1 U1668 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n2260), .Y(n1954) );
  MUX2X1 U1669 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n2260), .Y(n1953) );
  MUX2X1 U1670 ( .B(n1952), .A(n1949), .S(n2228), .Y(n1963) );
  MUX2X1 U1671 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n2261), .Y(n1957) );
  MUX2X1 U1672 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n2261), .Y(n1956) );
  MUX2X1 U1673 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n2261), .Y(n1960) );
  MUX2X1 U1674 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n2261), .Y(n1959) );
  MUX2X1 U1675 ( .B(n1958), .A(n1955), .S(n2228), .Y(n1962) );
  MUX2X1 U1676 ( .B(n1961), .A(n1946), .S(n2221), .Y(n2211) );
  MUX2X1 U1677 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n2261), .Y(n1966) );
  MUX2X1 U1678 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n2261), .Y(n1965) );
  MUX2X1 U1679 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n2261), .Y(n1969) );
  MUX2X1 U1680 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n2261), .Y(n1968) );
  MUX2X1 U1681 ( .B(n1967), .A(n1964), .S(n2228), .Y(n1978) );
  MUX2X1 U1682 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n2261), .Y(n1972) );
  MUX2X1 U1683 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n2261), .Y(n1971) );
  MUX2X1 U1684 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n2261), .Y(n1975) );
  MUX2X1 U1685 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n2261), .Y(n1974) );
  MUX2X1 U1686 ( .B(n1973), .A(n1970), .S(n2228), .Y(n1977) );
  MUX2X1 U1687 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n2262), .Y(n1981) );
  MUX2X1 U1688 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n2262), .Y(n1980) );
  MUX2X1 U1689 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n2262), .Y(n1984) );
  MUX2X1 U1690 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n2262), .Y(n1983) );
  MUX2X1 U1691 ( .B(n1982), .A(n1979), .S(n2228), .Y(n1993) );
  MUX2X1 U1692 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n2262), .Y(n1987) );
  MUX2X1 U1693 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n2262), .Y(n1986) );
  MUX2X1 U1694 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n2262), .Y(n1990) );
  MUX2X1 U1695 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n2262), .Y(n1989) );
  MUX2X1 U1696 ( .B(n1988), .A(n1985), .S(n2228), .Y(n1992) );
  MUX2X1 U1697 ( .B(n1991), .A(n1976), .S(n2221), .Y(n2212) );
  MUX2X1 U1698 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n2262), .Y(n1996) );
  MUX2X1 U1699 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n2262), .Y(n1995) );
  MUX2X1 U1700 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n2262), .Y(n1999) );
  MUX2X1 U1701 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n2262), .Y(n1998) );
  MUX2X1 U1702 ( .B(n1997), .A(n1994), .S(n2227), .Y(n2008) );
  MUX2X1 U1703 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n2263), .Y(n2002) );
  MUX2X1 U1704 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n2263), .Y(n2001) );
  MUX2X1 U1705 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n2263), .Y(n2005) );
  MUX2X1 U1706 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n2263), .Y(n2004) );
  MUX2X1 U1707 ( .B(n2003), .A(n2000), .S(n2227), .Y(n2007) );
  MUX2X1 U1708 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n2263), .Y(n2011) );
  MUX2X1 U1709 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n2263), .Y(n2010) );
  MUX2X1 U1710 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n2263), .Y(n2014) );
  MUX2X1 U1711 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n2263), .Y(n2013) );
  MUX2X1 U1712 ( .B(n2012), .A(n2009), .S(n2227), .Y(n2023) );
  MUX2X1 U1713 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n2263), .Y(n2017) );
  MUX2X1 U1714 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n2263), .Y(n2016) );
  MUX2X1 U1715 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n2263), .Y(n2020) );
  MUX2X1 U1716 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n2263), .Y(n2019) );
  MUX2X1 U1717 ( .B(n2018), .A(n2015), .S(n2227), .Y(n2022) );
  MUX2X1 U1718 ( .B(n2021), .A(n2006), .S(n2221), .Y(n2213) );
  MUX2X1 U1719 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n2264), .Y(n2026) );
  MUX2X1 U1720 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n2264), .Y(n2025) );
  MUX2X1 U1721 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n2264), .Y(n2029) );
  MUX2X1 U1722 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n2264), .Y(n2028) );
  MUX2X1 U1723 ( .B(n2027), .A(n2024), .S(n2227), .Y(n2038) );
  MUX2X1 U1724 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n2264), .Y(n2032) );
  MUX2X1 U1725 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n2264), .Y(n2031) );
  MUX2X1 U1726 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n2264), .Y(n2035) );
  MUX2X1 U1727 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n2264), .Y(n2034) );
  MUX2X1 U1728 ( .B(n2033), .A(n2030), .S(n2227), .Y(n2037) );
  MUX2X1 U1729 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n2264), .Y(n2041) );
  MUX2X1 U1730 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n2264), .Y(n2040) );
  MUX2X1 U1731 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n2264), .Y(n2044) );
  MUX2X1 U1732 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n2264), .Y(n2043) );
  MUX2X1 U1733 ( .B(n2042), .A(n2039), .S(n2227), .Y(n2053) );
  MUX2X1 U1734 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n2265), .Y(n2047) );
  MUX2X1 U1735 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n2265), .Y(n2046) );
  MUX2X1 U1736 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n2265), .Y(n2050) );
  MUX2X1 U1737 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n2265), .Y(n2049) );
  MUX2X1 U1738 ( .B(n2048), .A(n2045), .S(n2227), .Y(n2052) );
  MUX2X1 U1739 ( .B(n2051), .A(n2036), .S(n2221), .Y(n2214) );
  MUX2X1 U1740 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n2265), .Y(n2056) );
  MUX2X1 U1741 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n2265), .Y(n2055) );
  MUX2X1 U1742 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n2265), .Y(n2059) );
  MUX2X1 U1743 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n2265), .Y(n2058) );
  MUX2X1 U1744 ( .B(n2057), .A(n2054), .S(n2227), .Y(n2068) );
  MUX2X1 U1745 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n2265), .Y(n2062) );
  MUX2X1 U1746 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n2265), .Y(n2061) );
  MUX2X1 U1747 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n2265), .Y(n2065) );
  MUX2X1 U1748 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n2265), .Y(n2064) );
  MUX2X1 U1749 ( .B(n2063), .A(n2060), .S(n2227), .Y(n2067) );
  MUX2X1 U1750 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n2266), .Y(n2071) );
  MUX2X1 U1751 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n2266), .Y(n2070) );
  MUX2X1 U1752 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n2266), .Y(n2074) );
  MUX2X1 U1753 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n2266), .Y(n2073) );
  MUX2X1 U1754 ( .B(n2072), .A(n2069), .S(n2227), .Y(n2083) );
  MUX2X1 U1755 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n2266), .Y(n2077) );
  MUX2X1 U1756 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n2266), .Y(n2076) );
  MUX2X1 U1757 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n2266), .Y(n2080) );
  MUX2X1 U1758 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n2266), .Y(n2079) );
  MUX2X1 U1759 ( .B(n2078), .A(n2075), .S(n2227), .Y(n2082) );
  MUX2X1 U1760 ( .B(n2081), .A(n2066), .S(n2221), .Y(n2215) );
  MUX2X1 U1761 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n2266), .Y(n2086) );
  MUX2X1 U1762 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n2266), .Y(n2085) );
  MUX2X1 U1763 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n2266), .Y(n2089) );
  MUX2X1 U1764 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n2266), .Y(n2088) );
  MUX2X1 U1765 ( .B(n2087), .A(n2084), .S(n2226), .Y(n2098) );
  MUX2X1 U1766 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n2267), .Y(n2092) );
  MUX2X1 U1767 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n2267), .Y(n2091) );
  MUX2X1 U1768 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n2267), .Y(n2095) );
  MUX2X1 U1769 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n2267), .Y(n2094) );
  MUX2X1 U1770 ( .B(n2093), .A(n2090), .S(n2226), .Y(n2097) );
  MUX2X1 U1771 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n2267), .Y(n2101) );
  MUX2X1 U1772 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n2267), .Y(n2100) );
  MUX2X1 U1773 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n2267), .Y(n2104) );
  MUX2X1 U1774 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n2267), .Y(n2103) );
  MUX2X1 U1775 ( .B(n2102), .A(n2099), .S(n2226), .Y(n2113) );
  MUX2X1 U1776 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n2267), .Y(n2107) );
  MUX2X1 U1777 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n2267), .Y(n2106) );
  MUX2X1 U1778 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n2267), .Y(n2110) );
  MUX2X1 U1779 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n2267), .Y(n2109) );
  MUX2X1 U1780 ( .B(n2108), .A(n2105), .S(n2226), .Y(n2112) );
  MUX2X1 U1781 ( .B(n2111), .A(n2096), .S(n2220), .Y(n2216) );
  MUX2X1 U1782 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n2268), .Y(n2116) );
  MUX2X1 U1783 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n2268), .Y(n2115) );
  MUX2X1 U1784 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n2268), .Y(n2119) );
  MUX2X1 U1785 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n2268), .Y(n2118) );
  MUX2X1 U1786 ( .B(n2117), .A(n2114), .S(n2226), .Y(n2128) );
  MUX2X1 U1787 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n2268), .Y(n2122) );
  MUX2X1 U1788 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n2268), .Y(n2121) );
  MUX2X1 U1789 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n2268), .Y(n2125) );
  MUX2X1 U1790 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n2268), .Y(n2124) );
  MUX2X1 U1791 ( .B(n2123), .A(n2120), .S(n2226), .Y(n2127) );
  MUX2X1 U1792 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n2268), .Y(n2131) );
  MUX2X1 U1793 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n2268), .Y(n2130) );
  MUX2X1 U1794 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n2268), .Y(n2134) );
  MUX2X1 U1795 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n2268), .Y(n2133) );
  MUX2X1 U1796 ( .B(n2132), .A(n2129), .S(n2226), .Y(n2143) );
  MUX2X1 U1797 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n2269), .Y(n2137) );
  MUX2X1 U1798 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n2269), .Y(n2136) );
  MUX2X1 U1799 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n2269), .Y(n2140) );
  MUX2X1 U1800 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n2269), .Y(n2139) );
  MUX2X1 U1801 ( .B(n2138), .A(n2135), .S(n2226), .Y(n2142) );
  MUX2X1 U1802 ( .B(n2141), .A(n2126), .S(n2220), .Y(n2217) );
  MUX2X1 U1803 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n2269), .Y(n2146) );
  MUX2X1 U1804 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n2269), .Y(n2145) );
  MUX2X1 U1805 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n2269), .Y(n2149) );
  MUX2X1 U1806 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n2269), .Y(n2148) );
  MUX2X1 U1807 ( .B(n2147), .A(n2144), .S(n2226), .Y(n2158) );
  MUX2X1 U1808 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n2269), .Y(n2152) );
  MUX2X1 U1809 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n2269), .Y(n2151) );
  MUX2X1 U1810 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n2269), .Y(n2155) );
  MUX2X1 U1811 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n2269), .Y(n2154) );
  MUX2X1 U1812 ( .B(n2153), .A(n2150), .S(n2226), .Y(n2157) );
  MUX2X1 U1813 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n2270), .Y(n2161) );
  MUX2X1 U1814 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n2270), .Y(n2160) );
  MUX2X1 U1815 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n2270), .Y(n2164) );
  MUX2X1 U1816 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n2270), .Y(n2163) );
  MUX2X1 U1817 ( .B(n2162), .A(n2159), .S(n2226), .Y(n2173) );
  MUX2X1 U1818 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n2270), .Y(n2167) );
  MUX2X1 U1819 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n2270), .Y(n2166) );
  MUX2X1 U1820 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n2270), .Y(n2170) );
  MUX2X1 U1821 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n2270), .Y(n2169) );
  MUX2X1 U1822 ( .B(n2168), .A(n2165), .S(n2226), .Y(n2172) );
  MUX2X1 U1823 ( .B(n2171), .A(n2156), .S(n2220), .Y(n2218) );
  MUX2X1 U1824 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n2270), .Y(n2176) );
  MUX2X1 U1825 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n2270), .Y(n2175) );
  MUX2X1 U1826 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n2270), .Y(n2179) );
  MUX2X1 U1827 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n2270), .Y(n2178) );
  MUX2X1 U1828 ( .B(n2177), .A(n2174), .S(n2225), .Y(n2188) );
  MUX2X1 U1829 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n2271), .Y(n2182) );
  MUX2X1 U1830 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n2271), .Y(n2181) );
  MUX2X1 U1831 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n2271), .Y(n2185) );
  MUX2X1 U1832 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n2271), .Y(n2184) );
  MUX2X1 U1833 ( .B(n2183), .A(n2180), .S(n2225), .Y(n2187) );
  MUX2X1 U1834 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n2271), .Y(n2191) );
  MUX2X1 U1835 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n2271), .Y(n2190) );
  MUX2X1 U1836 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n2271), .Y(n2194) );
  MUX2X1 U1837 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n2271), .Y(n2193) );
  MUX2X1 U1838 ( .B(n2192), .A(n2189), .S(n2225), .Y(n2203) );
  MUX2X1 U1839 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n2271), .Y(n2197) );
  MUX2X1 U1840 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n2271), .Y(n2196) );
  MUX2X1 U1841 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n2271), .Y(n2200) );
  MUX2X1 U1842 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n2271), .Y(n2199) );
  MUX2X1 U1843 ( .B(n2198), .A(n2195), .S(n2225), .Y(n2202) );
  MUX2X1 U1844 ( .B(n2201), .A(n2186), .S(n2220), .Y(n2219) );
  INVX8 U1845 ( .A(n2242), .Y(n2231) );
  INVX8 U1846 ( .A(n2231), .Y(n2233) );
  INVX8 U1847 ( .A(n2273), .Y(n2243) );
  INVX8 U1848 ( .A(n2273), .Y(n2244) );
  INVX8 U1849 ( .A(n2273), .Y(n2245) );
  INVX8 U1850 ( .A(n2273), .Y(n2246) );
  INVX8 U1851 ( .A(n2274), .Y(n2247) );
  INVX8 U1852 ( .A(n2274), .Y(n2248) );
  INVX8 U1853 ( .A(n2274), .Y(n2249) );
  INVX8 U1854 ( .A(n2249), .Y(n2250) );
  INVX8 U1855 ( .A(n2249), .Y(n2251) );
  INVX8 U1856 ( .A(n2249), .Y(n2252) );
  INVX8 U1857 ( .A(n2248), .Y(n2253) );
  INVX8 U1858 ( .A(n2248), .Y(n2254) );
  INVX8 U1859 ( .A(n2248), .Y(n2255) );
  INVX8 U1860 ( .A(n2247), .Y(n2256) );
  INVX8 U1861 ( .A(n2247), .Y(n2257) );
  INVX8 U1862 ( .A(n2247), .Y(n2258) );
  INVX8 U1863 ( .A(n2246), .Y(n2259) );
  INVX8 U1864 ( .A(n2246), .Y(n2260) );
  INVX8 U1865 ( .A(n2246), .Y(n2261) );
  INVX8 U1866 ( .A(n2245), .Y(n2262) );
  INVX8 U1867 ( .A(n2245), .Y(n2263) );
  INVX8 U1868 ( .A(n2245), .Y(n2264) );
  INVX8 U1869 ( .A(n2244), .Y(n2265) );
  INVX8 U1870 ( .A(n2244), .Y(n2266) );
  INVX8 U1871 ( .A(n2244), .Y(n2267) );
  INVX8 U1872 ( .A(n2243), .Y(n2268) );
  INVX8 U1873 ( .A(n2243), .Y(n2269) );
  INVX8 U1874 ( .A(n2243), .Y(n2270) );
  INVX8 U1875 ( .A(n2243), .Y(n2271) );
  INVX8 U1876 ( .A(n2272), .Y(n2274) );
  AND2X2 U1877 ( .A(n3), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U1878 ( .A(N25), .B(n3), .Y(\data_out<7> ) );
  AND2X2 U1879 ( .A(N24), .B(n110), .Y(\data_out<8> ) );
  AND2X2 U1880 ( .A(n110), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U1881 ( .A(N22), .B(n109), .Y(\data_out<10> ) );
  AND2X2 U1882 ( .A(n1), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U1883 ( .A(n1), .B(N20), .Y(\data_out<12> ) );
  INVX1 U1884 ( .A(N11), .Y(n2378) );
  INVX1 U1885 ( .A(N10), .Y(n2377) );
  INVX8 U1886 ( .A(n2341), .Y(n2339) );
  INVX8 U1887 ( .A(n2341), .Y(n2340) );
  INVX8 U1888 ( .A(n37), .Y(n2343) );
  INVX8 U1889 ( .A(n38), .Y(n2345) );
  INVX8 U1890 ( .A(n39), .Y(n2347) );
  INVX8 U1891 ( .A(n40), .Y(n2349) );
  INVX8 U1892 ( .A(n41), .Y(n2351) );
  INVX8 U1893 ( .A(n42), .Y(n2353) );
  INVX8 U1894 ( .A(n43), .Y(n2355) );
  INVX8 U1895 ( .A(n44), .Y(n2357) );
  INVX8 U1896 ( .A(n45), .Y(n2359) );
  INVX8 U1897 ( .A(n46), .Y(n2361) );
  INVX8 U1898 ( .A(n47), .Y(n2363) );
  INVX8 U1899 ( .A(n48), .Y(n2365) );
  INVX8 U1900 ( .A(n49), .Y(n2367) );
  INVX8 U1901 ( .A(n50), .Y(n2369) );
  INVX8 U1902 ( .A(n51), .Y(n2371) );
  INVX8 U1903 ( .A(n52), .Y(n2373) );
  AND2X2 U1904 ( .A(n110), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U1905 ( .A(N30), .B(n2), .Y(\data_out<2> ) );
  AND2X2 U1906 ( .A(N29), .B(n112), .Y(\data_out<3> ) );
  AND2X2 U1907 ( .A(N28), .B(n114), .Y(\data_out<4> ) );
  AND2X2 U1908 ( .A(N27), .B(n114), .Y(\data_out<5> ) );
  AND2X2 U1909 ( .A(n1), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U1910 ( .A(n112), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U1911 ( .A(N17), .B(n2), .Y(\data_out<15> ) );
  OAI21X1 U1912 ( .A(n2276), .B(n2343), .C(n184), .Y(n2911) );
  OAI21X1 U1913 ( .A(n2346), .B(n2275), .C(n186), .Y(n2910) );
  OAI21X1 U1914 ( .A(n2348), .B(n2275), .C(n188), .Y(n2909) );
  OAI21X1 U1915 ( .A(n2350), .B(n2275), .C(n190), .Y(n2908) );
  OAI21X1 U1916 ( .A(n2352), .B(n2275), .C(n192), .Y(n2907) );
  OAI21X1 U1917 ( .A(n2354), .B(n2275), .C(n194), .Y(n2906) );
  OAI21X1 U1918 ( .A(n2356), .B(n2275), .C(n196), .Y(n2905) );
  OAI21X1 U1919 ( .A(n2358), .B(n2275), .C(n198), .Y(n2904) );
  OAI21X1 U1920 ( .A(n2360), .B(n2275), .C(n200), .Y(n2903) );
  OAI21X1 U1921 ( .A(n2362), .B(n2276), .C(n202), .Y(n2902) );
  OAI21X1 U1922 ( .A(n2364), .B(n2276), .C(n204), .Y(n2901) );
  OAI21X1 U1923 ( .A(n2366), .B(n2276), .C(n206), .Y(n2900) );
  OAI21X1 U1924 ( .A(n2368), .B(n2276), .C(n208), .Y(n2899) );
  OAI21X1 U1925 ( .A(n2370), .B(n2276), .C(n210), .Y(n2898) );
  OAI21X1 U1926 ( .A(n2372), .B(n2276), .C(n212), .Y(n2897) );
  OAI21X1 U1927 ( .A(n2374), .B(n2276), .C(n215), .Y(n2896) );
  OAI21X1 U1928 ( .A(n2277), .B(n2343), .C(n32), .Y(n2895) );
  OAI21X1 U1929 ( .A(n2277), .B(n2346), .C(n217), .Y(n2894) );
  OAI21X1 U1930 ( .A(n2277), .B(n2348), .C(n219), .Y(n2893) );
  OAI21X1 U1931 ( .A(n2277), .B(n2350), .C(n221), .Y(n2892) );
  OAI21X1 U1932 ( .A(n2277), .B(n2352), .C(n223), .Y(n2891) );
  OAI21X1 U1933 ( .A(n2277), .B(n2354), .C(n225), .Y(n2890) );
  OAI21X1 U1934 ( .A(n2277), .B(n2356), .C(n227), .Y(n2889) );
  OAI21X1 U1935 ( .A(n2277), .B(n2358), .C(n229), .Y(n2888) );
  OAI21X1 U1936 ( .A(n2278), .B(n2360), .C(n231), .Y(n2887) );
  OAI21X1 U1937 ( .A(n2278), .B(n2362), .C(n233), .Y(n2886) );
  OAI21X1 U1938 ( .A(n2278), .B(n2364), .C(n235), .Y(n2885) );
  OAI21X1 U1939 ( .A(n2278), .B(n2366), .C(n237), .Y(n2884) );
  OAI21X1 U1940 ( .A(n2278), .B(n2368), .C(n239), .Y(n2883) );
  OAI21X1 U1941 ( .A(n2278), .B(n2370), .C(n241), .Y(n2882) );
  OAI21X1 U1942 ( .A(n2278), .B(n2372), .C(n243), .Y(n2881) );
  OAI21X1 U1943 ( .A(n2278), .B(n2374), .C(n245), .Y(n2880) );
  NAND3X1 U1944 ( .A(n2376), .B(n2379), .C(n2378), .Y(n2385) );
  OAI21X1 U1945 ( .A(n2279), .B(n2344), .C(n34), .Y(n2879) );
  OAI21X1 U1946 ( .A(n2279), .B(n2346), .C(n247), .Y(n2878) );
  OAI21X1 U1947 ( .A(n2279), .B(n2348), .C(n249), .Y(n2877) );
  OAI21X1 U1948 ( .A(n2279), .B(n2350), .C(n251), .Y(n2876) );
  OAI21X1 U1949 ( .A(n2279), .B(n2352), .C(n253), .Y(n2875) );
  OAI21X1 U1950 ( .A(n2279), .B(n2354), .C(n255), .Y(n2874) );
  OAI21X1 U1951 ( .A(n2279), .B(n2356), .C(n257), .Y(n2873) );
  OAI21X1 U1952 ( .A(n2279), .B(n2358), .C(n259), .Y(n2872) );
  OAI21X1 U1953 ( .A(n2280), .B(n2360), .C(n261), .Y(n2871) );
  OAI21X1 U1954 ( .A(n2280), .B(n2362), .C(n263), .Y(n2870) );
  OAI21X1 U1955 ( .A(n2280), .B(n2364), .C(n265), .Y(n2869) );
  OAI21X1 U1956 ( .A(n2280), .B(n2366), .C(n267), .Y(n2868) );
  OAI21X1 U1957 ( .A(n2280), .B(n2368), .C(n269), .Y(n2867) );
  OAI21X1 U1958 ( .A(n2280), .B(n2370), .C(n271), .Y(n2866) );
  OAI21X1 U1959 ( .A(n2280), .B(n2372), .C(n273), .Y(n2865) );
  OAI21X1 U1960 ( .A(n2280), .B(n2374), .C(n275), .Y(n2864) );
  NAND3X1 U1961 ( .A(n2379), .B(n2378), .C(n2377), .Y(n2386) );
  OAI21X1 U1962 ( .A(n2281), .B(n2343), .C(n36), .Y(n2863) );
  OAI21X1 U1963 ( .A(n2281), .B(n2346), .C(n277), .Y(n2862) );
  OAI21X1 U1964 ( .A(n2281), .B(n2348), .C(n279), .Y(n2861) );
  OAI21X1 U1965 ( .A(n2281), .B(n2350), .C(n281), .Y(n2860) );
  OAI21X1 U1966 ( .A(n2281), .B(n2352), .C(n283), .Y(n2859) );
  OAI21X1 U1967 ( .A(n2281), .B(n2354), .C(n285), .Y(n2858) );
  OAI21X1 U1968 ( .A(n2281), .B(n2356), .C(n287), .Y(n2857) );
  OAI21X1 U1969 ( .A(n2281), .B(n2358), .C(n289), .Y(n2856) );
  OAI21X1 U1970 ( .A(n2282), .B(n2360), .C(n291), .Y(n2855) );
  OAI21X1 U1971 ( .A(n2282), .B(n2362), .C(n293), .Y(n2854) );
  OAI21X1 U1972 ( .A(n2282), .B(n2364), .C(n295), .Y(n2853) );
  OAI21X1 U1973 ( .A(n2282), .B(n2366), .C(n297), .Y(n2852) );
  OAI21X1 U1974 ( .A(n2282), .B(n2368), .C(n299), .Y(n2851) );
  OAI21X1 U1975 ( .A(n2282), .B(n2370), .C(n301), .Y(n2850) );
  OAI21X1 U1976 ( .A(n2282), .B(n2372), .C(n303), .Y(n2849) );
  OAI21X1 U1977 ( .A(n2282), .B(n2374), .C(n305), .Y(n2848) );
  NAND3X1 U1978 ( .A(n2376), .B(n2233), .C(n2380), .Y(n2387) );
  OAI21X1 U1979 ( .A(n2283), .B(n2343), .C(n307), .Y(n2847) );
  OAI21X1 U1980 ( .A(n2283), .B(n2346), .C(n309), .Y(n2846) );
  OAI21X1 U1981 ( .A(n2283), .B(n2348), .C(n311), .Y(n2845) );
  OAI21X1 U1982 ( .A(n2283), .B(n2350), .C(n313), .Y(n2844) );
  OAI21X1 U1983 ( .A(n2283), .B(n2352), .C(n315), .Y(n2843) );
  OAI21X1 U1984 ( .A(n2283), .B(n2354), .C(n317), .Y(n2842) );
  OAI21X1 U1985 ( .A(n2283), .B(n2356), .C(n319), .Y(n2841) );
  OAI21X1 U1986 ( .A(n2283), .B(n2358), .C(n321), .Y(n2840) );
  OAI21X1 U1987 ( .A(n2284), .B(n2360), .C(n323), .Y(n2839) );
  OAI21X1 U1988 ( .A(n2284), .B(n2362), .C(n325), .Y(n2838) );
  OAI21X1 U1989 ( .A(n2284), .B(n2364), .C(n327), .Y(n2837) );
  OAI21X1 U1990 ( .A(n2284), .B(n2366), .C(n329), .Y(n2836) );
  OAI21X1 U1991 ( .A(n2284), .B(n2368), .C(n331), .Y(n2835) );
  OAI21X1 U1992 ( .A(n2284), .B(n2370), .C(n333), .Y(n2834) );
  OAI21X1 U1993 ( .A(n2284), .B(n2372), .C(n335), .Y(n2833) );
  OAI21X1 U1994 ( .A(n2284), .B(n2374), .C(n337), .Y(n2832) );
  NAND3X1 U1995 ( .A(n2380), .B(n2233), .C(n2377), .Y(n2388) );
  OAI21X1 U1996 ( .A(n2285), .B(n2344), .C(n339), .Y(n2831) );
  OAI21X1 U1997 ( .A(n2285), .B(n2346), .C(n341), .Y(n2830) );
  OAI21X1 U1998 ( .A(n2285), .B(n2348), .C(n343), .Y(n2829) );
  OAI21X1 U1999 ( .A(n2285), .B(n2350), .C(n345), .Y(n2828) );
  OAI21X1 U2000 ( .A(n2285), .B(n2352), .C(n347), .Y(n2827) );
  OAI21X1 U2001 ( .A(n2285), .B(n2354), .C(n349), .Y(n2826) );
  OAI21X1 U2002 ( .A(n2285), .B(n2356), .C(n351), .Y(n2825) );
  OAI21X1 U2003 ( .A(n2285), .B(n2358), .C(n353), .Y(n2824) );
  OAI21X1 U2004 ( .A(n2286), .B(n2360), .C(n355), .Y(n2823) );
  OAI21X1 U2005 ( .A(n2286), .B(n2362), .C(n357), .Y(n2822) );
  OAI21X1 U2006 ( .A(n2286), .B(n2364), .C(n359), .Y(n2821) );
  OAI21X1 U2007 ( .A(n2286), .B(n2366), .C(n361), .Y(n2820) );
  OAI21X1 U2008 ( .A(n2286), .B(n2368), .C(n363), .Y(n2819) );
  OAI21X1 U2009 ( .A(n2286), .B(n2370), .C(n365), .Y(n2818) );
  OAI21X1 U2010 ( .A(n2286), .B(n2372), .C(n367), .Y(n2817) );
  OAI21X1 U2011 ( .A(n2286), .B(n2374), .C(n369), .Y(n2816) );
  NAND3X1 U2012 ( .A(n2376), .B(n2380), .C(n2378), .Y(n2389) );
  OAI21X1 U2013 ( .A(n2288), .B(n2343), .C(n371), .Y(n2815) );
  OAI21X1 U2014 ( .A(n2288), .B(n2346), .C(n373), .Y(n2814) );
  OAI21X1 U2015 ( .A(n2288), .B(n2348), .C(n375), .Y(n2813) );
  OAI21X1 U2016 ( .A(n2288), .B(n2350), .C(n377), .Y(n2812) );
  OAI21X1 U2017 ( .A(n2288), .B(n2352), .C(n379), .Y(n2811) );
  OAI21X1 U2018 ( .A(n2288), .B(n2354), .C(n381), .Y(n2810) );
  OAI21X1 U2019 ( .A(n2288), .B(n2356), .C(n383), .Y(n2809) );
  OAI21X1 U2020 ( .A(n2288), .B(n2358), .C(n385), .Y(n2808) );
  OAI21X1 U2021 ( .A(n2289), .B(n2360), .C(n387), .Y(n2807) );
  OAI21X1 U2022 ( .A(n2289), .B(n2362), .C(n389), .Y(n2806) );
  OAI21X1 U2023 ( .A(n2289), .B(n2364), .C(n391), .Y(n2805) );
  OAI21X1 U2024 ( .A(n2289), .B(n2366), .C(n393), .Y(n2804) );
  OAI21X1 U2025 ( .A(n2289), .B(n2368), .C(n395), .Y(n2803) );
  OAI21X1 U2026 ( .A(n2289), .B(n2370), .C(n397), .Y(n2802) );
  OAI21X1 U2027 ( .A(n2289), .B(n2372), .C(n399), .Y(n2801) );
  OAI21X1 U2028 ( .A(n2289), .B(n2374), .C(n401), .Y(n2800) );
  NOR3X1 U2029 ( .A(n2376), .B(n2233), .C(n2379), .Y(n2399) );
  OAI21X1 U2030 ( .A(n1662), .B(n2343), .C(n403), .Y(n2799) );
  OAI21X1 U2031 ( .A(n1662), .B(n2346), .C(n405), .Y(n2798) );
  OAI21X1 U2032 ( .A(n1662), .B(n2348), .C(n407), .Y(n2797) );
  OAI21X1 U2033 ( .A(n1662), .B(n2350), .C(n409), .Y(n2796) );
  OAI21X1 U2034 ( .A(n1662), .B(n2352), .C(n411), .Y(n2795) );
  OAI21X1 U2035 ( .A(n1662), .B(n2354), .C(n413), .Y(n2794) );
  OAI21X1 U2036 ( .A(n1662), .B(n2356), .C(n415), .Y(n2793) );
  OAI21X1 U2037 ( .A(n1662), .B(n2358), .C(n417), .Y(n2792) );
  OAI21X1 U2038 ( .A(n1662), .B(n2360), .C(n419), .Y(n2791) );
  OAI21X1 U2039 ( .A(n1662), .B(n2362), .C(n421), .Y(n2790) );
  OAI21X1 U2040 ( .A(n1662), .B(n2364), .C(n423), .Y(n2789) );
  OAI21X1 U2041 ( .A(n1662), .B(n2366), .C(n425), .Y(n2788) );
  OAI21X1 U2042 ( .A(n1662), .B(n2368), .C(n427), .Y(n2787) );
  OAI21X1 U2043 ( .A(n1662), .B(n2370), .C(n429), .Y(n2786) );
  OAI21X1 U2044 ( .A(n1662), .B(n2372), .C(n431), .Y(n2785) );
  OAI21X1 U2045 ( .A(n1662), .B(n2374), .C(n433), .Y(n2784) );
  OAI21X1 U2046 ( .A(n2290), .B(n2343), .C(n116), .Y(n2783) );
  OAI21X1 U2047 ( .A(n2290), .B(n2345), .C(n118), .Y(n2782) );
  OAI21X1 U2048 ( .A(n2290), .B(n2347), .C(n120), .Y(n2781) );
  OAI21X1 U2049 ( .A(n2290), .B(n2349), .C(n122), .Y(n2780) );
  OAI21X1 U2050 ( .A(n2290), .B(n2351), .C(n124), .Y(n2779) );
  OAI21X1 U2051 ( .A(n2290), .B(n2353), .C(n126), .Y(n2778) );
  OAI21X1 U2052 ( .A(n2290), .B(n2355), .C(n128), .Y(n2777) );
  OAI21X1 U2053 ( .A(n2290), .B(n2357), .C(n130), .Y(n2776) );
  OAI21X1 U2054 ( .A(n2291), .B(n2359), .C(n435), .Y(n2775) );
  OAI21X1 U2055 ( .A(n2291), .B(n2361), .C(n437), .Y(n2774) );
  OAI21X1 U2056 ( .A(n2291), .B(n2363), .C(n439), .Y(n2773) );
  OAI21X1 U2057 ( .A(n2291), .B(n2365), .C(n441), .Y(n2772) );
  OAI21X1 U2058 ( .A(n2291), .B(n2367), .C(n443), .Y(n2771) );
  OAI21X1 U2059 ( .A(n2291), .B(n2369), .C(n445), .Y(n2770) );
  OAI21X1 U2060 ( .A(n2291), .B(n2371), .C(n447), .Y(n2769) );
  OAI21X1 U2061 ( .A(n2291), .B(n2373), .C(n449), .Y(n2768) );
  OAI21X1 U2062 ( .A(n2292), .B(n2343), .C(n132), .Y(n2767) );
  OAI21X1 U2063 ( .A(n2292), .B(n2345), .C(n134), .Y(n2766) );
  OAI21X1 U2064 ( .A(n2292), .B(n2347), .C(n136), .Y(n2765) );
  OAI21X1 U2065 ( .A(n2292), .B(n2349), .C(n138), .Y(n2764) );
  OAI21X1 U2066 ( .A(n2292), .B(n2351), .C(n140), .Y(n2763) );
  OAI21X1 U2067 ( .A(n2292), .B(n2353), .C(n142), .Y(n2762) );
  OAI21X1 U2068 ( .A(n2292), .B(n2355), .C(n144), .Y(n2761) );
  OAI21X1 U2069 ( .A(n2292), .B(n2357), .C(n146), .Y(n2760) );
  OAI21X1 U2070 ( .A(n2293), .B(n2359), .C(n451), .Y(n2759) );
  OAI21X1 U2071 ( .A(n2293), .B(n2361), .C(n453), .Y(n2758) );
  OAI21X1 U2072 ( .A(n2293), .B(n2363), .C(n455), .Y(n2757) );
  OAI21X1 U2073 ( .A(n2293), .B(n2365), .C(n457), .Y(n2756) );
  OAI21X1 U2074 ( .A(n2293), .B(n2367), .C(n459), .Y(n2755) );
  OAI21X1 U2075 ( .A(n2293), .B(n2369), .C(n461), .Y(n2754) );
  OAI21X1 U2076 ( .A(n2293), .B(n2371), .C(n463), .Y(n2753) );
  OAI21X1 U2077 ( .A(n2293), .B(n2373), .C(n465), .Y(n2752) );
  OAI21X1 U2078 ( .A(n2295), .B(n2343), .C(n148), .Y(n2751) );
  OAI21X1 U2079 ( .A(n2295), .B(n2345), .C(n150), .Y(n2750) );
  OAI21X1 U2080 ( .A(n2295), .B(n2347), .C(n152), .Y(n2749) );
  OAI21X1 U2081 ( .A(n2295), .B(n2349), .C(n154), .Y(n2748) );
  OAI21X1 U2082 ( .A(n2295), .B(n2351), .C(n156), .Y(n2747) );
  OAI21X1 U2083 ( .A(n2295), .B(n2353), .C(n158), .Y(n2746) );
  OAI21X1 U2084 ( .A(n2295), .B(n2355), .C(n160), .Y(n2745) );
  OAI21X1 U2085 ( .A(n2295), .B(n2357), .C(n162), .Y(n2744) );
  OAI21X1 U2086 ( .A(n2296), .B(n2359), .C(n467), .Y(n2743) );
  OAI21X1 U2087 ( .A(n2296), .B(n2361), .C(n469), .Y(n2742) );
  OAI21X1 U2088 ( .A(n2296), .B(n2363), .C(n471), .Y(n2741) );
  OAI21X1 U2089 ( .A(n2296), .B(n2365), .C(n473), .Y(n2740) );
  OAI21X1 U2090 ( .A(n2296), .B(n2367), .C(n475), .Y(n2739) );
  OAI21X1 U2091 ( .A(n2296), .B(n2369), .C(n477), .Y(n2738) );
  OAI21X1 U2092 ( .A(n2296), .B(n2371), .C(n479), .Y(n2737) );
  OAI21X1 U2093 ( .A(n2296), .B(n2373), .C(n481), .Y(n2736) );
  OAI21X1 U2094 ( .A(n2297), .B(n2343), .C(n164), .Y(n2735) );
  OAI21X1 U2095 ( .A(n2297), .B(n2345), .C(n166), .Y(n2734) );
  OAI21X1 U2096 ( .A(n2297), .B(n2347), .C(n168), .Y(n2733) );
  OAI21X1 U2097 ( .A(n2297), .B(n2349), .C(n170), .Y(n2732) );
  OAI21X1 U2098 ( .A(n2297), .B(n2351), .C(n172), .Y(n2731) );
  OAI21X1 U2099 ( .A(n2297), .B(n2353), .C(n174), .Y(n2730) );
  OAI21X1 U2100 ( .A(n2297), .B(n2355), .C(n176), .Y(n2729) );
  OAI21X1 U2101 ( .A(n2297), .B(n2357), .C(n178), .Y(n2728) );
  OAI21X1 U2102 ( .A(n2298), .B(n2359), .C(n483), .Y(n2727) );
  OAI21X1 U2103 ( .A(n2298), .B(n2361), .C(n485), .Y(n2726) );
  OAI21X1 U2104 ( .A(n2298), .B(n2363), .C(n487), .Y(n2725) );
  OAI21X1 U2105 ( .A(n2298), .B(n2365), .C(n489), .Y(n2724) );
  OAI21X1 U2106 ( .A(n2298), .B(n2367), .C(n491), .Y(n2723) );
  OAI21X1 U2107 ( .A(n2298), .B(n2369), .C(n493), .Y(n2722) );
  OAI21X1 U2108 ( .A(n2298), .B(n2371), .C(n495), .Y(n2721) );
  OAI21X1 U2109 ( .A(n2298), .B(n2373), .C(n497), .Y(n2720) );
  OAI21X1 U2110 ( .A(n2300), .B(n2343), .C(n499), .Y(n2719) );
  OAI21X1 U2111 ( .A(n2300), .B(n2345), .C(n501), .Y(n2718) );
  OAI21X1 U2112 ( .A(n2300), .B(n2347), .C(n503), .Y(n2717) );
  OAI21X1 U2113 ( .A(n2300), .B(n2349), .C(n505), .Y(n2716) );
  OAI21X1 U2114 ( .A(n2300), .B(n2351), .C(n507), .Y(n2715) );
  OAI21X1 U2115 ( .A(n2300), .B(n2353), .C(n509), .Y(n2714) );
  OAI21X1 U2116 ( .A(n2300), .B(n2355), .C(n511), .Y(n2713) );
  OAI21X1 U2117 ( .A(n2300), .B(n2357), .C(n513), .Y(n2712) );
  OAI21X1 U2118 ( .A(n2301), .B(n2359), .C(n515), .Y(n2711) );
  OAI21X1 U2119 ( .A(n2301), .B(n2361), .C(n517), .Y(n2710) );
  OAI21X1 U2120 ( .A(n2301), .B(n2363), .C(n519), .Y(n2709) );
  OAI21X1 U2121 ( .A(n2301), .B(n2365), .C(n521), .Y(n2708) );
  OAI21X1 U2122 ( .A(n2301), .B(n2367), .C(n523), .Y(n2707) );
  OAI21X1 U2123 ( .A(n2301), .B(n2369), .C(n525), .Y(n2706) );
  OAI21X1 U2124 ( .A(n2301), .B(n2371), .C(n527), .Y(n2705) );
  OAI21X1 U2125 ( .A(n2301), .B(n2373), .C(n529), .Y(n2704) );
  OAI21X1 U2126 ( .A(n2303), .B(n2343), .C(n531), .Y(n2703) );
  OAI21X1 U2127 ( .A(n2303), .B(n2345), .C(n533), .Y(n2702) );
  OAI21X1 U2128 ( .A(n2303), .B(n2347), .C(n535), .Y(n2701) );
  OAI21X1 U2129 ( .A(n2303), .B(n2349), .C(n537), .Y(n2700) );
  OAI21X1 U2130 ( .A(n2303), .B(n2351), .C(n539), .Y(n2699) );
  OAI21X1 U2131 ( .A(n2303), .B(n2353), .C(n541), .Y(n2698) );
  OAI21X1 U2132 ( .A(n2303), .B(n2355), .C(n543), .Y(n2697) );
  OAI21X1 U2133 ( .A(n2303), .B(n2357), .C(n545), .Y(n2696) );
  OAI21X1 U2134 ( .A(n2304), .B(n2359), .C(n547), .Y(n2695) );
  OAI21X1 U2135 ( .A(n2304), .B(n2361), .C(n549), .Y(n2694) );
  OAI21X1 U2136 ( .A(n2304), .B(n2363), .C(n551), .Y(n2693) );
  OAI21X1 U2137 ( .A(n2304), .B(n2365), .C(n553), .Y(n2692) );
  OAI21X1 U2138 ( .A(n2304), .B(n2367), .C(n555), .Y(n2691) );
  OAI21X1 U2139 ( .A(n2304), .B(n2369), .C(n557), .Y(n2690) );
  OAI21X1 U2140 ( .A(n2304), .B(n2371), .C(n559), .Y(n2689) );
  OAI21X1 U2141 ( .A(n2304), .B(n2373), .C(n561), .Y(n2688) );
  OAI21X1 U2142 ( .A(n2305), .B(n2343), .C(n563), .Y(n2687) );
  OAI21X1 U2143 ( .A(n2305), .B(n2345), .C(n565), .Y(n2686) );
  OAI21X1 U2144 ( .A(n2305), .B(n2347), .C(n567), .Y(n2685) );
  OAI21X1 U2145 ( .A(n2305), .B(n2349), .C(n569), .Y(n2684) );
  OAI21X1 U2146 ( .A(n2305), .B(n2351), .C(n571), .Y(n2683) );
  OAI21X1 U2147 ( .A(n2305), .B(n2353), .C(n573), .Y(n2682) );
  OAI21X1 U2148 ( .A(n2305), .B(n2355), .C(n575), .Y(n2681) );
  OAI21X1 U2149 ( .A(n2305), .B(n2357), .C(n577), .Y(n2680) );
  OAI21X1 U2150 ( .A(n2306), .B(n2359), .C(n579), .Y(n2679) );
  OAI21X1 U2151 ( .A(n2306), .B(n2361), .C(n581), .Y(n2678) );
  OAI21X1 U2152 ( .A(n2306), .B(n2363), .C(n583), .Y(n2677) );
  OAI21X1 U2153 ( .A(n2306), .B(n2365), .C(n585), .Y(n2676) );
  OAI21X1 U2154 ( .A(n2306), .B(n2367), .C(n587), .Y(n2675) );
  OAI21X1 U2155 ( .A(n2306), .B(n2369), .C(n589), .Y(n2674) );
  OAI21X1 U2156 ( .A(n2306), .B(n2371), .C(n591), .Y(n2673) );
  OAI21X1 U2157 ( .A(n2306), .B(n2373), .C(n593), .Y(n2672) );
  OAI21X1 U2158 ( .A(n2307), .B(n2343), .C(n595), .Y(n2671) );
  OAI21X1 U2159 ( .A(n2307), .B(n2345), .C(n597), .Y(n2670) );
  OAI21X1 U2160 ( .A(n2307), .B(n2347), .C(n599), .Y(n2669) );
  OAI21X1 U2161 ( .A(n2307), .B(n2349), .C(n601), .Y(n2668) );
  OAI21X1 U2162 ( .A(n2307), .B(n2351), .C(n603), .Y(n2667) );
  OAI21X1 U2163 ( .A(n2307), .B(n2353), .C(n605), .Y(n2666) );
  OAI21X1 U2164 ( .A(n2307), .B(n2355), .C(n607), .Y(n2665) );
  OAI21X1 U2165 ( .A(n2307), .B(n2357), .C(n609), .Y(n2664) );
  OAI21X1 U2166 ( .A(n2307), .B(n2359), .C(n611), .Y(n2663) );
  OAI21X1 U2167 ( .A(n2307), .B(n2361), .C(n613), .Y(n2662) );
  OAI21X1 U2168 ( .A(n2307), .B(n2363), .C(n615), .Y(n2661) );
  OAI21X1 U2169 ( .A(n2307), .B(n2365), .C(n617), .Y(n2660) );
  OAI21X1 U2170 ( .A(n2307), .B(n2367), .C(n619), .Y(n2659) );
  OAI21X1 U2171 ( .A(n2307), .B(n2369), .C(n621), .Y(n2658) );
  OAI21X1 U2172 ( .A(n2307), .B(n2371), .C(n623), .Y(n2657) );
  OAI21X1 U2173 ( .A(n2307), .B(n2373), .C(n625), .Y(n2656) );
  NAND3X1 U2174 ( .A(n2381), .B(n2912), .C(n2384), .Y(n2390) );
  OAI21X1 U2175 ( .A(n2308), .B(n2343), .C(n627), .Y(n2655) );
  OAI21X1 U2176 ( .A(n2308), .B(n2345), .C(n629), .Y(n2654) );
  OAI21X1 U2177 ( .A(n2308), .B(n2347), .C(n631), .Y(n2653) );
  OAI21X1 U2178 ( .A(n2308), .B(n2349), .C(n633), .Y(n2652) );
  OAI21X1 U2179 ( .A(n2308), .B(n2351), .C(n635), .Y(n2651) );
  OAI21X1 U2180 ( .A(n2308), .B(n2353), .C(n637), .Y(n2650) );
  OAI21X1 U2181 ( .A(n2308), .B(n2355), .C(n639), .Y(n2649) );
  OAI21X1 U2182 ( .A(n2308), .B(n2357), .C(n641), .Y(n2648) );
  OAI21X1 U2183 ( .A(n2309), .B(n2359), .C(n643), .Y(n2647) );
  OAI21X1 U2184 ( .A(n2309), .B(n2361), .C(n645), .Y(n2646) );
  OAI21X1 U2185 ( .A(n2309), .B(n2363), .C(n647), .Y(n2645) );
  OAI21X1 U2186 ( .A(n2309), .B(n2365), .C(n649), .Y(n2644) );
  OAI21X1 U2187 ( .A(n2309), .B(n2367), .C(n1163), .Y(n2643) );
  OAI21X1 U2188 ( .A(n2309), .B(n2369), .C(n1165), .Y(n2642) );
  OAI21X1 U2189 ( .A(n2309), .B(n2371), .C(n1167), .Y(n2641) );
  OAI21X1 U2190 ( .A(n2309), .B(n2373), .C(n1169), .Y(n2640) );
  OAI21X1 U2191 ( .A(n2310), .B(n2343), .C(n1171), .Y(n2639) );
  OAI21X1 U2192 ( .A(n2310), .B(n2345), .C(n1173), .Y(n2638) );
  OAI21X1 U2193 ( .A(n2310), .B(n2347), .C(n1175), .Y(n2637) );
  OAI21X1 U2194 ( .A(n2310), .B(n2349), .C(n1177), .Y(n2636) );
  OAI21X1 U2195 ( .A(n2310), .B(n2351), .C(n1179), .Y(n2635) );
  OAI21X1 U2196 ( .A(n2310), .B(n2353), .C(n1181), .Y(n2634) );
  OAI21X1 U2197 ( .A(n2310), .B(n2355), .C(n1183), .Y(n2633) );
  OAI21X1 U2198 ( .A(n2310), .B(n2357), .C(n1185), .Y(n2632) );
  OAI21X1 U2199 ( .A(n2311), .B(n2359), .C(n1187), .Y(n2631) );
  OAI21X1 U2200 ( .A(n2311), .B(n2361), .C(n1189), .Y(n2630) );
  OAI21X1 U2201 ( .A(n2311), .B(n2363), .C(n1191), .Y(n2629) );
  OAI21X1 U2202 ( .A(n2311), .B(n2365), .C(n1193), .Y(n2628) );
  OAI21X1 U2203 ( .A(n2311), .B(n2367), .C(n1195), .Y(n2627) );
  OAI21X1 U2204 ( .A(n2311), .B(n2369), .C(n1197), .Y(n2626) );
  OAI21X1 U2205 ( .A(n2311), .B(n2371), .C(n1199), .Y(n2625) );
  OAI21X1 U2206 ( .A(n2311), .B(n2373), .C(n1201), .Y(n2624) );
  OAI21X1 U2207 ( .A(n2312), .B(n2343), .C(n1203), .Y(n2623) );
  OAI21X1 U2208 ( .A(n2312), .B(n2345), .C(n1205), .Y(n2622) );
  OAI21X1 U2209 ( .A(n2312), .B(n2347), .C(n1207), .Y(n2621) );
  OAI21X1 U2210 ( .A(n2312), .B(n2349), .C(n1209), .Y(n2620) );
  OAI21X1 U2211 ( .A(n2312), .B(n2351), .C(n1211), .Y(n2619) );
  OAI21X1 U2212 ( .A(n2312), .B(n2353), .C(n1213), .Y(n2618) );
  OAI21X1 U2213 ( .A(n2312), .B(n2355), .C(n1215), .Y(n2617) );
  OAI21X1 U2214 ( .A(n2312), .B(n2357), .C(n1217), .Y(n2616) );
  OAI21X1 U2215 ( .A(n2313), .B(n2359), .C(n1219), .Y(n2615) );
  OAI21X1 U2216 ( .A(n2313), .B(n2361), .C(n1221), .Y(n2614) );
  OAI21X1 U2217 ( .A(n2313), .B(n2363), .C(n1223), .Y(n2613) );
  OAI21X1 U2218 ( .A(n2313), .B(n2365), .C(n1225), .Y(n2612) );
  OAI21X1 U2219 ( .A(n2313), .B(n2367), .C(n1227), .Y(n2611) );
  OAI21X1 U2220 ( .A(n2313), .B(n2369), .C(n1229), .Y(n2610) );
  OAI21X1 U2221 ( .A(n2313), .B(n2371), .C(n1231), .Y(n2609) );
  OAI21X1 U2222 ( .A(n2313), .B(n2373), .C(n1233), .Y(n2608) );
  OAI21X1 U2223 ( .A(n2314), .B(n2343), .C(n1235), .Y(n2607) );
  OAI21X1 U2224 ( .A(n2314), .B(n2345), .C(n1237), .Y(n2606) );
  OAI21X1 U2225 ( .A(n2314), .B(n2347), .C(n1239), .Y(n2605) );
  OAI21X1 U2226 ( .A(n2314), .B(n2349), .C(n1241), .Y(n2604) );
  OAI21X1 U2227 ( .A(n2314), .B(n2351), .C(n1243), .Y(n2603) );
  OAI21X1 U2228 ( .A(n2314), .B(n2353), .C(n1245), .Y(n2602) );
  OAI21X1 U2229 ( .A(n2314), .B(n2355), .C(n1247), .Y(n2601) );
  OAI21X1 U2230 ( .A(n2314), .B(n2357), .C(n1249), .Y(n2600) );
  OAI21X1 U2231 ( .A(n2315), .B(n2359), .C(n1251), .Y(n2599) );
  OAI21X1 U2232 ( .A(n2315), .B(n2361), .C(n1253), .Y(n2598) );
  OAI21X1 U2233 ( .A(n2315), .B(n2363), .C(n1255), .Y(n2597) );
  OAI21X1 U2234 ( .A(n2315), .B(n2365), .C(n1257), .Y(n2596) );
  OAI21X1 U2235 ( .A(n2315), .B(n2367), .C(n1259), .Y(n2595) );
  OAI21X1 U2236 ( .A(n2315), .B(n2369), .C(n1261), .Y(n2594) );
  OAI21X1 U2237 ( .A(n2315), .B(n2371), .C(n1263), .Y(n2593) );
  OAI21X1 U2238 ( .A(n2315), .B(n2373), .C(n1265), .Y(n2592) );
  OAI21X1 U2239 ( .A(n2316), .B(n2343), .C(n1267), .Y(n2591) );
  OAI21X1 U2240 ( .A(n2316), .B(n2345), .C(n1269), .Y(n2590) );
  OAI21X1 U2241 ( .A(n2316), .B(n2347), .C(n1271), .Y(n2589) );
  OAI21X1 U2242 ( .A(n2316), .B(n2349), .C(n1273), .Y(n2588) );
  OAI21X1 U2243 ( .A(n2316), .B(n2351), .C(n1275), .Y(n2587) );
  OAI21X1 U2244 ( .A(n2316), .B(n2353), .C(n1277), .Y(n2586) );
  OAI21X1 U2245 ( .A(n2316), .B(n2355), .C(n1279), .Y(n2585) );
  OAI21X1 U2246 ( .A(n2316), .B(n2357), .C(n1281), .Y(n2584) );
  OAI21X1 U2247 ( .A(n2317), .B(n2359), .C(n1283), .Y(n2583) );
  OAI21X1 U2248 ( .A(n2317), .B(n2361), .C(n1285), .Y(n2582) );
  OAI21X1 U2249 ( .A(n2317), .B(n2363), .C(n1287), .Y(n2581) );
  OAI21X1 U2250 ( .A(n2317), .B(n2365), .C(n1289), .Y(n2580) );
  OAI21X1 U2251 ( .A(n2317), .B(n2367), .C(n1291), .Y(n2579) );
  OAI21X1 U2252 ( .A(n2317), .B(n2369), .C(n1293), .Y(n2578) );
  OAI21X1 U2253 ( .A(n2317), .B(n2371), .C(n1295), .Y(n2577) );
  OAI21X1 U2254 ( .A(n2317), .B(n2373), .C(n1297), .Y(n2576) );
  OAI21X1 U2255 ( .A(n2318), .B(n2343), .C(n1299), .Y(n2575) );
  OAI21X1 U2256 ( .A(n2318), .B(n2345), .C(n1301), .Y(n2574) );
  OAI21X1 U2257 ( .A(n2318), .B(n2347), .C(n1303), .Y(n2573) );
  OAI21X1 U2258 ( .A(n2318), .B(n2349), .C(n1305), .Y(n2572) );
  OAI21X1 U2259 ( .A(n2318), .B(n2351), .C(n1307), .Y(n2571) );
  OAI21X1 U2260 ( .A(n2318), .B(n2353), .C(n1309), .Y(n2570) );
  OAI21X1 U2261 ( .A(n2318), .B(n2355), .C(n1311), .Y(n2569) );
  OAI21X1 U2262 ( .A(n2318), .B(n2357), .C(n1313), .Y(n2568) );
  OAI21X1 U2263 ( .A(n2319), .B(n2359), .C(n1315), .Y(n2567) );
  OAI21X1 U2264 ( .A(n2319), .B(n2361), .C(n1317), .Y(n2566) );
  OAI21X1 U2265 ( .A(n2319), .B(n2363), .C(n1319), .Y(n2565) );
  OAI21X1 U2266 ( .A(n2319), .B(n2365), .C(n1321), .Y(n2564) );
  OAI21X1 U2267 ( .A(n2319), .B(n2367), .C(n1323), .Y(n2563) );
  OAI21X1 U2268 ( .A(n2319), .B(n2369), .C(n1325), .Y(n2562) );
  OAI21X1 U2269 ( .A(n2319), .B(n2371), .C(n1327), .Y(n2561) );
  OAI21X1 U2270 ( .A(n2319), .B(n2373), .C(n1329), .Y(n2560) );
  OAI21X1 U2271 ( .A(n2320), .B(n2343), .C(n1331), .Y(n2559) );
  OAI21X1 U2272 ( .A(n2320), .B(n2345), .C(n1333), .Y(n2558) );
  OAI21X1 U2273 ( .A(n2320), .B(n2347), .C(n1335), .Y(n2557) );
  OAI21X1 U2274 ( .A(n2320), .B(n2349), .C(n1337), .Y(n2556) );
  OAI21X1 U2275 ( .A(n2320), .B(n2351), .C(n1339), .Y(n2555) );
  OAI21X1 U2276 ( .A(n2320), .B(n2353), .C(n1341), .Y(n2554) );
  OAI21X1 U2277 ( .A(n2320), .B(n2355), .C(n1343), .Y(n2553) );
  OAI21X1 U2278 ( .A(n2320), .B(n2357), .C(n1345), .Y(n2552) );
  OAI21X1 U2279 ( .A(n2321), .B(n2359), .C(n1347), .Y(n2551) );
  OAI21X1 U2280 ( .A(n2321), .B(n2361), .C(n1349), .Y(n2550) );
  OAI21X1 U2281 ( .A(n2321), .B(n2363), .C(n1351), .Y(n2549) );
  OAI21X1 U2282 ( .A(n2321), .B(n2365), .C(n1353), .Y(n2548) );
  OAI21X1 U2283 ( .A(n2321), .B(n2367), .C(n1355), .Y(n2547) );
  OAI21X1 U2284 ( .A(n2321), .B(n2369), .C(n1357), .Y(n2546) );
  OAI21X1 U2285 ( .A(n2321), .B(n2371), .C(n1359), .Y(n2545) );
  OAI21X1 U2286 ( .A(n2321), .B(n2373), .C(n1361), .Y(n2544) );
  OAI21X1 U2287 ( .A(n2322), .B(n2343), .C(n1363), .Y(n2543) );
  OAI21X1 U2288 ( .A(n2322), .B(n2345), .C(n1365), .Y(n2542) );
  OAI21X1 U2289 ( .A(n2322), .B(n2347), .C(n1367), .Y(n2541) );
  OAI21X1 U2290 ( .A(n2322), .B(n2349), .C(n1369), .Y(n2540) );
  OAI21X1 U2291 ( .A(n2322), .B(n2351), .C(n1371), .Y(n2539) );
  OAI21X1 U2292 ( .A(n2322), .B(n2353), .C(n1373), .Y(n2538) );
  OAI21X1 U2293 ( .A(n2322), .B(n2355), .C(n1375), .Y(n2537) );
  OAI21X1 U2294 ( .A(n2322), .B(n2357), .C(n1377), .Y(n2536) );
  OAI21X1 U2295 ( .A(n2322), .B(n2360), .C(n1379), .Y(n2535) );
  OAI21X1 U2296 ( .A(n2322), .B(n2362), .C(n1381), .Y(n2534) );
  OAI21X1 U2297 ( .A(n2322), .B(n2364), .C(n1383), .Y(n2533) );
  OAI21X1 U2298 ( .A(n2322), .B(n2366), .C(n1385), .Y(n2532) );
  OAI21X1 U2299 ( .A(n2322), .B(n2368), .C(n1387), .Y(n2531) );
  OAI21X1 U2300 ( .A(n2322), .B(n2370), .C(n1389), .Y(n2530) );
  OAI21X1 U2301 ( .A(n2322), .B(n2372), .C(n1391), .Y(n2529) );
  OAI21X1 U2302 ( .A(n2322), .B(n2374), .C(n1393), .Y(n2528) );
  NAND3X1 U2303 ( .A(n2382), .B(n2912), .C(n2384), .Y(n2392) );
  OAI21X1 U2304 ( .A(n2323), .B(n2344), .C(n1395), .Y(n2527) );
  OAI21X1 U2305 ( .A(n2323), .B(n2345), .C(n1397), .Y(n2526) );
  OAI21X1 U2306 ( .A(n2323), .B(n2347), .C(n1399), .Y(n2525) );
  OAI21X1 U2307 ( .A(n2323), .B(n2349), .C(n1401), .Y(n2524) );
  OAI21X1 U2308 ( .A(n2323), .B(n2351), .C(n1403), .Y(n2523) );
  OAI21X1 U2309 ( .A(n2323), .B(n2353), .C(n1405), .Y(n2522) );
  OAI21X1 U2310 ( .A(n2323), .B(n2355), .C(n1407), .Y(n2521) );
  OAI21X1 U2311 ( .A(n2323), .B(n2357), .C(n1409), .Y(n2520) );
  OAI21X1 U2312 ( .A(n2324), .B(n2359), .C(n1411), .Y(n2519) );
  OAI21X1 U2313 ( .A(n2324), .B(n2361), .C(n1413), .Y(n2518) );
  OAI21X1 U2314 ( .A(n2324), .B(n2363), .C(n1415), .Y(n2517) );
  OAI21X1 U2315 ( .A(n2324), .B(n2365), .C(n1417), .Y(n2516) );
  OAI21X1 U2316 ( .A(n2324), .B(n2367), .C(n1419), .Y(n2515) );
  OAI21X1 U2317 ( .A(n2324), .B(n2369), .C(n1421), .Y(n2514) );
  OAI21X1 U2318 ( .A(n2324), .B(n2371), .C(n1423), .Y(n2513) );
  OAI21X1 U2319 ( .A(n2324), .B(n2373), .C(n1425), .Y(n2512) );
  OAI21X1 U2320 ( .A(n2325), .B(n2344), .C(n1427), .Y(n2511) );
  OAI21X1 U2321 ( .A(n2325), .B(n2345), .C(n1429), .Y(n2510) );
  OAI21X1 U2322 ( .A(n2325), .B(n2347), .C(n1431), .Y(n2509) );
  OAI21X1 U2323 ( .A(n2325), .B(n2349), .C(n1433), .Y(n2508) );
  OAI21X1 U2324 ( .A(n2325), .B(n2351), .C(n1435), .Y(n2507) );
  OAI21X1 U2325 ( .A(n2325), .B(n2353), .C(n1437), .Y(n2506) );
  OAI21X1 U2326 ( .A(n2325), .B(n2355), .C(n1439), .Y(n2505) );
  OAI21X1 U2327 ( .A(n2325), .B(n2357), .C(n1441), .Y(n2504) );
  OAI21X1 U2328 ( .A(n2326), .B(n2359), .C(n1443), .Y(n2503) );
  OAI21X1 U2329 ( .A(n2326), .B(n2361), .C(n1445), .Y(n2502) );
  OAI21X1 U2330 ( .A(n2326), .B(n2363), .C(n1447), .Y(n2501) );
  OAI21X1 U2331 ( .A(n2326), .B(n2365), .C(n1449), .Y(n2500) );
  OAI21X1 U2332 ( .A(n2326), .B(n2367), .C(n1451), .Y(n2499) );
  OAI21X1 U2333 ( .A(n2326), .B(n2369), .C(n1453), .Y(n2498) );
  OAI21X1 U2334 ( .A(n2326), .B(n2371), .C(n1455), .Y(n2497) );
  OAI21X1 U2335 ( .A(n2326), .B(n2373), .C(n1457), .Y(n2496) );
  OAI21X1 U2336 ( .A(n2327), .B(n2344), .C(n1459), .Y(n2495) );
  OAI21X1 U2337 ( .A(n2327), .B(n2346), .C(n1461), .Y(n2494) );
  OAI21X1 U2338 ( .A(n2327), .B(n2348), .C(n1463), .Y(n2493) );
  OAI21X1 U2339 ( .A(n2327), .B(n2350), .C(n1465), .Y(n2492) );
  OAI21X1 U2340 ( .A(n2327), .B(n2352), .C(n1467), .Y(n2491) );
  OAI21X1 U2341 ( .A(n2327), .B(n2354), .C(n1469), .Y(n2490) );
  OAI21X1 U2342 ( .A(n2327), .B(n2356), .C(n1471), .Y(n2489) );
  OAI21X1 U2343 ( .A(n2327), .B(n2358), .C(n1473), .Y(n2488) );
  OAI21X1 U2344 ( .A(n2328), .B(n2359), .C(n1475), .Y(n2487) );
  OAI21X1 U2345 ( .A(n2328), .B(n2361), .C(n1477), .Y(n2486) );
  OAI21X1 U2346 ( .A(n2328), .B(n2363), .C(n1479), .Y(n2485) );
  OAI21X1 U2347 ( .A(n2328), .B(n2365), .C(n1481), .Y(n2484) );
  OAI21X1 U2348 ( .A(n2328), .B(n2367), .C(n1483), .Y(n2483) );
  OAI21X1 U2349 ( .A(n2328), .B(n2369), .C(n1485), .Y(n2482) );
  OAI21X1 U2350 ( .A(n2328), .B(n2371), .C(n1487), .Y(n2481) );
  OAI21X1 U2351 ( .A(n2328), .B(n2373), .C(n1489), .Y(n2480) );
  OAI21X1 U2352 ( .A(n2329), .B(n2344), .C(n1491), .Y(n2479) );
  OAI21X1 U2353 ( .A(n2329), .B(n2345), .C(n1493), .Y(n2478) );
  OAI21X1 U2354 ( .A(n2329), .B(n2347), .C(n1495), .Y(n2477) );
  OAI21X1 U2355 ( .A(n2329), .B(n2349), .C(n1497), .Y(n2476) );
  OAI21X1 U2356 ( .A(n2329), .B(n2351), .C(n1499), .Y(n2475) );
  OAI21X1 U2357 ( .A(n2329), .B(n2353), .C(n1501), .Y(n2474) );
  OAI21X1 U2358 ( .A(n2329), .B(n2355), .C(n1503), .Y(n2473) );
  OAI21X1 U2359 ( .A(n2329), .B(n2357), .C(n1505), .Y(n2472) );
  OAI21X1 U2360 ( .A(n2330), .B(n2359), .C(n1507), .Y(n2471) );
  OAI21X1 U2361 ( .A(n2330), .B(n2361), .C(n1509), .Y(n2470) );
  OAI21X1 U2362 ( .A(n2330), .B(n2363), .C(n1511), .Y(n2469) );
  OAI21X1 U2363 ( .A(n2330), .B(n2365), .C(n1513), .Y(n2468) );
  OAI21X1 U2364 ( .A(n2330), .B(n2367), .C(n1515), .Y(n2467) );
  OAI21X1 U2365 ( .A(n2330), .B(n2369), .C(n1517), .Y(n2466) );
  OAI21X1 U2366 ( .A(n2330), .B(n2371), .C(n1519), .Y(n2465) );
  OAI21X1 U2367 ( .A(n2330), .B(n2373), .C(n1521), .Y(n2464) );
  OAI21X1 U2368 ( .A(n2331), .B(n2344), .C(n1523), .Y(n2463) );
  OAI21X1 U2369 ( .A(n2331), .B(n2345), .C(n1525), .Y(n2462) );
  OAI21X1 U2370 ( .A(n2331), .B(n2347), .C(n1527), .Y(n2461) );
  OAI21X1 U2371 ( .A(n2331), .B(n2349), .C(n1529), .Y(n2460) );
  OAI21X1 U2372 ( .A(n2331), .B(n2351), .C(n1531), .Y(n2459) );
  OAI21X1 U2373 ( .A(n2331), .B(n2353), .C(n1533), .Y(n2458) );
  OAI21X1 U2374 ( .A(n2331), .B(n2355), .C(n1535), .Y(n2457) );
  OAI21X1 U2375 ( .A(n2331), .B(n2357), .C(n1537), .Y(n2456) );
  OAI21X1 U2376 ( .A(n2332), .B(n2360), .C(n1539), .Y(n2455) );
  OAI21X1 U2377 ( .A(n2332), .B(n2362), .C(n1541), .Y(n2454) );
  OAI21X1 U2378 ( .A(n2332), .B(n2364), .C(n1543), .Y(n2453) );
  OAI21X1 U2379 ( .A(n2332), .B(n2366), .C(n1545), .Y(n2452) );
  OAI21X1 U2380 ( .A(n2332), .B(n2368), .C(n1547), .Y(n2451) );
  OAI21X1 U2381 ( .A(n2332), .B(n2370), .C(n1549), .Y(n2450) );
  OAI21X1 U2382 ( .A(n2332), .B(n2372), .C(n1551), .Y(n2449) );
  OAI21X1 U2383 ( .A(n2332), .B(n2374), .C(n1553), .Y(n2448) );
  OAI21X1 U2384 ( .A(n2333), .B(n2344), .C(n1555), .Y(n2447) );
  OAI21X1 U2385 ( .A(n2333), .B(n2346), .C(n1557), .Y(n2446) );
  OAI21X1 U2386 ( .A(n2333), .B(n2348), .C(n1559), .Y(n2445) );
  OAI21X1 U2387 ( .A(n2333), .B(n2350), .C(n1561), .Y(n2444) );
  OAI21X1 U2388 ( .A(n2333), .B(n2352), .C(n1563), .Y(n2443) );
  OAI21X1 U2389 ( .A(n2333), .B(n2354), .C(n1565), .Y(n2442) );
  OAI21X1 U2390 ( .A(n2333), .B(n2356), .C(n1567), .Y(n2441) );
  OAI21X1 U2391 ( .A(n2333), .B(n2358), .C(n1569), .Y(n2440) );
  OAI21X1 U2392 ( .A(n2334), .B(n2359), .C(n1571), .Y(n2439) );
  OAI21X1 U2393 ( .A(n2334), .B(n2361), .C(n1573), .Y(n2438) );
  OAI21X1 U2394 ( .A(n2334), .B(n2363), .C(n1575), .Y(n2437) );
  OAI21X1 U2395 ( .A(n2334), .B(n2365), .C(n1577), .Y(n2436) );
  OAI21X1 U2396 ( .A(n2334), .B(n2367), .C(n1579), .Y(n2435) );
  OAI21X1 U2397 ( .A(n2334), .B(n2369), .C(n1581), .Y(n2434) );
  OAI21X1 U2398 ( .A(n2334), .B(n2371), .C(n1583), .Y(n2433) );
  OAI21X1 U2399 ( .A(n2334), .B(n2373), .C(n1585), .Y(n2432) );
  OAI21X1 U2400 ( .A(n2335), .B(n2344), .C(n1587), .Y(n2431) );
  OAI21X1 U2401 ( .A(n2335), .B(n2345), .C(n1589), .Y(n2430) );
  OAI21X1 U2402 ( .A(n2335), .B(n2347), .C(n1591), .Y(n2429) );
  OAI21X1 U2403 ( .A(n2335), .B(n2349), .C(n1593), .Y(n2428) );
  OAI21X1 U2404 ( .A(n2335), .B(n2351), .C(n1595), .Y(n2427) );
  OAI21X1 U2405 ( .A(n2335), .B(n2353), .C(n1597), .Y(n2426) );
  OAI21X1 U2406 ( .A(n2335), .B(n2355), .C(n1599), .Y(n2425) );
  OAI21X1 U2407 ( .A(n2335), .B(n2357), .C(n1601), .Y(n2424) );
  OAI21X1 U2408 ( .A(n2336), .B(n2359), .C(n1603), .Y(n2423) );
  OAI21X1 U2409 ( .A(n2336), .B(n2361), .C(n1605), .Y(n2422) );
  OAI21X1 U2410 ( .A(n2336), .B(n2363), .C(n1607), .Y(n2421) );
  OAI21X1 U2411 ( .A(n2336), .B(n2365), .C(n1609), .Y(n2420) );
  OAI21X1 U2412 ( .A(n2336), .B(n2367), .C(n1611), .Y(n2419) );
  OAI21X1 U2413 ( .A(n2336), .B(n2369), .C(n1613), .Y(n2418) );
  OAI21X1 U2414 ( .A(n2336), .B(n2371), .C(n1615), .Y(n2417) );
  OAI21X1 U2415 ( .A(n2336), .B(n2373), .C(n1617), .Y(n2416) );
  OAI21X1 U2416 ( .A(n2337), .B(n2344), .C(n1619), .Y(n2415) );
  OAI21X1 U2417 ( .A(n2337), .B(n2345), .C(n1621), .Y(n2414) );
  OAI21X1 U2418 ( .A(n2337), .B(n2347), .C(n1623), .Y(n2413) );
  OAI21X1 U2419 ( .A(n2337), .B(n2349), .C(n1625), .Y(n2412) );
  OAI21X1 U2420 ( .A(n2337), .B(n2351), .C(n1627), .Y(n2411) );
  OAI21X1 U2421 ( .A(n2337), .B(n2353), .C(n1629), .Y(n2410) );
  OAI21X1 U2422 ( .A(n2337), .B(n2355), .C(n1631), .Y(n2409) );
  OAI21X1 U2423 ( .A(n2337), .B(n2357), .C(n1633), .Y(n2408) );
  OAI21X1 U2424 ( .A(n2337), .B(n2359), .C(n1635), .Y(n2407) );
  OAI21X1 U2425 ( .A(n2337), .B(n2361), .C(n1637), .Y(n2406) );
  OAI21X1 U2426 ( .A(n2337), .B(n2363), .C(n1639), .Y(n2405) );
  OAI21X1 U2427 ( .A(n2337), .B(n2365), .C(n1641), .Y(n2404) );
  OAI21X1 U2428 ( .A(n2337), .B(n2367), .C(n1643), .Y(n2403) );
  OAI21X1 U2429 ( .A(n2337), .B(n2369), .C(n1645), .Y(n2402) );
  OAI21X1 U2430 ( .A(n2337), .B(n2371), .C(n1647), .Y(n2401) );
  OAI21X1 U2431 ( .A(n2337), .B(n2373), .C(n1649), .Y(n2400) );
endmodule


module memc_Size16_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2189), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2190), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2191), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2192), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2193), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2194), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2195), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2196), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2197), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2198), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2199), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2200), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2201), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2202), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2203), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2204), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2205), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2206), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2207), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2208), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2209), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2210), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2211), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2212), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2213), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2214), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2215), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2216), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2217), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2218), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2219), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2220), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2221), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2222), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2223), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2224), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2225), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2226), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2227), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2228), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2229), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2230), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2231), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2232), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2233), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2234), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2235), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2236), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2237), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2238), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2239), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2240), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2241), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2242), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2243), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2244), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2245), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2246), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2247), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2248), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2249), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2250), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2251), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2252), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2253), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2254), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2255), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2256), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2257), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2258), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2259), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2260), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2261), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2262), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2263), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2264), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2265), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2266), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2267), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2268), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2269), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2270), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2271), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2272), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2273), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2274), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2275), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2276), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2277), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2278), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2279), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2280), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2281), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2282), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2283), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2284), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2285), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2286), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2287), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2288), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2289), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2290), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2291), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2292), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2293), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2294), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2295), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2296), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2297), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2298), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2299), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2300), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2301), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2302), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2303), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2304), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2305), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2306), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2307), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2308), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2309), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2310), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2311), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2312), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2313), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2314), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2315), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2316), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2317), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2318), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2319), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2320), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2321), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2322), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2323), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2324), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2325), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2326), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2327), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2328), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2329), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2330), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2331), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2332), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2333), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2334), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2335), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2336), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2337), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2338), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2339), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2340), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2341), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2342), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2343), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2344), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2345), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2346), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2347), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2348), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2349), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2350), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2351), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2352), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2353), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2354), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2355), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2356), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2357), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2358), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2359), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2360), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2361), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2362), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2363), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2364), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2365), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2366), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2367), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2368), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2369), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2370), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2371), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2372), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2373), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2374), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2375), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2376), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2377), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2378), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2379), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2380), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2381), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2382), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2383), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2384), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2385), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2386), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2387), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2388), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2389), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2390), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2391), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2392), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2393), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2394), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2395), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2396), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2397), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2398), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2399), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2400), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2401), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2402), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2403), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2404), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2405), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2406), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2407), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2408), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2409), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2410), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2411), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2412), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2413), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2414), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2415), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2416), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2417), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2418), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2419), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2420), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2421), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2422), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2423), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2424), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2425), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2426), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2427), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2428), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2429), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2430), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2431), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2432), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2433), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2434), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2435), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2436), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2437), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2438), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2439), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2440), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2441), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2442), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2443), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2444), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2445), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2446), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2447), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2448), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2449), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2450), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2451), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2452), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2453), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2454), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2455), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2456), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2457), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2458), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2459), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2460), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2461), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2462), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2463), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2464), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2465), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2466), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2467), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2468), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2469), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2470), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2471), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2472), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2473), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2474), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2475), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2476), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2477), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2478), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2479), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2480), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2481), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2482), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2483), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2484), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2485), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2486), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2487), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2488), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2489), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2490), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2491), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2492), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2493), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2494), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2495), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2496), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2497), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2498), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2499), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2500), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2501), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2502), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2503), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2504), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2505), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2506), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2507), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2508), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2509), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2510), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2511), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2512), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2513), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2514), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2515), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2516), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2517), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2518), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2519), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2520), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2521), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2522), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2523), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2524), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2525), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2526), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2527), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2528), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2529), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2530), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2531), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2532), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2533), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2534), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2535), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2536), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2537), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2538), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2539), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2540), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2541), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2542), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2543), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2544), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2545), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2546), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2547), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2548), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2549), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2550), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2551), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2552), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2553), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2554), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2555), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2556), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2557), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2558), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2559), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2560), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2561), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2562), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2563), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2564), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2565), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2566), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2567), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2568), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2569), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2570), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2571), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2572), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2573), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2574), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2575), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2576), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2577), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2578), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2579), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2580), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2581), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2582), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2583), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2584), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2585), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2586), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2587), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2588), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2589), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2590), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2591), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2592), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2593), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2594), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2595), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2596), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2597), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2598), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2599), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2600), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2601), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2602), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2603), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2604), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2605), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2606), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2607), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2608), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2609), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2610), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2611), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2612), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2613), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2614), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2615), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2616), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2617), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2618), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2619), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2620), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2621), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2622), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2623), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2624), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2625), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2626), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2627), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2628), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2629), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2630), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2631), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2632), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2633), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2634), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2635), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2636), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2637), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2638), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2639), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2640), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2641), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2642), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2643), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2644), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2645), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2646), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2647), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2648), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2649), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2650), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2651), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2652), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2653), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2654), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2655), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2656), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2657), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2658), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2659), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2660), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2661), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2662), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2663), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2664), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2665), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2666), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2667), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2668), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2669), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2670), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2671), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2672), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2673), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2674), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2675), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2676), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2677), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2678), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2679), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2680), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2681), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2682), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2683), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2684), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2685), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2686), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2687), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2688), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2689), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2690), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2691), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2692), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2693), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2694), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2695), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2696), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2697), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2698), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2699), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2700), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2701) );
  INVX4 U2 ( .A(n1210), .Y(n1211) );
  INVX4 U3 ( .A(n618), .Y(n619) );
  INVX4 U4 ( .A(n1184), .Y(n1185) );
  INVX4 U5 ( .A(n1182), .Y(n1183) );
  INVX4 U6 ( .A(n620), .Y(n621) );
  INVX4 U7 ( .A(n616), .Y(n617) );
  INVX4 U8 ( .A(n641), .Y(n642) );
  INVX4 U9 ( .A(n639), .Y(n640) );
  INVX4 U10 ( .A(n614), .Y(n615) );
  INVX2 U11 ( .A(n1230), .Y(n1231) );
  INVX1 U12 ( .A(n1965), .Y(n1810) );
  INVX1 U13 ( .A(n1965), .Y(n1809) );
  INVX2 U14 ( .A(n1812), .Y(n1813) );
  INVX1 U15 ( .A(n1965), .Y(n1811) );
  INVX1 U16 ( .A(n1801), .Y(N23) );
  INVX1 U17 ( .A(n1804), .Y(N20) );
  INVX1 U18 ( .A(n1960), .Y(n1819) );
  INVX2 U19 ( .A(n1820), .Y(n1821) );
  INVX2 U20 ( .A(n1819), .Y(n1824) );
  INVX2 U21 ( .A(n1819), .Y(n1825) );
  INVX2 U22 ( .A(n1819), .Y(n1826) );
  INVX2 U23 ( .A(n1819), .Y(n1829) );
  INVX1 U24 ( .A(n1792), .Y(N32) );
  INVX1 U25 ( .A(n1793), .Y(N31) );
  INVX1 U26 ( .A(n1794), .Y(N30) );
  INVX1 U27 ( .A(n1795), .Y(N29) );
  INVX1 U28 ( .A(n1796), .Y(N28) );
  INVX1 U29 ( .A(n1797), .Y(N27) );
  INVX1 U30 ( .A(n1799), .Y(N25) );
  INVX1 U31 ( .A(n1802), .Y(N22) );
  INVX1 U32 ( .A(n1803), .Y(N21) );
  INVX1 U33 ( .A(n1805), .Y(N19) );
  INVX1 U34 ( .A(n1806), .Y(N18) );
  INVX1 U35 ( .A(n1807), .Y(N17) );
  INVX1 U36 ( .A(n1798), .Y(N26) );
  INVX1 U37 ( .A(n1800), .Y(N24) );
  BUFX2 U38 ( .A(n1255), .Y(n1862) );
  BUFX2 U39 ( .A(n1257), .Y(n1864) );
  BUFX2 U40 ( .A(n1259), .Y(n1866) );
  BUFX2 U41 ( .A(n1261), .Y(n1868) );
  BUFX2 U42 ( .A(n1263), .Y(n1870) );
  BUFX2 U43 ( .A(n1265), .Y(n1872) );
  BUFX2 U44 ( .A(n1267), .Y(n1874) );
  BUFX2 U45 ( .A(n1269), .Y(n1876) );
  BUFX2 U46 ( .A(n1271), .Y(n1878) );
  BUFX2 U47 ( .A(n1273), .Y(n1880) );
  BUFX2 U48 ( .A(n1275), .Y(n1882) );
  BUFX2 U49 ( .A(n1277), .Y(n1884) );
  BUFX2 U50 ( .A(n1279), .Y(n1886) );
  BUFX2 U51 ( .A(n1281), .Y(n1888) );
  BUFX2 U52 ( .A(n1283), .Y(n1891) );
  BUFX2 U53 ( .A(n1285), .Y(n1893) );
  BUFX2 U54 ( .A(n1287), .Y(n1895) );
  BUFX2 U55 ( .A(n1289), .Y(n1897) );
  BUFX2 U56 ( .A(n1291), .Y(n1899) );
  BUFX2 U57 ( .A(n1293), .Y(n1901) );
  BUFX2 U58 ( .A(n1295), .Y(n1903) );
  BUFX2 U59 ( .A(n1297), .Y(n1906) );
  BUFX2 U60 ( .A(n1299), .Y(n1908) );
  BUFX2 U61 ( .A(n1301), .Y(n1910) );
  BUFX2 U62 ( .A(n1303), .Y(n1912) );
  BUFX2 U63 ( .A(n1305), .Y(n1914) );
  BUFX2 U64 ( .A(n1307), .Y(n1916) );
  BUFX2 U65 ( .A(n1309), .Y(n1918) );
  INVX2 U66 ( .A(n1860), .Y(n1832) );
  INVX2 U67 ( .A(n1960), .Y(n1820) );
  INVX1 U68 ( .A(n1962), .Y(n1812) );
  INVX1 U69 ( .A(n1958), .Y(n1859) );
  INVX1 U70 ( .A(n1967), .Y(n1966) );
  INVX1 U71 ( .A(N14), .Y(n1967) );
  INVX1 U72 ( .A(n1859), .Y(n1860) );
  BUFX2 U73 ( .A(n1255), .Y(n1863) );
  BUFX2 U74 ( .A(n1269), .Y(n1877) );
  BUFX2 U75 ( .A(n1271), .Y(n1879) );
  BUFX2 U76 ( .A(n1273), .Y(n1881) );
  BUFX2 U77 ( .A(n1261), .Y(n1869) );
  BUFX2 U78 ( .A(n1263), .Y(n1871) );
  BUFX2 U79 ( .A(n1267), .Y(n1875) );
  BUFX2 U80 ( .A(n1257), .Y(n1865) );
  INVX1 U81 ( .A(n1965), .Y(n1964) );
  INVX1 U82 ( .A(N13), .Y(n1965) );
  BUFX2 U83 ( .A(n1275), .Y(n1883) );
  BUFX2 U84 ( .A(n1279), .Y(n1887) );
  BUFX2 U85 ( .A(n1281), .Y(n1889) );
  BUFX2 U86 ( .A(n1259), .Y(n1867) );
  BUFX2 U87 ( .A(n1265), .Y(n1873) );
  BUFX2 U88 ( .A(n1283), .Y(n1892) );
  BUFX2 U89 ( .A(n1285), .Y(n1894) );
  BUFX2 U90 ( .A(n1287), .Y(n1896) );
  BUFX2 U91 ( .A(n1289), .Y(n1898) );
  BUFX2 U92 ( .A(n1291), .Y(n1900) );
  BUFX2 U93 ( .A(n1293), .Y(n1902) );
  BUFX2 U94 ( .A(n1295), .Y(n1904) );
  INVX1 U95 ( .A(n1967), .Y(n1808) );
  INVX1 U96 ( .A(n1252), .Y(n1905) );
  INVX1 U97 ( .A(n1253), .Y(n1920) );
  BUFX2 U98 ( .A(n1277), .Y(n1885) );
  BUFX2 U99 ( .A(n1297), .Y(n1907) );
  BUFX2 U100 ( .A(n1301), .Y(n1911) );
  BUFX2 U101 ( .A(n1303), .Y(n1913) );
  BUFX2 U102 ( .A(n1305), .Y(n1915) );
  BUFX2 U103 ( .A(n1307), .Y(n1917) );
  BUFX2 U104 ( .A(n1309), .Y(n1919) );
  BUFX2 U105 ( .A(n1299), .Y(n1909) );
  INVX1 U106 ( .A(n1251), .Y(n1890) );
  INVX4 U107 ( .A(n622), .Y(n1924) );
  INVX1 U108 ( .A(rst), .Y(n1957) );
  AND2X2 U109 ( .A(\mem<31><0> ), .B(n640), .Y(n1) );
  INVX1 U110 ( .A(n1), .Y(n2) );
  AND2X2 U111 ( .A(\mem<31><15> ), .B(n640), .Y(n3) );
  INVX1 U112 ( .A(n3), .Y(n4) );
  AND2X2 U113 ( .A(\mem<30><0> ), .B(n642), .Y(n5) );
  INVX1 U114 ( .A(n5), .Y(n6) );
  AND2X2 U115 ( .A(\mem<30><15> ), .B(n642), .Y(n7) );
  INVX1 U116 ( .A(n7), .Y(n8) );
  AND2X2 U117 ( .A(\mem<29><15> ), .B(n644), .Y(n9) );
  INVX1 U118 ( .A(n9), .Y(n10) );
  AND2X2 U119 ( .A(\mem<28><0> ), .B(n648), .Y(n11) );
  INVX1 U120 ( .A(n11), .Y(n12) );
  AND2X2 U121 ( .A(\mem<28><15> ), .B(n647), .Y(n13) );
  INVX1 U122 ( .A(n13), .Y(n14) );
  AND2X2 U123 ( .A(\mem<27><0> ), .B(n1163), .Y(n15) );
  INVX1 U124 ( .A(n15), .Y(n16) );
  AND2X2 U125 ( .A(\mem<27><15> ), .B(n650), .Y(n17) );
  INVX1 U126 ( .A(n17), .Y(n18) );
  AND2X2 U127 ( .A(\mem<26><15> ), .B(n1165), .Y(n19) );
  INVX1 U128 ( .A(n19), .Y(n20) );
  AND2X2 U129 ( .A(\mem<25><0> ), .B(n1169), .Y(n21) );
  INVX1 U130 ( .A(n21), .Y(n22) );
  AND2X2 U131 ( .A(\mem<25><15> ), .B(n1168), .Y(n23) );
  INVX1 U132 ( .A(n23), .Y(n24) );
  AND2X2 U133 ( .A(\mem<24><0> ), .B(n1172), .Y(n25) );
  INVX1 U134 ( .A(n25), .Y(n26) );
  AND2X2 U135 ( .A(\mem<24><15> ), .B(n1171), .Y(n27) );
  INVX1 U136 ( .A(n27), .Y(n28) );
  AND2X2 U137 ( .A(\mem<23><0> ), .B(n1175), .Y(n29) );
  INVX1 U138 ( .A(n29), .Y(n30) );
  AND2X2 U139 ( .A(\mem<23><1> ), .B(n1175), .Y(n31) );
  INVX1 U140 ( .A(n31), .Y(n32) );
  AND2X2 U141 ( .A(\mem<23><2> ), .B(n1175), .Y(n33) );
  INVX1 U142 ( .A(n33), .Y(n34) );
  AND2X2 U143 ( .A(\mem<23><3> ), .B(n1175), .Y(n35) );
  INVX1 U144 ( .A(n35), .Y(n36) );
  AND2X2 U145 ( .A(\mem<23><4> ), .B(n1175), .Y(n37) );
  INVX1 U146 ( .A(n37), .Y(n38) );
  AND2X2 U147 ( .A(\mem<23><5> ), .B(n1175), .Y(n39) );
  INVX1 U148 ( .A(n39), .Y(n40) );
  AND2X2 U149 ( .A(\mem<23><6> ), .B(n1175), .Y(n41) );
  INVX1 U150 ( .A(n41), .Y(n42) );
  AND2X2 U151 ( .A(\mem<23><7> ), .B(n1175), .Y(n43) );
  INVX1 U152 ( .A(n43), .Y(n44) );
  AND2X2 U153 ( .A(\mem<23><8> ), .B(n1174), .Y(n45) );
  INVX1 U154 ( .A(n45), .Y(n46) );
  AND2X2 U155 ( .A(\mem<23><9> ), .B(n1174), .Y(n47) );
  INVX1 U156 ( .A(n47), .Y(n48) );
  AND2X2 U157 ( .A(\mem<23><10> ), .B(n1174), .Y(n49) );
  INVX1 U158 ( .A(n49), .Y(n50) );
  AND2X2 U159 ( .A(\mem<23><11> ), .B(n1174), .Y(n51) );
  INVX1 U160 ( .A(n51), .Y(n52) );
  AND2X2 U161 ( .A(\mem<23><12> ), .B(n1174), .Y(n53) );
  INVX1 U162 ( .A(n53), .Y(n54) );
  AND2X2 U163 ( .A(\mem<23><13> ), .B(n1174), .Y(n55) );
  INVX1 U164 ( .A(n55), .Y(n56) );
  AND2X2 U165 ( .A(\mem<23><14> ), .B(n1174), .Y(n57) );
  INVX1 U166 ( .A(n57), .Y(n58) );
  AND2X2 U167 ( .A(\mem<23><15> ), .B(n1174), .Y(n59) );
  INVX1 U168 ( .A(n59), .Y(n60) );
  AND2X2 U169 ( .A(\mem<22><0> ), .B(n1178), .Y(n61) );
  INVX1 U170 ( .A(n61), .Y(n62) );
  AND2X2 U171 ( .A(\mem<22><1> ), .B(n1178), .Y(n63) );
  INVX1 U172 ( .A(n63), .Y(n64) );
  AND2X2 U173 ( .A(\mem<22><2> ), .B(n1178), .Y(n65) );
  INVX1 U174 ( .A(n65), .Y(n66) );
  AND2X2 U175 ( .A(\mem<22><3> ), .B(n1178), .Y(n67) );
  INVX1 U176 ( .A(n67), .Y(n68) );
  AND2X2 U177 ( .A(\mem<22><4> ), .B(n1178), .Y(n69) );
  INVX1 U178 ( .A(n69), .Y(n70) );
  AND2X2 U179 ( .A(\mem<22><5> ), .B(n1178), .Y(n71) );
  INVX1 U180 ( .A(n71), .Y(n72) );
  AND2X2 U181 ( .A(\mem<22><6> ), .B(n1178), .Y(n73) );
  INVX1 U182 ( .A(n73), .Y(n74) );
  AND2X2 U183 ( .A(\mem<22><7> ), .B(n1178), .Y(n75) );
  INVX1 U184 ( .A(n75), .Y(n76) );
  AND2X2 U185 ( .A(\mem<22><8> ), .B(n1177), .Y(n77) );
  INVX1 U186 ( .A(n77), .Y(n78) );
  AND2X2 U187 ( .A(\mem<22><9> ), .B(n1177), .Y(n79) );
  INVX1 U188 ( .A(n79), .Y(n80) );
  AND2X2 U189 ( .A(\mem<22><10> ), .B(n1177), .Y(n81) );
  INVX1 U190 ( .A(n81), .Y(n82) );
  AND2X2 U191 ( .A(\mem<22><11> ), .B(n1177), .Y(n83) );
  INVX1 U192 ( .A(n83), .Y(n84) );
  AND2X2 U193 ( .A(\mem<22><12> ), .B(n1177), .Y(n85) );
  INVX1 U194 ( .A(n85), .Y(n86) );
  AND2X2 U195 ( .A(\mem<22><13> ), .B(n1177), .Y(n87) );
  INVX1 U196 ( .A(n87), .Y(n88) );
  AND2X2 U197 ( .A(\mem<22><14> ), .B(n1177), .Y(n89) );
  INVX1 U198 ( .A(n89), .Y(n90) );
  AND2X2 U199 ( .A(\mem<22><15> ), .B(n1177), .Y(n91) );
  INVX1 U200 ( .A(n91), .Y(n92) );
  AND2X2 U201 ( .A(\mem<21><0> ), .B(n1181), .Y(n93) );
  INVX1 U202 ( .A(n93), .Y(n94) );
  AND2X2 U203 ( .A(\mem<21><1> ), .B(n1181), .Y(n95) );
  INVX1 U204 ( .A(n95), .Y(n96) );
  AND2X2 U205 ( .A(\mem<21><2> ), .B(n1181), .Y(n97) );
  INVX1 U206 ( .A(n97), .Y(n98) );
  AND2X2 U207 ( .A(\mem<21><3> ), .B(n1181), .Y(n99) );
  INVX1 U208 ( .A(n99), .Y(n100) );
  AND2X2 U209 ( .A(\mem<21><4> ), .B(n1181), .Y(n101) );
  INVX1 U210 ( .A(n101), .Y(n102) );
  AND2X2 U211 ( .A(\mem<21><5> ), .B(n1181), .Y(n103) );
  INVX1 U212 ( .A(n103), .Y(n104) );
  AND2X2 U213 ( .A(\mem<21><6> ), .B(n1181), .Y(n105) );
  INVX1 U214 ( .A(n105), .Y(n106) );
  AND2X2 U215 ( .A(\mem<21><7> ), .B(n1181), .Y(n107) );
  INVX1 U216 ( .A(n107), .Y(n108) );
  AND2X2 U217 ( .A(\mem<21><8> ), .B(n1180), .Y(n109) );
  INVX1 U218 ( .A(n109), .Y(n110) );
  AND2X2 U219 ( .A(\mem<21><9> ), .B(n1180), .Y(n111) );
  INVX1 U220 ( .A(n111), .Y(n112) );
  AND2X2 U221 ( .A(\mem<21><10> ), .B(n1180), .Y(n113) );
  INVX1 U222 ( .A(n113), .Y(n114) );
  AND2X2 U223 ( .A(\mem<21><11> ), .B(n1180), .Y(n115) );
  INVX1 U224 ( .A(n115), .Y(n116) );
  AND2X2 U225 ( .A(\mem<21><12> ), .B(n1180), .Y(n117) );
  INVX1 U226 ( .A(n117), .Y(n118) );
  AND2X2 U227 ( .A(\mem<21><13> ), .B(n1180), .Y(n119) );
  INVX1 U228 ( .A(n119), .Y(n120) );
  AND2X2 U229 ( .A(\mem<21><14> ), .B(n1180), .Y(n121) );
  INVX1 U230 ( .A(n121), .Y(n122) );
  AND2X2 U231 ( .A(\mem<21><15> ), .B(n1180), .Y(n123) );
  INVX1 U232 ( .A(n123), .Y(n124) );
  AND2X2 U233 ( .A(\mem<18><0> ), .B(n1183), .Y(n125) );
  INVX1 U234 ( .A(n125), .Y(n126) );
  AND2X2 U235 ( .A(\mem<18><1> ), .B(n1183), .Y(n127) );
  INVX1 U236 ( .A(n127), .Y(n128) );
  AND2X2 U237 ( .A(\mem<18><2> ), .B(n1183), .Y(n129) );
  INVX1 U238 ( .A(n129), .Y(n130) );
  AND2X2 U239 ( .A(\mem<18><3> ), .B(n1183), .Y(n131) );
  INVX1 U240 ( .A(n131), .Y(n132) );
  AND2X2 U241 ( .A(\mem<18><4> ), .B(n1183), .Y(n133) );
  INVX1 U242 ( .A(n133), .Y(n134) );
  AND2X2 U243 ( .A(\mem<18><5> ), .B(n1183), .Y(n135) );
  INVX1 U244 ( .A(n135), .Y(n136) );
  AND2X2 U245 ( .A(\mem<18><6> ), .B(n1183), .Y(n137) );
  INVX1 U246 ( .A(n137), .Y(n138) );
  AND2X2 U247 ( .A(\mem<18><7> ), .B(n1183), .Y(n139) );
  INVX1 U248 ( .A(n139), .Y(n140) );
  AND2X2 U249 ( .A(\mem<18><8> ), .B(n1183), .Y(n141) );
  INVX1 U250 ( .A(n141), .Y(n142) );
  AND2X2 U251 ( .A(\mem<18><9> ), .B(n1183), .Y(n143) );
  INVX1 U252 ( .A(n143), .Y(n144) );
  AND2X2 U253 ( .A(\mem<18><10> ), .B(n1183), .Y(n145) );
  INVX1 U254 ( .A(n145), .Y(n146) );
  AND2X2 U255 ( .A(\mem<18><11> ), .B(n1183), .Y(n147) );
  INVX1 U256 ( .A(n147), .Y(n148) );
  AND2X2 U257 ( .A(\mem<18><12> ), .B(n1183), .Y(n149) );
  INVX1 U258 ( .A(n149), .Y(n150) );
  AND2X2 U259 ( .A(\mem<18><13> ), .B(n1183), .Y(n151) );
  INVX1 U260 ( .A(n151), .Y(n152) );
  AND2X2 U261 ( .A(\mem<18><14> ), .B(n1183), .Y(n153) );
  INVX1 U262 ( .A(n153), .Y(n154) );
  AND2X2 U263 ( .A(\mem<18><15> ), .B(n1183), .Y(n155) );
  INVX1 U264 ( .A(n155), .Y(n156) );
  AND2X2 U265 ( .A(\mem<17><0> ), .B(n1185), .Y(n157) );
  INVX1 U266 ( .A(n157), .Y(n158) );
  AND2X2 U267 ( .A(\mem<17><1> ), .B(n1185), .Y(n159) );
  INVX1 U268 ( .A(n159), .Y(n160) );
  AND2X2 U269 ( .A(\mem<17><2> ), .B(n1185), .Y(n161) );
  INVX1 U270 ( .A(n161), .Y(n162) );
  AND2X2 U271 ( .A(\mem<17><3> ), .B(n1185), .Y(n163) );
  INVX1 U272 ( .A(n163), .Y(n164) );
  AND2X2 U273 ( .A(\mem<17><4> ), .B(n1185), .Y(n165) );
  INVX1 U274 ( .A(n165), .Y(n166) );
  AND2X2 U275 ( .A(\mem<17><5> ), .B(n1185), .Y(n167) );
  INVX1 U276 ( .A(n167), .Y(n168) );
  AND2X2 U277 ( .A(\mem<17><6> ), .B(n1185), .Y(n169) );
  INVX1 U278 ( .A(n169), .Y(n170) );
  AND2X2 U279 ( .A(\mem<17><7> ), .B(n1185), .Y(n171) );
  INVX1 U280 ( .A(n171), .Y(n172) );
  AND2X2 U281 ( .A(\mem<17><8> ), .B(n1185), .Y(n173) );
  INVX1 U282 ( .A(n173), .Y(n174) );
  AND2X2 U283 ( .A(\mem<17><9> ), .B(n1185), .Y(n175) );
  INVX1 U284 ( .A(n175), .Y(n176) );
  AND2X2 U285 ( .A(\mem<17><10> ), .B(n1185), .Y(n177) );
  INVX1 U286 ( .A(n177), .Y(n178) );
  AND2X2 U287 ( .A(\mem<17><11> ), .B(n1185), .Y(n179) );
  INVX1 U288 ( .A(n179), .Y(n180) );
  AND2X2 U289 ( .A(\mem<17><12> ), .B(n1185), .Y(n181) );
  INVX1 U290 ( .A(n181), .Y(n182) );
  AND2X2 U291 ( .A(\mem<17><13> ), .B(n1185), .Y(n183) );
  INVX1 U292 ( .A(n183), .Y(n184) );
  AND2X2 U293 ( .A(\mem<17><14> ), .B(n1185), .Y(n185) );
  INVX1 U294 ( .A(n185), .Y(n186) );
  AND2X2 U295 ( .A(\mem<17><15> ), .B(n1185), .Y(n187) );
  INVX1 U296 ( .A(n187), .Y(n188) );
  AND2X2 U297 ( .A(\mem<16><0> ), .B(n1188), .Y(n189) );
  INVX1 U298 ( .A(n189), .Y(n190) );
  AND2X2 U299 ( .A(\mem<16><1> ), .B(n1188), .Y(n191) );
  INVX1 U300 ( .A(n191), .Y(n192) );
  AND2X2 U301 ( .A(\mem<16><2> ), .B(n1188), .Y(n193) );
  INVX1 U302 ( .A(n193), .Y(n194) );
  AND2X2 U303 ( .A(\mem<16><3> ), .B(n1188), .Y(n195) );
  INVX1 U304 ( .A(n195), .Y(n196) );
  AND2X2 U305 ( .A(\mem<16><4> ), .B(n1188), .Y(n197) );
  INVX1 U306 ( .A(n197), .Y(n198) );
  AND2X2 U307 ( .A(\mem<16><5> ), .B(n1188), .Y(n199) );
  INVX1 U308 ( .A(n199), .Y(n200) );
  AND2X2 U309 ( .A(\mem<16><6> ), .B(n1188), .Y(n201) );
  INVX1 U310 ( .A(n201), .Y(n202) );
  AND2X2 U311 ( .A(\mem<16><7> ), .B(n1188), .Y(n203) );
  INVX1 U312 ( .A(n203), .Y(n204) );
  AND2X2 U313 ( .A(\mem<16><8> ), .B(n1187), .Y(n205) );
  INVX1 U314 ( .A(n205), .Y(n206) );
  AND2X2 U315 ( .A(\mem<16><9> ), .B(n1187), .Y(n207) );
  INVX1 U316 ( .A(n207), .Y(n208) );
  AND2X2 U317 ( .A(\mem<16><10> ), .B(n1187), .Y(n209) );
  INVX1 U318 ( .A(n209), .Y(n210) );
  AND2X2 U319 ( .A(\mem<16><11> ), .B(n1187), .Y(n211) );
  INVX1 U320 ( .A(n211), .Y(n212) );
  AND2X2 U321 ( .A(\mem<16><12> ), .B(n1187), .Y(n213) );
  INVX1 U322 ( .A(n213), .Y(n215) );
  AND2X2 U323 ( .A(\mem<16><13> ), .B(n1187), .Y(n216) );
  INVX1 U324 ( .A(n216), .Y(n217) );
  AND2X2 U325 ( .A(\mem<16><14> ), .B(n1187), .Y(n218) );
  INVX1 U326 ( .A(n218), .Y(n219) );
  AND2X2 U327 ( .A(\mem<16><15> ), .B(n1187), .Y(n220) );
  INVX1 U328 ( .A(n220), .Y(n221) );
  AND2X2 U329 ( .A(\mem<15><0> ), .B(n1191), .Y(n222) );
  INVX1 U330 ( .A(n222), .Y(n223) );
  AND2X2 U331 ( .A(\mem<15><1> ), .B(n1191), .Y(n224) );
  INVX1 U332 ( .A(n224), .Y(n225) );
  AND2X2 U333 ( .A(\mem<15><2> ), .B(n1191), .Y(n226) );
  INVX1 U334 ( .A(n226), .Y(n227) );
  AND2X2 U335 ( .A(\mem<15><3> ), .B(n1191), .Y(n228) );
  INVX1 U336 ( .A(n228), .Y(n229) );
  AND2X2 U337 ( .A(\mem<15><4> ), .B(n1191), .Y(n230) );
  INVX1 U338 ( .A(n230), .Y(n231) );
  AND2X2 U339 ( .A(\mem<15><5> ), .B(n1191), .Y(n232) );
  INVX1 U340 ( .A(n232), .Y(n233) );
  AND2X2 U341 ( .A(\mem<15><6> ), .B(n1191), .Y(n234) );
  INVX1 U342 ( .A(n234), .Y(n235) );
  AND2X2 U343 ( .A(\mem<15><7> ), .B(n1191), .Y(n236) );
  INVX1 U344 ( .A(n236), .Y(n237) );
  AND2X2 U345 ( .A(\mem<15><8> ), .B(n1190), .Y(n238) );
  INVX1 U346 ( .A(n238), .Y(n239) );
  AND2X2 U347 ( .A(\mem<15><9> ), .B(n1190), .Y(n240) );
  INVX1 U348 ( .A(n240), .Y(n241) );
  AND2X2 U349 ( .A(\mem<15><10> ), .B(n1190), .Y(n242) );
  INVX1 U350 ( .A(n242), .Y(n243) );
  AND2X2 U351 ( .A(\mem<15><11> ), .B(n1190), .Y(n244) );
  INVX1 U352 ( .A(n244), .Y(n245) );
  AND2X2 U353 ( .A(\mem<15><12> ), .B(n1190), .Y(n246) );
  INVX1 U354 ( .A(n246), .Y(n247) );
  AND2X2 U355 ( .A(\mem<15><13> ), .B(n1190), .Y(n248) );
  INVX1 U356 ( .A(n248), .Y(n249) );
  AND2X2 U357 ( .A(\mem<15><14> ), .B(n1190), .Y(n250) );
  INVX1 U358 ( .A(n250), .Y(n251) );
  AND2X2 U359 ( .A(\mem<15><15> ), .B(n1190), .Y(n252) );
  INVX1 U360 ( .A(n252), .Y(n253) );
  AND2X2 U361 ( .A(\mem<14><0> ), .B(n1194), .Y(n254) );
  INVX1 U362 ( .A(n254), .Y(n255) );
  AND2X2 U363 ( .A(\mem<14><1> ), .B(n1194), .Y(n256) );
  INVX1 U364 ( .A(n256), .Y(n257) );
  AND2X2 U365 ( .A(\mem<14><2> ), .B(n1194), .Y(n258) );
  INVX1 U366 ( .A(n258), .Y(n259) );
  AND2X2 U367 ( .A(\mem<14><3> ), .B(n1194), .Y(n260) );
  INVX1 U368 ( .A(n260), .Y(n261) );
  AND2X2 U369 ( .A(\mem<14><4> ), .B(n1194), .Y(n262) );
  INVX1 U370 ( .A(n262), .Y(n263) );
  AND2X2 U371 ( .A(\mem<14><5> ), .B(n1194), .Y(n264) );
  INVX1 U372 ( .A(n264), .Y(n265) );
  AND2X2 U373 ( .A(\mem<14><6> ), .B(n1194), .Y(n266) );
  INVX1 U374 ( .A(n266), .Y(n267) );
  AND2X2 U375 ( .A(\mem<14><7> ), .B(n1194), .Y(n268) );
  INVX1 U376 ( .A(n268), .Y(n269) );
  AND2X2 U377 ( .A(\mem<14><8> ), .B(n1193), .Y(n270) );
  INVX1 U378 ( .A(n270), .Y(n271) );
  AND2X2 U379 ( .A(\mem<14><9> ), .B(n1193), .Y(n272) );
  INVX1 U380 ( .A(n272), .Y(n273) );
  AND2X2 U381 ( .A(\mem<14><10> ), .B(n1193), .Y(n274) );
  INVX1 U382 ( .A(n274), .Y(n275) );
  AND2X2 U383 ( .A(\mem<14><11> ), .B(n1193), .Y(n276) );
  INVX1 U384 ( .A(n276), .Y(n277) );
  AND2X2 U385 ( .A(\mem<14><12> ), .B(n1193), .Y(n278) );
  INVX1 U386 ( .A(n278), .Y(n279) );
  AND2X2 U387 ( .A(\mem<14><13> ), .B(n1193), .Y(n280) );
  INVX1 U388 ( .A(n280), .Y(n281) );
  AND2X2 U389 ( .A(\mem<14><14> ), .B(n1193), .Y(n282) );
  INVX1 U390 ( .A(n282), .Y(n283) );
  AND2X2 U391 ( .A(\mem<14><15> ), .B(n1193), .Y(n284) );
  INVX1 U392 ( .A(n284), .Y(n285) );
  AND2X2 U393 ( .A(\mem<13><0> ), .B(n1197), .Y(n286) );
  INVX1 U394 ( .A(n286), .Y(n287) );
  AND2X2 U395 ( .A(\mem<13><1> ), .B(n1197), .Y(n288) );
  INVX1 U396 ( .A(n288), .Y(n289) );
  AND2X2 U397 ( .A(\mem<13><2> ), .B(n1197), .Y(n290) );
  INVX1 U398 ( .A(n290), .Y(n291) );
  AND2X2 U399 ( .A(\mem<13><3> ), .B(n1197), .Y(n292) );
  INVX1 U400 ( .A(n292), .Y(n293) );
  AND2X2 U401 ( .A(\mem<13><4> ), .B(n1197), .Y(n294) );
  INVX1 U402 ( .A(n294), .Y(n295) );
  AND2X2 U403 ( .A(\mem<13><5> ), .B(n1197), .Y(n296) );
  INVX1 U404 ( .A(n296), .Y(n297) );
  AND2X2 U405 ( .A(\mem<13><6> ), .B(n1197), .Y(n298) );
  INVX1 U406 ( .A(n298), .Y(n299) );
  AND2X2 U407 ( .A(\mem<13><7> ), .B(n1197), .Y(n300) );
  INVX1 U408 ( .A(n300), .Y(n301) );
  AND2X2 U409 ( .A(\mem<13><8> ), .B(n1196), .Y(n302) );
  INVX1 U410 ( .A(n302), .Y(n303) );
  AND2X2 U411 ( .A(\mem<13><9> ), .B(n1196), .Y(n304) );
  INVX1 U412 ( .A(n304), .Y(n305) );
  AND2X2 U413 ( .A(\mem<13><10> ), .B(n1196), .Y(n306) );
  INVX1 U414 ( .A(n306), .Y(n307) );
  AND2X2 U415 ( .A(\mem<13><11> ), .B(n1196), .Y(n308) );
  INVX1 U416 ( .A(n308), .Y(n309) );
  AND2X2 U417 ( .A(\mem<13><12> ), .B(n1196), .Y(n310) );
  INVX1 U418 ( .A(n310), .Y(n311) );
  AND2X2 U419 ( .A(\mem<13><13> ), .B(n1196), .Y(n312) );
  INVX1 U420 ( .A(n312), .Y(n313) );
  AND2X2 U421 ( .A(\mem<13><14> ), .B(n1196), .Y(n314) );
  INVX1 U422 ( .A(n314), .Y(n315) );
  AND2X2 U423 ( .A(\mem<13><15> ), .B(n1196), .Y(n316) );
  INVX1 U424 ( .A(n316), .Y(n317) );
  AND2X2 U425 ( .A(\mem<12><0> ), .B(n1200), .Y(n318) );
  INVX1 U426 ( .A(n318), .Y(n319) );
  AND2X2 U427 ( .A(\mem<12><1> ), .B(n1200), .Y(n320) );
  INVX1 U428 ( .A(n320), .Y(n321) );
  AND2X2 U429 ( .A(\mem<12><2> ), .B(n1200), .Y(n322) );
  INVX1 U430 ( .A(n322), .Y(n323) );
  AND2X2 U431 ( .A(\mem<12><3> ), .B(n1200), .Y(n324) );
  INVX1 U432 ( .A(n324), .Y(n325) );
  AND2X2 U433 ( .A(\mem<12><4> ), .B(n1200), .Y(n326) );
  INVX1 U434 ( .A(n326), .Y(n327) );
  AND2X2 U435 ( .A(\mem<12><5> ), .B(n1200), .Y(n328) );
  INVX1 U436 ( .A(n328), .Y(n329) );
  AND2X2 U437 ( .A(\mem<12><6> ), .B(n1200), .Y(n330) );
  INVX1 U438 ( .A(n330), .Y(n331) );
  AND2X2 U439 ( .A(\mem<12><7> ), .B(n1200), .Y(n332) );
  INVX1 U440 ( .A(n332), .Y(n333) );
  AND2X2 U441 ( .A(\mem<12><8> ), .B(n1199), .Y(n334) );
  INVX1 U442 ( .A(n334), .Y(n335) );
  AND2X2 U443 ( .A(\mem<12><9> ), .B(n1199), .Y(n336) );
  INVX1 U444 ( .A(n336), .Y(n337) );
  AND2X2 U445 ( .A(\mem<12><10> ), .B(n1199), .Y(n338) );
  INVX1 U446 ( .A(n338), .Y(n339) );
  AND2X2 U447 ( .A(\mem<12><11> ), .B(n1199), .Y(n340) );
  INVX1 U448 ( .A(n340), .Y(n341) );
  AND2X2 U449 ( .A(\mem<12><12> ), .B(n1199), .Y(n342) );
  INVX1 U450 ( .A(n342), .Y(n343) );
  AND2X2 U451 ( .A(\mem<12><13> ), .B(n1199), .Y(n344) );
  INVX1 U452 ( .A(n344), .Y(n345) );
  AND2X2 U453 ( .A(\mem<12><14> ), .B(n1199), .Y(n346) );
  INVX1 U454 ( .A(n346), .Y(n347) );
  AND2X2 U455 ( .A(\mem<12><15> ), .B(n1199), .Y(n348) );
  INVX1 U456 ( .A(n348), .Y(n349) );
  AND2X2 U457 ( .A(\mem<11><0> ), .B(n1203), .Y(n350) );
  INVX1 U458 ( .A(n350), .Y(n351) );
  AND2X2 U459 ( .A(\mem<11><1> ), .B(n1203), .Y(n352) );
  INVX1 U460 ( .A(n352), .Y(n353) );
  AND2X2 U461 ( .A(\mem<11><2> ), .B(n1203), .Y(n354) );
  INVX1 U462 ( .A(n354), .Y(n355) );
  AND2X2 U463 ( .A(\mem<11><3> ), .B(n1203), .Y(n356) );
  INVX1 U464 ( .A(n356), .Y(n357) );
  AND2X2 U465 ( .A(\mem<11><4> ), .B(n1203), .Y(n358) );
  INVX1 U466 ( .A(n358), .Y(n359) );
  AND2X2 U467 ( .A(\mem<11><5> ), .B(n1203), .Y(n360) );
  INVX1 U468 ( .A(n360), .Y(n361) );
  AND2X2 U469 ( .A(\mem<11><6> ), .B(n1203), .Y(n362) );
  INVX1 U470 ( .A(n362), .Y(n363) );
  AND2X2 U471 ( .A(\mem<11><7> ), .B(n1203), .Y(n364) );
  INVX1 U472 ( .A(n364), .Y(n365) );
  AND2X2 U473 ( .A(\mem<11><8> ), .B(n1202), .Y(n366) );
  INVX1 U474 ( .A(n366), .Y(n367) );
  AND2X2 U475 ( .A(\mem<11><9> ), .B(n1202), .Y(n368) );
  INVX1 U476 ( .A(n368), .Y(n369) );
  AND2X2 U477 ( .A(\mem<11><10> ), .B(n1202), .Y(n370) );
  INVX1 U478 ( .A(n370), .Y(n371) );
  AND2X2 U479 ( .A(\mem<11><11> ), .B(n1202), .Y(n372) );
  INVX1 U480 ( .A(n372), .Y(n373) );
  AND2X2 U481 ( .A(\mem<11><12> ), .B(n1202), .Y(n374) );
  INVX1 U482 ( .A(n374), .Y(n375) );
  AND2X2 U483 ( .A(\mem<11><13> ), .B(n1202), .Y(n376) );
  INVX1 U484 ( .A(n376), .Y(n377) );
  AND2X2 U485 ( .A(\mem<11><14> ), .B(n1202), .Y(n378) );
  INVX1 U486 ( .A(n378), .Y(n379) );
  AND2X2 U487 ( .A(\mem<11><15> ), .B(n1202), .Y(n380) );
  INVX1 U488 ( .A(n380), .Y(n381) );
  AND2X2 U489 ( .A(\mem<10><0> ), .B(n1206), .Y(n382) );
  INVX1 U490 ( .A(n382), .Y(n383) );
  AND2X2 U491 ( .A(\mem<10><1> ), .B(n1206), .Y(n384) );
  INVX1 U492 ( .A(n384), .Y(n385) );
  AND2X2 U493 ( .A(\mem<10><2> ), .B(n1206), .Y(n386) );
  INVX1 U494 ( .A(n386), .Y(n387) );
  AND2X2 U495 ( .A(\mem<10><3> ), .B(n1206), .Y(n388) );
  INVX1 U496 ( .A(n388), .Y(n389) );
  AND2X2 U497 ( .A(\mem<10><4> ), .B(n1206), .Y(n390) );
  INVX1 U498 ( .A(n390), .Y(n391) );
  AND2X2 U499 ( .A(\mem<10><5> ), .B(n1206), .Y(n392) );
  INVX1 U500 ( .A(n392), .Y(n393) );
  AND2X2 U501 ( .A(\mem<10><6> ), .B(n1206), .Y(n394) );
  INVX1 U502 ( .A(n394), .Y(n395) );
  AND2X2 U503 ( .A(\mem<10><7> ), .B(n1206), .Y(n396) );
  INVX1 U504 ( .A(n396), .Y(n397) );
  AND2X2 U505 ( .A(\mem<10><8> ), .B(n1205), .Y(n398) );
  INVX1 U506 ( .A(n398), .Y(n399) );
  AND2X2 U507 ( .A(\mem<10><9> ), .B(n1205), .Y(n400) );
  INVX1 U508 ( .A(n400), .Y(n401) );
  AND2X2 U509 ( .A(\mem<10><10> ), .B(n1205), .Y(n402) );
  INVX1 U510 ( .A(n402), .Y(n403) );
  AND2X2 U511 ( .A(\mem<10><11> ), .B(n1205), .Y(n404) );
  INVX1 U512 ( .A(n404), .Y(n405) );
  AND2X2 U513 ( .A(\mem<10><12> ), .B(n1205), .Y(n406) );
  INVX1 U514 ( .A(n406), .Y(n407) );
  AND2X2 U515 ( .A(\mem<10><13> ), .B(n1205), .Y(n408) );
  INVX1 U516 ( .A(n408), .Y(n409) );
  AND2X2 U517 ( .A(\mem<10><14> ), .B(n1205), .Y(n410) );
  INVX1 U518 ( .A(n410), .Y(n411) );
  AND2X2 U519 ( .A(\mem<10><15> ), .B(n1205), .Y(n412) );
  INVX1 U520 ( .A(n412), .Y(n413) );
  AND2X2 U521 ( .A(\mem<9><0> ), .B(n1209), .Y(n414) );
  INVX1 U522 ( .A(n414), .Y(n415) );
  AND2X2 U523 ( .A(\mem<9><1> ), .B(n1209), .Y(n416) );
  INVX1 U524 ( .A(n416), .Y(n417) );
  AND2X2 U525 ( .A(\mem<9><2> ), .B(n1209), .Y(n418) );
  INVX1 U526 ( .A(n418), .Y(n419) );
  AND2X2 U527 ( .A(\mem<9><3> ), .B(n1209), .Y(n420) );
  INVX1 U528 ( .A(n420), .Y(n421) );
  AND2X2 U529 ( .A(\mem<9><4> ), .B(n1209), .Y(n422) );
  INVX1 U530 ( .A(n422), .Y(n423) );
  AND2X2 U531 ( .A(\mem<9><5> ), .B(n1209), .Y(n424) );
  INVX1 U532 ( .A(n424), .Y(n425) );
  AND2X2 U533 ( .A(\mem<9><6> ), .B(n1209), .Y(n426) );
  INVX1 U534 ( .A(n426), .Y(n427) );
  AND2X2 U535 ( .A(\mem<9><7> ), .B(n1209), .Y(n428) );
  INVX1 U536 ( .A(n428), .Y(n429) );
  AND2X2 U537 ( .A(\mem<9><8> ), .B(n1208), .Y(n430) );
  INVX1 U538 ( .A(n430), .Y(n431) );
  AND2X2 U539 ( .A(\mem<9><9> ), .B(n1208), .Y(n432) );
  INVX1 U540 ( .A(n432), .Y(n433) );
  AND2X2 U541 ( .A(\mem<9><10> ), .B(n1208), .Y(n434) );
  INVX1 U542 ( .A(n434), .Y(n435) );
  AND2X2 U543 ( .A(\mem<9><11> ), .B(n1208), .Y(n436) );
  INVX1 U544 ( .A(n436), .Y(n437) );
  AND2X2 U545 ( .A(\mem<9><12> ), .B(n1208), .Y(n438) );
  INVX1 U546 ( .A(n438), .Y(n439) );
  AND2X2 U547 ( .A(\mem<9><13> ), .B(n1208), .Y(n440) );
  INVX1 U548 ( .A(n440), .Y(n441) );
  AND2X2 U549 ( .A(\mem<9><14> ), .B(n1208), .Y(n442) );
  INVX1 U550 ( .A(n442), .Y(n443) );
  AND2X2 U551 ( .A(\mem<9><15> ), .B(n1208), .Y(n444) );
  INVX1 U552 ( .A(n444), .Y(n445) );
  AND2X2 U553 ( .A(\mem<7><1> ), .B(n1211), .Y(n446) );
  INVX1 U554 ( .A(n446), .Y(n447) );
  AND2X2 U555 ( .A(\mem<7><2> ), .B(n1211), .Y(n448) );
  INVX1 U556 ( .A(n448), .Y(n449) );
  AND2X2 U557 ( .A(\mem<7><3> ), .B(n1211), .Y(n450) );
  INVX1 U558 ( .A(n450), .Y(n451) );
  AND2X2 U559 ( .A(\mem<7><4> ), .B(n1211), .Y(n452) );
  INVX1 U560 ( .A(n452), .Y(n453) );
  AND2X2 U561 ( .A(\mem<7><5> ), .B(n1211), .Y(n454) );
  INVX1 U562 ( .A(n454), .Y(n455) );
  AND2X2 U563 ( .A(\mem<7><6> ), .B(n1211), .Y(n456) );
  INVX1 U564 ( .A(n456), .Y(n457) );
  AND2X2 U565 ( .A(\mem<7><7> ), .B(n1211), .Y(n458) );
  INVX1 U566 ( .A(n458), .Y(n459) );
  AND2X2 U567 ( .A(\mem<7><8> ), .B(n1211), .Y(n460) );
  INVX1 U568 ( .A(n460), .Y(n461) );
  AND2X2 U569 ( .A(\mem<7><9> ), .B(n1211), .Y(n462) );
  INVX1 U570 ( .A(n462), .Y(n463) );
  AND2X2 U571 ( .A(\mem<7><10> ), .B(n1211), .Y(n464) );
  INVX1 U572 ( .A(n464), .Y(n465) );
  AND2X2 U573 ( .A(\mem<7><11> ), .B(n1211), .Y(n466) );
  INVX1 U574 ( .A(n466), .Y(n467) );
  AND2X2 U575 ( .A(\mem<7><12> ), .B(n1211), .Y(n468) );
  INVX1 U576 ( .A(n468), .Y(n469) );
  AND2X2 U577 ( .A(\mem<7><13> ), .B(n1211), .Y(n470) );
  INVX1 U578 ( .A(n470), .Y(n471) );
  AND2X2 U579 ( .A(\mem<7><14> ), .B(n1211), .Y(n472) );
  INVX1 U580 ( .A(n472), .Y(n473) );
  AND2X2 U581 ( .A(\mem<7><15> ), .B(n1211), .Y(n474) );
  INVX1 U582 ( .A(n474), .Y(n475) );
  AND2X2 U583 ( .A(\mem<6><1> ), .B(n1214), .Y(n476) );
  INVX1 U584 ( .A(n476), .Y(n477) );
  AND2X2 U585 ( .A(\mem<6><2> ), .B(n1214), .Y(n478) );
  INVX1 U586 ( .A(n478), .Y(n479) );
  AND2X2 U587 ( .A(\mem<6><3> ), .B(n1214), .Y(n480) );
  INVX1 U588 ( .A(n480), .Y(n481) );
  AND2X2 U589 ( .A(\mem<6><4> ), .B(n1214), .Y(n482) );
  INVX1 U590 ( .A(n482), .Y(n483) );
  AND2X2 U591 ( .A(\mem<6><5> ), .B(n1214), .Y(n484) );
  INVX1 U592 ( .A(n484), .Y(n485) );
  AND2X2 U593 ( .A(\mem<6><6> ), .B(n1214), .Y(n486) );
  INVX1 U594 ( .A(n486), .Y(n487) );
  AND2X2 U595 ( .A(\mem<6><7> ), .B(n1214), .Y(n488) );
  INVX1 U596 ( .A(n488), .Y(n489) );
  AND2X2 U597 ( .A(\mem<6><8> ), .B(n1213), .Y(n490) );
  INVX1 U598 ( .A(n490), .Y(n491) );
  AND2X2 U599 ( .A(\mem<6><9> ), .B(n1213), .Y(n492) );
  INVX1 U600 ( .A(n492), .Y(n493) );
  AND2X2 U601 ( .A(\mem<6><10> ), .B(n1213), .Y(n494) );
  INVX1 U602 ( .A(n494), .Y(n495) );
  AND2X2 U603 ( .A(\mem<6><11> ), .B(n1213), .Y(n496) );
  INVX1 U604 ( .A(n496), .Y(n497) );
  AND2X2 U605 ( .A(\mem<6><12> ), .B(n1213), .Y(n498) );
  INVX1 U606 ( .A(n498), .Y(n499) );
  AND2X2 U607 ( .A(\mem<6><13> ), .B(n1213), .Y(n500) );
  INVX1 U608 ( .A(n500), .Y(n501) );
  AND2X2 U609 ( .A(\mem<6><14> ), .B(n1213), .Y(n502) );
  INVX1 U610 ( .A(n502), .Y(n503) );
  AND2X2 U611 ( .A(\mem<6><15> ), .B(n1213), .Y(n504) );
  INVX1 U612 ( .A(n504), .Y(n505) );
  AND2X2 U613 ( .A(\mem<5><8> ), .B(n1216), .Y(n506) );
  INVX1 U614 ( .A(n506), .Y(n507) );
  AND2X2 U615 ( .A(\mem<5><9> ), .B(n1216), .Y(n508) );
  INVX1 U616 ( .A(n508), .Y(n509) );
  AND2X2 U617 ( .A(\mem<5><10> ), .B(n1216), .Y(n510) );
  INVX1 U618 ( .A(n510), .Y(n511) );
  AND2X2 U619 ( .A(\mem<5><11> ), .B(n1216), .Y(n512) );
  INVX1 U620 ( .A(n512), .Y(n513) );
  AND2X2 U621 ( .A(\mem<5><12> ), .B(n1216), .Y(n514) );
  INVX1 U622 ( .A(n514), .Y(n515) );
  AND2X2 U623 ( .A(\mem<5><13> ), .B(n1216), .Y(n516) );
  INVX1 U624 ( .A(n516), .Y(n517) );
  AND2X2 U625 ( .A(\mem<5><14> ), .B(n1216), .Y(n518) );
  INVX1 U626 ( .A(n518), .Y(n519) );
  AND2X2 U627 ( .A(\mem<5><15> ), .B(n1216), .Y(n520) );
  INVX1 U628 ( .A(n520), .Y(n521) );
  AND2X2 U629 ( .A(\mem<4><1> ), .B(n1220), .Y(n522) );
  INVX1 U630 ( .A(n522), .Y(n523) );
  AND2X2 U631 ( .A(\mem<4><2> ), .B(n1220), .Y(n524) );
  INVX1 U632 ( .A(n524), .Y(n525) );
  AND2X2 U633 ( .A(\mem<4><3> ), .B(n1220), .Y(n526) );
  INVX1 U634 ( .A(n526), .Y(n527) );
  AND2X2 U635 ( .A(\mem<4><4> ), .B(n1220), .Y(n528) );
  INVX1 U636 ( .A(n528), .Y(n529) );
  AND2X2 U637 ( .A(\mem<4><5> ), .B(n1220), .Y(n530) );
  INVX1 U638 ( .A(n530), .Y(n531) );
  AND2X2 U639 ( .A(\mem<4><6> ), .B(n1220), .Y(n532) );
  INVX1 U640 ( .A(n532), .Y(n533) );
  AND2X2 U641 ( .A(\mem<4><7> ), .B(n1220), .Y(n534) );
  INVX1 U642 ( .A(n534), .Y(n535) );
  AND2X2 U643 ( .A(\mem<4><8> ), .B(n1219), .Y(n536) );
  INVX1 U644 ( .A(n536), .Y(n537) );
  AND2X2 U645 ( .A(\mem<4><9> ), .B(n1219), .Y(n538) );
  INVX1 U646 ( .A(n538), .Y(n539) );
  AND2X2 U647 ( .A(\mem<4><10> ), .B(n1219), .Y(n540) );
  INVX1 U648 ( .A(n540), .Y(n541) );
  AND2X2 U649 ( .A(\mem<4><11> ), .B(n1219), .Y(n542) );
  INVX1 U650 ( .A(n542), .Y(n543) );
  AND2X2 U651 ( .A(\mem<4><12> ), .B(n1219), .Y(n544) );
  INVX1 U652 ( .A(n544), .Y(n545) );
  AND2X2 U653 ( .A(\mem<4><13> ), .B(n1219), .Y(n546) );
  INVX1 U654 ( .A(n546), .Y(n547) );
  AND2X2 U655 ( .A(\mem<4><14> ), .B(n1219), .Y(n548) );
  INVX1 U656 ( .A(n548), .Y(n549) );
  AND2X2 U657 ( .A(\mem<4><15> ), .B(n1219), .Y(n550) );
  INVX1 U658 ( .A(n550), .Y(n551) );
  AND2X2 U659 ( .A(\mem<3><1> ), .B(n1223), .Y(n552) );
  INVX1 U660 ( .A(n552), .Y(n553) );
  AND2X2 U661 ( .A(\mem<3><2> ), .B(n1223), .Y(n554) );
  INVX1 U662 ( .A(n554), .Y(n555) );
  AND2X2 U663 ( .A(\mem<3><3> ), .B(n1223), .Y(n556) );
  INVX1 U664 ( .A(n556), .Y(n557) );
  AND2X2 U665 ( .A(\mem<3><4> ), .B(n1223), .Y(n558) );
  INVX1 U666 ( .A(n558), .Y(n559) );
  AND2X2 U667 ( .A(\mem<3><5> ), .B(n1223), .Y(n560) );
  INVX1 U668 ( .A(n560), .Y(n561) );
  AND2X2 U669 ( .A(\mem<3><6> ), .B(n1223), .Y(n562) );
  INVX1 U670 ( .A(n562), .Y(n563) );
  AND2X2 U671 ( .A(\mem<3><7> ), .B(n1223), .Y(n564) );
  INVX1 U672 ( .A(n564), .Y(n565) );
  AND2X2 U673 ( .A(\mem<3><15> ), .B(n1222), .Y(n566) );
  INVX1 U674 ( .A(n566), .Y(n567) );
  AND2X2 U675 ( .A(\mem<2><8> ), .B(n1225), .Y(n568) );
  INVX1 U676 ( .A(n568), .Y(n569) );
  AND2X2 U677 ( .A(\mem<2><9> ), .B(n1225), .Y(n570) );
  INVX1 U678 ( .A(n570), .Y(n571) );
  AND2X2 U679 ( .A(\mem<2><10> ), .B(n1225), .Y(n572) );
  INVX1 U680 ( .A(n572), .Y(n573) );
  AND2X2 U681 ( .A(\mem<2><11> ), .B(n1225), .Y(n574) );
  INVX1 U682 ( .A(n574), .Y(n575) );
  AND2X2 U683 ( .A(\mem<2><12> ), .B(n1225), .Y(n576) );
  INVX1 U684 ( .A(n576), .Y(n577) );
  AND2X2 U685 ( .A(\mem<2><13> ), .B(n1225), .Y(n578) );
  INVX1 U686 ( .A(n578), .Y(n579) );
  AND2X2 U687 ( .A(\mem<2><14> ), .B(n1225), .Y(n580) );
  INVX1 U688 ( .A(n580), .Y(n581) );
  AND2X2 U689 ( .A(\mem<2><15> ), .B(n1225), .Y(n582) );
  INVX1 U690 ( .A(n582), .Y(n583) );
  AND2X2 U691 ( .A(\mem<1><1> ), .B(n1229), .Y(n584) );
  INVX1 U692 ( .A(n584), .Y(n585) );
  AND2X2 U693 ( .A(\mem<1><2> ), .B(n1229), .Y(n586) );
  INVX1 U694 ( .A(n586), .Y(n587) );
  AND2X2 U695 ( .A(\mem<1><3> ), .B(n1229), .Y(n588) );
  INVX1 U696 ( .A(n588), .Y(n589) );
  AND2X2 U697 ( .A(\mem<1><4> ), .B(n1229), .Y(n590) );
  INVX1 U698 ( .A(n590), .Y(n591) );
  AND2X2 U699 ( .A(\mem<1><5> ), .B(n1229), .Y(n592) );
  INVX1 U700 ( .A(n592), .Y(n593) );
  AND2X2 U701 ( .A(\mem<1><6> ), .B(n1229), .Y(n594) );
  INVX1 U702 ( .A(n594), .Y(n595) );
  AND2X2 U703 ( .A(\mem<1><7> ), .B(n1229), .Y(n596) );
  INVX1 U704 ( .A(n596), .Y(n597) );
  AND2X2 U705 ( .A(\mem<1><8> ), .B(n1228), .Y(n598) );
  INVX1 U706 ( .A(n598), .Y(n599) );
  AND2X2 U707 ( .A(\mem<1><9> ), .B(n1228), .Y(n600) );
  INVX1 U708 ( .A(n600), .Y(n601) );
  AND2X2 U709 ( .A(\mem<1><10> ), .B(n1228), .Y(n602) );
  INVX1 U710 ( .A(n602), .Y(n603) );
  AND2X2 U711 ( .A(\mem<1><11> ), .B(n1228), .Y(n604) );
  INVX1 U712 ( .A(n604), .Y(n605) );
  AND2X2 U713 ( .A(\mem<1><12> ), .B(n1228), .Y(n606) );
  INVX1 U714 ( .A(n606), .Y(n607) );
  AND2X2 U715 ( .A(\mem<1><13> ), .B(n1228), .Y(n608) );
  INVX1 U716 ( .A(n608), .Y(n609) );
  AND2X2 U717 ( .A(\mem<1><14> ), .B(n1228), .Y(n610) );
  INVX1 U718 ( .A(n610), .Y(n611) );
  AND2X2 U719 ( .A(\mem<1><15> ), .B(n1228), .Y(n612) );
  INVX1 U720 ( .A(n612), .Y(n613) );
  AND2X2 U721 ( .A(n1921), .B(n1274), .Y(n614) );
  AND2X2 U722 ( .A(n1922), .B(n1276), .Y(n616) );
  AND2X2 U723 ( .A(n1923), .B(n1252), .Y(n618) );
  AND2X2 U724 ( .A(n1922), .B(n1253), .Y(n620) );
  AND2X2 U725 ( .A(n1957), .B(n1311), .Y(n622) );
  AND2X2 U726 ( .A(\data_in<0> ), .B(n1922), .Y(n623) );
  AND2X2 U727 ( .A(\data_in<1> ), .B(n1923), .Y(n624) );
  AND2X2 U728 ( .A(\data_in<2> ), .B(n1922), .Y(n625) );
  AND2X2 U729 ( .A(\data_in<3> ), .B(n1922), .Y(n626) );
  AND2X2 U730 ( .A(\data_in<4> ), .B(n1922), .Y(n627) );
  AND2X2 U731 ( .A(\data_in<5> ), .B(n1923), .Y(n628) );
  AND2X2 U732 ( .A(\data_in<6> ), .B(n1923), .Y(n629) );
  AND2X2 U733 ( .A(\data_in<7> ), .B(n1923), .Y(n630) );
  AND2X2 U734 ( .A(\data_in<8> ), .B(n1922), .Y(n631) );
  AND2X2 U735 ( .A(\data_in<9> ), .B(n1922), .Y(n632) );
  AND2X2 U736 ( .A(\data_in<10> ), .B(n1923), .Y(n633) );
  AND2X2 U737 ( .A(\data_in<11> ), .B(n1923), .Y(n634) );
  AND2X2 U738 ( .A(\data_in<12> ), .B(n1923), .Y(n635) );
  AND2X2 U739 ( .A(\data_in<13> ), .B(n1923), .Y(n636) );
  AND2X2 U740 ( .A(\data_in<14> ), .B(n1923), .Y(n637) );
  AND2X2 U741 ( .A(\data_in<15> ), .B(n1923), .Y(n638) );
  AND2X2 U742 ( .A(n1921), .B(n1254), .Y(n639) );
  AND2X2 U743 ( .A(n1921), .B(n1256), .Y(n641) );
  AND2X2 U744 ( .A(n1921), .B(n1258), .Y(n643) );
  INVX1 U745 ( .A(n643), .Y(n644) );
  INVX1 U746 ( .A(n643), .Y(n645) );
  AND2X2 U747 ( .A(n1921), .B(n1260), .Y(n646) );
  INVX1 U748 ( .A(n646), .Y(n647) );
  INVX1 U749 ( .A(n646), .Y(n648) );
  AND2X2 U750 ( .A(n1921), .B(n1262), .Y(n649) );
  INVX1 U751 ( .A(n649), .Y(n650) );
  INVX1 U752 ( .A(n649), .Y(n1163) );
  AND2X2 U753 ( .A(n1921), .B(n1264), .Y(n1164) );
  INVX1 U754 ( .A(n1164), .Y(n1165) );
  INVX1 U755 ( .A(n1164), .Y(n1166) );
  AND2X2 U756 ( .A(n1921), .B(n1266), .Y(n1167) );
  INVX1 U757 ( .A(n1167), .Y(n1168) );
  INVX1 U758 ( .A(n1167), .Y(n1169) );
  AND2X2 U759 ( .A(n1921), .B(n1249), .Y(n1170) );
  INVX1 U760 ( .A(n1170), .Y(n1171) );
  INVX1 U761 ( .A(n1170), .Y(n1172) );
  AND2X2 U762 ( .A(n1921), .B(n1268), .Y(n1173) );
  INVX1 U763 ( .A(n1173), .Y(n1174) );
  INVX1 U764 ( .A(n1173), .Y(n1175) );
  AND2X2 U765 ( .A(n1921), .B(n1270), .Y(n1176) );
  INVX1 U766 ( .A(n1176), .Y(n1177) );
  INVX1 U767 ( .A(n1176), .Y(n1178) );
  AND2X2 U768 ( .A(n1921), .B(n1272), .Y(n1179) );
  INVX1 U769 ( .A(n1179), .Y(n1180) );
  INVX1 U770 ( .A(n1179), .Y(n1181) );
  AND2X2 U771 ( .A(n1922), .B(n1278), .Y(n1182) );
  AND2X2 U772 ( .A(n1922), .B(n1280), .Y(n1184) );
  AND2X2 U773 ( .A(n1922), .B(n1251), .Y(n1186) );
  INVX1 U774 ( .A(n1186), .Y(n1187) );
  INVX1 U775 ( .A(n1186), .Y(n1188) );
  AND2X2 U776 ( .A(n1922), .B(n1282), .Y(n1189) );
  INVX1 U777 ( .A(n1189), .Y(n1190) );
  INVX1 U778 ( .A(n1189), .Y(n1191) );
  AND2X2 U779 ( .A(n1922), .B(n1284), .Y(n1192) );
  INVX1 U780 ( .A(n1192), .Y(n1193) );
  INVX1 U781 ( .A(n1192), .Y(n1194) );
  AND2X2 U782 ( .A(n1922), .B(n1286), .Y(n1195) );
  INVX1 U783 ( .A(n1195), .Y(n1196) );
  INVX1 U784 ( .A(n1195), .Y(n1197) );
  AND2X2 U785 ( .A(n1922), .B(n1288), .Y(n1198) );
  INVX1 U786 ( .A(n1198), .Y(n1199) );
  INVX1 U787 ( .A(n1198), .Y(n1200) );
  AND2X2 U788 ( .A(n1922), .B(n1290), .Y(n1201) );
  INVX1 U789 ( .A(n1201), .Y(n1202) );
  INVX1 U790 ( .A(n1201), .Y(n1203) );
  AND2X2 U791 ( .A(n1922), .B(n1292), .Y(n1204) );
  INVX1 U792 ( .A(n1204), .Y(n1205) );
  INVX1 U793 ( .A(n1204), .Y(n1206) );
  AND2X2 U794 ( .A(n1922), .B(n1294), .Y(n1207) );
  INVX1 U795 ( .A(n1207), .Y(n1208) );
  INVX1 U796 ( .A(n1207), .Y(n1209) );
  AND2X2 U797 ( .A(n1923), .B(n1296), .Y(n1210) );
  AND2X2 U798 ( .A(n1923), .B(n1298), .Y(n1212) );
  INVX1 U799 ( .A(n1212), .Y(n1213) );
  INVX1 U800 ( .A(n1212), .Y(n1214) );
  AND2X2 U801 ( .A(n1923), .B(n1300), .Y(n1215) );
  INVX1 U802 ( .A(n1215), .Y(n1216) );
  INVX1 U803 ( .A(n1215), .Y(n1217) );
  AND2X2 U804 ( .A(n1923), .B(n1302), .Y(n1218) );
  INVX1 U805 ( .A(n1218), .Y(n1219) );
  INVX1 U806 ( .A(n1218), .Y(n1220) );
  AND2X2 U807 ( .A(n1923), .B(n1304), .Y(n1221) );
  INVX1 U808 ( .A(n1221), .Y(n1222) );
  INVX1 U809 ( .A(n1221), .Y(n1223) );
  AND2X2 U810 ( .A(n1923), .B(n1306), .Y(n1224) );
  INVX1 U811 ( .A(n1224), .Y(n1225) );
  INVX1 U812 ( .A(n1224), .Y(n1226) );
  AND2X2 U813 ( .A(n1923), .B(n1308), .Y(n1227) );
  INVX1 U814 ( .A(n1227), .Y(n1228) );
  INVX1 U815 ( .A(n1227), .Y(n1229) );
  OR2X2 U816 ( .A(write), .B(rst), .Y(n1230) );
  OR2X2 U817 ( .A(write), .B(rst), .Y(n1232) );
  INVX1 U818 ( .A(n1232), .Y(n1233) );
  INVX1 U819 ( .A(n1232), .Y(n1234) );
  INVX1 U820 ( .A(n1232), .Y(n1235) );
  INVX1 U821 ( .A(n1959), .Y(n1958) );
  INVX4 U822 ( .A(n623), .Y(n1926) );
  INVX4 U823 ( .A(n624), .Y(n1928) );
  INVX4 U824 ( .A(n625), .Y(n1930) );
  INVX4 U825 ( .A(n626), .Y(n1932) );
  INVX4 U826 ( .A(n627), .Y(n1934) );
  INVX4 U827 ( .A(n628), .Y(n1936) );
  INVX4 U828 ( .A(n629), .Y(n1938) );
  INVX4 U829 ( .A(n630), .Y(n1940) );
  INVX4 U830 ( .A(n631), .Y(n1942) );
  INVX4 U831 ( .A(n632), .Y(n1944) );
  INVX4 U832 ( .A(n633), .Y(n1946) );
  INVX4 U833 ( .A(n634), .Y(n1948) );
  INVX4 U834 ( .A(n635), .Y(n1950) );
  INVX4 U835 ( .A(n636), .Y(n1952) );
  INVX4 U836 ( .A(n637), .Y(n1954) );
  INVX4 U837 ( .A(n638), .Y(n1956) );
  INVX1 U838 ( .A(n1963), .Y(n1962) );
  AND2X1 U839 ( .A(n1962), .B(n1960), .Y(n1236) );
  INVX1 U840 ( .A(n1961), .Y(n1960) );
  AND2X1 U841 ( .A(n2701), .B(n1966), .Y(n1237) );
  BUFX2 U842 ( .A(n1996), .Y(n1238) );
  INVX1 U843 ( .A(n1238), .Y(n2140) );
  BUFX2 U844 ( .A(n2012), .Y(n1239) );
  INVX1 U845 ( .A(n1239), .Y(n2149) );
  BUFX2 U846 ( .A(n2027), .Y(n1240) );
  INVX1 U847 ( .A(n1240), .Y(n2151) );
  BUFX2 U848 ( .A(n2042), .Y(n1241) );
  INVX1 U849 ( .A(n1241), .Y(n2160) );
  BUFX2 U850 ( .A(n2058), .Y(n1242) );
  INVX1 U851 ( .A(n1242), .Y(n2169) );
  BUFX2 U852 ( .A(n2119), .Y(n1243) );
  INVX1 U853 ( .A(n1243), .Y(n2120) );
  BUFX2 U854 ( .A(n2137), .Y(n1244) );
  INVX1 U855 ( .A(n1244), .Y(n2171) );
  AND2X1 U856 ( .A(n1958), .B(n1236), .Y(n1245) );
  AND2X1 U857 ( .A(n1964), .B(n1237), .Y(n1246) );
  AND2X1 U858 ( .A(n1959), .B(n1236), .Y(n1247) );
  AND2X1 U859 ( .A(n1965), .B(n1237), .Y(n1248) );
  AND2X1 U860 ( .A(n1246), .B(n2172), .Y(n1249) );
  INVX1 U861 ( .A(n1249), .Y(n1250) );
  AND2X1 U862 ( .A(n2172), .B(n1248), .Y(n1251) );
  AND2X1 U863 ( .A(n2172), .B(n2120), .Y(n1252) );
  AND2X1 U864 ( .A(n2172), .B(n2171), .Y(n1253) );
  AND2X1 U865 ( .A(n1245), .B(n1246), .Y(n1254) );
  INVX1 U866 ( .A(n1254), .Y(n1255) );
  AND2X1 U867 ( .A(n1246), .B(n1247), .Y(n1256) );
  INVX1 U868 ( .A(n1256), .Y(n1257) );
  AND2X1 U869 ( .A(n1246), .B(n2140), .Y(n1258) );
  INVX1 U870 ( .A(n1258), .Y(n1259) );
  AND2X1 U871 ( .A(n1246), .B(n2149), .Y(n1260) );
  INVX1 U872 ( .A(n1260), .Y(n1261) );
  AND2X1 U873 ( .A(n1246), .B(n2151), .Y(n1262) );
  INVX1 U874 ( .A(n1262), .Y(n1263) );
  AND2X1 U875 ( .A(n1246), .B(n2160), .Y(n1264) );
  INVX1 U876 ( .A(n1264), .Y(n1265) );
  AND2X1 U877 ( .A(n1246), .B(n2169), .Y(n1266) );
  INVX1 U878 ( .A(n1266), .Y(n1267) );
  AND2X1 U879 ( .A(n1245), .B(n1248), .Y(n1268) );
  INVX1 U880 ( .A(n1268), .Y(n1269) );
  AND2X1 U881 ( .A(n1247), .B(n1248), .Y(n1270) );
  INVX1 U882 ( .A(n1270), .Y(n1271) );
  AND2X1 U883 ( .A(n2140), .B(n1248), .Y(n1272) );
  INVX1 U884 ( .A(n1272), .Y(n1273) );
  AND2X1 U885 ( .A(n2149), .B(n1248), .Y(n1274) );
  INVX1 U886 ( .A(n1274), .Y(n1275) );
  AND2X1 U887 ( .A(n2151), .B(n1248), .Y(n1276) );
  INVX1 U888 ( .A(n1276), .Y(n1277) );
  AND2X1 U889 ( .A(n2160), .B(n1248), .Y(n1278) );
  INVX1 U890 ( .A(n1278), .Y(n1279) );
  AND2X1 U891 ( .A(n2169), .B(n1248), .Y(n1280) );
  INVX1 U892 ( .A(n1280), .Y(n1281) );
  AND2X1 U893 ( .A(n1245), .B(n2120), .Y(n1282) );
  INVX1 U894 ( .A(n1282), .Y(n1283) );
  AND2X1 U895 ( .A(n1247), .B(n2120), .Y(n1284) );
  INVX1 U896 ( .A(n1284), .Y(n1285) );
  AND2X1 U897 ( .A(n2140), .B(n2120), .Y(n1286) );
  INVX1 U898 ( .A(n1286), .Y(n1287) );
  AND2X1 U899 ( .A(n2149), .B(n2120), .Y(n1288) );
  INVX1 U900 ( .A(n1288), .Y(n1289) );
  AND2X1 U901 ( .A(n2151), .B(n2120), .Y(n1290) );
  INVX1 U902 ( .A(n1290), .Y(n1291) );
  AND2X1 U903 ( .A(n2160), .B(n2120), .Y(n1292) );
  INVX1 U904 ( .A(n1292), .Y(n1293) );
  AND2X1 U905 ( .A(n2169), .B(n2120), .Y(n1294) );
  INVX1 U906 ( .A(n1294), .Y(n1295) );
  AND2X1 U907 ( .A(n1245), .B(n2171), .Y(n1296) );
  INVX1 U908 ( .A(n1296), .Y(n1297) );
  AND2X1 U909 ( .A(n1247), .B(n2171), .Y(n1298) );
  INVX1 U910 ( .A(n1298), .Y(n1299) );
  AND2X1 U911 ( .A(n2140), .B(n2171), .Y(n1300) );
  INVX1 U912 ( .A(n1300), .Y(n1301) );
  AND2X1 U913 ( .A(n2149), .B(n2171), .Y(n1302) );
  INVX1 U914 ( .A(n1302), .Y(n1303) );
  AND2X1 U915 ( .A(n2151), .B(n2171), .Y(n1304) );
  INVX1 U916 ( .A(n1304), .Y(n1305) );
  AND2X1 U917 ( .A(n2160), .B(n2171), .Y(n1306) );
  INVX1 U918 ( .A(n1306), .Y(n1307) );
  AND2X1 U919 ( .A(n2169), .B(n2171), .Y(n1308) );
  INVX1 U920 ( .A(n1308), .Y(n1309) );
  INVX1 U921 ( .A(N12), .Y(n1963) );
  INVX1 U922 ( .A(write), .Y(n1310) );
  INVX1 U923 ( .A(n1310), .Y(n1311) );
  MUX2X1 U924 ( .B(n1313), .A(n1314), .S(n1821), .Y(n1312) );
  MUX2X1 U925 ( .B(n1316), .A(n1317), .S(n1821), .Y(n1315) );
  MUX2X1 U926 ( .B(n1319), .A(n1320), .S(n1821), .Y(n1318) );
  MUX2X1 U927 ( .B(n1322), .A(n1323), .S(n1821), .Y(n1321) );
  MUX2X1 U928 ( .B(n1325), .A(n1326), .S(n1811), .Y(n1324) );
  MUX2X1 U929 ( .B(n1328), .A(n1329), .S(n1821), .Y(n1327) );
  MUX2X1 U930 ( .B(n1331), .A(n1332), .S(n1821), .Y(n1330) );
  MUX2X1 U931 ( .B(n1334), .A(n1335), .S(n1821), .Y(n1333) );
  MUX2X1 U932 ( .B(n1337), .A(n1338), .S(n1821), .Y(n1336) );
  MUX2X1 U933 ( .B(n1340), .A(n1341), .S(n1811), .Y(n1339) );
  MUX2X1 U934 ( .B(n1343), .A(n1344), .S(n1822), .Y(n1342) );
  MUX2X1 U935 ( .B(n1346), .A(n1347), .S(n1822), .Y(n1345) );
  MUX2X1 U936 ( .B(n1349), .A(n1350), .S(n1822), .Y(n1348) );
  MUX2X1 U937 ( .B(n1352), .A(n1353), .S(n1822), .Y(n1351) );
  MUX2X1 U938 ( .B(n1355), .A(n1356), .S(n1811), .Y(n1354) );
  MUX2X1 U939 ( .B(n1358), .A(n1359), .S(n1822), .Y(n1357) );
  MUX2X1 U940 ( .B(n1361), .A(n1362), .S(n1822), .Y(n1360) );
  MUX2X1 U941 ( .B(n1364), .A(n1365), .S(n1822), .Y(n1363) );
  MUX2X1 U942 ( .B(n1367), .A(n1368), .S(n1822), .Y(n1366) );
  MUX2X1 U943 ( .B(n1370), .A(n1371), .S(n1811), .Y(n1369) );
  MUX2X1 U944 ( .B(n1373), .A(n1374), .S(n1822), .Y(n1372) );
  MUX2X1 U945 ( .B(n1376), .A(n1377), .S(n1822), .Y(n1375) );
  MUX2X1 U946 ( .B(n1379), .A(n1380), .S(n1822), .Y(n1378) );
  MUX2X1 U947 ( .B(n1382), .A(n1383), .S(n1822), .Y(n1381) );
  MUX2X1 U948 ( .B(n1385), .A(n1386), .S(n1811), .Y(n1384) );
  MUX2X1 U949 ( .B(n1388), .A(n1389), .S(n1823), .Y(n1387) );
  MUX2X1 U950 ( .B(n1391), .A(n1392), .S(n1823), .Y(n1390) );
  MUX2X1 U951 ( .B(n1394), .A(n1395), .S(n1823), .Y(n1393) );
  MUX2X1 U952 ( .B(n1397), .A(n1398), .S(n1823), .Y(n1396) );
  MUX2X1 U953 ( .B(n1400), .A(n1401), .S(n1811), .Y(n1399) );
  MUX2X1 U954 ( .B(n1403), .A(n1404), .S(n1823), .Y(n1402) );
  MUX2X1 U955 ( .B(n1406), .A(n1407), .S(n1823), .Y(n1405) );
  MUX2X1 U956 ( .B(n1409), .A(n1410), .S(n1823), .Y(n1408) );
  MUX2X1 U957 ( .B(n1412), .A(n1413), .S(n1823), .Y(n1411) );
  MUX2X1 U958 ( .B(n1415), .A(n1416), .S(n1811), .Y(n1414) );
  MUX2X1 U959 ( .B(n1418), .A(n1419), .S(n1823), .Y(n1417) );
  MUX2X1 U960 ( .B(n1421), .A(n1422), .S(n1823), .Y(n1420) );
  MUX2X1 U961 ( .B(n1424), .A(n1425), .S(n1823), .Y(n1423) );
  MUX2X1 U962 ( .B(n1427), .A(n1428), .S(n1823), .Y(n1426) );
  MUX2X1 U963 ( .B(n1430), .A(n1431), .S(n1811), .Y(n1429) );
  MUX2X1 U964 ( .B(n1433), .A(n1434), .S(n1824), .Y(n1432) );
  MUX2X1 U965 ( .B(n1436), .A(n1437), .S(n1824), .Y(n1435) );
  MUX2X1 U966 ( .B(n1439), .A(n1440), .S(n1824), .Y(n1438) );
  MUX2X1 U967 ( .B(n1442), .A(n1443), .S(n1824), .Y(n1441) );
  MUX2X1 U968 ( .B(n1445), .A(n1446), .S(n1811), .Y(n1444) );
  MUX2X1 U969 ( .B(n1448), .A(n1449), .S(n1824), .Y(n1447) );
  MUX2X1 U970 ( .B(n1451), .A(n1452), .S(n1824), .Y(n1450) );
  MUX2X1 U971 ( .B(n1454), .A(n1455), .S(n1824), .Y(n1453) );
  MUX2X1 U972 ( .B(n1457), .A(n1458), .S(n1824), .Y(n1456) );
  MUX2X1 U973 ( .B(n1460), .A(n1461), .S(n1811), .Y(n1459) );
  MUX2X1 U974 ( .B(n1463), .A(n1464), .S(n1824), .Y(n1462) );
  MUX2X1 U975 ( .B(n1466), .A(n1467), .S(n1824), .Y(n1465) );
  MUX2X1 U976 ( .B(n1469), .A(n1470), .S(n1824), .Y(n1468) );
  MUX2X1 U977 ( .B(n1472), .A(n1473), .S(n1824), .Y(n1471) );
  MUX2X1 U978 ( .B(n1475), .A(n1476), .S(n1811), .Y(n1474) );
  MUX2X1 U979 ( .B(n1478), .A(n1479), .S(n1825), .Y(n1477) );
  MUX2X1 U980 ( .B(n1481), .A(n1482), .S(n1825), .Y(n1480) );
  MUX2X1 U981 ( .B(n1484), .A(n1485), .S(n1825), .Y(n1483) );
  MUX2X1 U982 ( .B(n1487), .A(n1488), .S(n1825), .Y(n1486) );
  MUX2X1 U983 ( .B(n1490), .A(n1491), .S(n1811), .Y(n1489) );
  MUX2X1 U984 ( .B(n1493), .A(n1494), .S(n1825), .Y(n1492) );
  MUX2X1 U985 ( .B(n1496), .A(n1497), .S(n1825), .Y(n1495) );
  MUX2X1 U986 ( .B(n1499), .A(n1500), .S(n1825), .Y(n1498) );
  MUX2X1 U987 ( .B(n1502), .A(n1503), .S(n1825), .Y(n1501) );
  MUX2X1 U988 ( .B(n1505), .A(n1506), .S(n1810), .Y(n1504) );
  MUX2X1 U989 ( .B(n1508), .A(n1509), .S(n1825), .Y(n1507) );
  MUX2X1 U990 ( .B(n1511), .A(n1512), .S(n1825), .Y(n1510) );
  MUX2X1 U991 ( .B(n1514), .A(n1515), .S(n1825), .Y(n1513) );
  MUX2X1 U992 ( .B(n1517), .A(n1518), .S(n1825), .Y(n1516) );
  MUX2X1 U993 ( .B(n1520), .A(n1521), .S(n1810), .Y(n1519) );
  MUX2X1 U994 ( .B(n1523), .A(n1524), .S(n1826), .Y(n1522) );
  MUX2X1 U995 ( .B(n1526), .A(n1527), .S(n1826), .Y(n1525) );
  MUX2X1 U996 ( .B(n1529), .A(n1530), .S(n1826), .Y(n1528) );
  MUX2X1 U997 ( .B(n1532), .A(n1533), .S(n1826), .Y(n1531) );
  MUX2X1 U998 ( .B(n1535), .A(n1536), .S(n1810), .Y(n1534) );
  MUX2X1 U999 ( .B(n1538), .A(n1539), .S(n1826), .Y(n1537) );
  MUX2X1 U1000 ( .B(n1541), .A(n1542), .S(n1826), .Y(n1540) );
  MUX2X1 U1001 ( .B(n1544), .A(n1545), .S(n1826), .Y(n1543) );
  MUX2X1 U1002 ( .B(n1547), .A(n1548), .S(n1826), .Y(n1546) );
  MUX2X1 U1003 ( .B(n1550), .A(n1551), .S(n1810), .Y(n1549) );
  MUX2X1 U1004 ( .B(n1553), .A(n1554), .S(n1826), .Y(n1552) );
  MUX2X1 U1005 ( .B(n1556), .A(n1557), .S(n1826), .Y(n1555) );
  MUX2X1 U1006 ( .B(n1559), .A(n1560), .S(n1826), .Y(n1558) );
  MUX2X1 U1007 ( .B(n1562), .A(n1563), .S(n1826), .Y(n1561) );
  MUX2X1 U1008 ( .B(n1565), .A(n1566), .S(n1810), .Y(n1564) );
  MUX2X1 U1009 ( .B(n1568), .A(n1569), .S(n1827), .Y(n1567) );
  MUX2X1 U1010 ( .B(n1571), .A(n1572), .S(n1827), .Y(n1570) );
  MUX2X1 U1011 ( .B(n1574), .A(n1575), .S(n1827), .Y(n1573) );
  MUX2X1 U1012 ( .B(n1577), .A(n1578), .S(n1827), .Y(n1576) );
  MUX2X1 U1013 ( .B(n1580), .A(n1581), .S(n1810), .Y(n1579) );
  MUX2X1 U1014 ( .B(n1583), .A(n1584), .S(n1827), .Y(n1582) );
  MUX2X1 U1015 ( .B(n1586), .A(n1587), .S(n1827), .Y(n1585) );
  MUX2X1 U1016 ( .B(n1589), .A(n1590), .S(n1827), .Y(n1588) );
  MUX2X1 U1017 ( .B(n1592), .A(n1593), .S(n1827), .Y(n1591) );
  MUX2X1 U1018 ( .B(n1595), .A(n1596), .S(n1810), .Y(n1594) );
  MUX2X1 U1019 ( .B(n1598), .A(n1599), .S(n1827), .Y(n1597) );
  MUX2X1 U1020 ( .B(n1601), .A(n1602), .S(n1827), .Y(n1600) );
  MUX2X1 U1021 ( .B(n1604), .A(n1605), .S(n1827), .Y(n1603) );
  MUX2X1 U1022 ( .B(n1607), .A(n1608), .S(n1827), .Y(n1606) );
  MUX2X1 U1023 ( .B(n1610), .A(n1611), .S(n1810), .Y(n1609) );
  MUX2X1 U1024 ( .B(n1613), .A(n1614), .S(n1828), .Y(n1612) );
  MUX2X1 U1025 ( .B(n1616), .A(n1617), .S(n1828), .Y(n1615) );
  MUX2X1 U1026 ( .B(n1619), .A(n1620), .S(n1828), .Y(n1618) );
  MUX2X1 U1027 ( .B(n1622), .A(n1623), .S(n1828), .Y(n1621) );
  MUX2X1 U1028 ( .B(n1625), .A(n1626), .S(n1810), .Y(n1624) );
  MUX2X1 U1029 ( .B(n1628), .A(n1629), .S(n1828), .Y(n1627) );
  MUX2X1 U1030 ( .B(n1631), .A(n1632), .S(n1828), .Y(n1630) );
  MUX2X1 U1031 ( .B(n1634), .A(n1635), .S(n1828), .Y(n1633) );
  MUX2X1 U1032 ( .B(n1637), .A(n1638), .S(n1828), .Y(n1636) );
  MUX2X1 U1033 ( .B(n1640), .A(n1641), .S(n1810), .Y(n1639) );
  MUX2X1 U1034 ( .B(n1643), .A(n1644), .S(n1828), .Y(n1642) );
  MUX2X1 U1035 ( .B(n1646), .A(n1647), .S(n1828), .Y(n1645) );
  MUX2X1 U1036 ( .B(n1649), .A(n1650), .S(n1828), .Y(n1648) );
  MUX2X1 U1037 ( .B(n1652), .A(n1653), .S(n1828), .Y(n1651) );
  MUX2X1 U1038 ( .B(n1655), .A(n1656), .S(n1810), .Y(n1654) );
  MUX2X1 U1039 ( .B(n1658), .A(n1659), .S(n1829), .Y(n1657) );
  MUX2X1 U1040 ( .B(n1661), .A(n1662), .S(n1829), .Y(n1660) );
  MUX2X1 U1041 ( .B(n1664), .A(n1665), .S(n1829), .Y(n1663) );
  MUX2X1 U1042 ( .B(n1667), .A(n1668), .S(n1829), .Y(n1666) );
  MUX2X1 U1043 ( .B(n1670), .A(n1671), .S(n1810), .Y(n1669) );
  MUX2X1 U1044 ( .B(n1673), .A(n1674), .S(n1829), .Y(n1672) );
  MUX2X1 U1045 ( .B(n1676), .A(n1677), .S(n1829), .Y(n1675) );
  MUX2X1 U1046 ( .B(n1679), .A(n1680), .S(n1829), .Y(n1678) );
  MUX2X1 U1047 ( .B(n1682), .A(n1683), .S(n1829), .Y(n1681) );
  MUX2X1 U1048 ( .B(n1685), .A(n1686), .S(n1809), .Y(n1684) );
  MUX2X1 U1049 ( .B(n1688), .A(n1689), .S(n1829), .Y(n1687) );
  MUX2X1 U1050 ( .B(n1691), .A(n1692), .S(n1829), .Y(n1690) );
  MUX2X1 U1051 ( .B(n1694), .A(n1695), .S(n1829), .Y(n1693) );
  MUX2X1 U1052 ( .B(n1697), .A(n1698), .S(n1829), .Y(n1696) );
  MUX2X1 U1053 ( .B(n1700), .A(n1701), .S(n1809), .Y(n1699) );
  MUX2X1 U1054 ( .B(n1703), .A(n1704), .S(n1830), .Y(n1702) );
  MUX2X1 U1055 ( .B(n1706), .A(n1707), .S(n1830), .Y(n1705) );
  MUX2X1 U1056 ( .B(n1709), .A(n1710), .S(n1830), .Y(n1708) );
  MUX2X1 U1057 ( .B(n1712), .A(n1713), .S(n1830), .Y(n1711) );
  MUX2X1 U1058 ( .B(n1715), .A(n1716), .S(n1809), .Y(n1714) );
  MUX2X1 U1059 ( .B(n1718), .A(n1719), .S(n1830), .Y(n1717) );
  MUX2X1 U1060 ( .B(n1721), .A(n1722), .S(n1830), .Y(n1720) );
  MUX2X1 U1061 ( .B(n1724), .A(n1725), .S(n1830), .Y(n1723) );
  MUX2X1 U1062 ( .B(n1727), .A(n1728), .S(n1830), .Y(n1726) );
  MUX2X1 U1063 ( .B(n1730), .A(n1731), .S(n1809), .Y(n1729) );
  MUX2X1 U1064 ( .B(n1733), .A(n1734), .S(n1830), .Y(n1732) );
  MUX2X1 U1065 ( .B(n1736), .A(n1737), .S(n1830), .Y(n1735) );
  MUX2X1 U1066 ( .B(n1739), .A(n1740), .S(n1830), .Y(n1738) );
  MUX2X1 U1067 ( .B(n1742), .A(n1743), .S(n1830), .Y(n1741) );
  MUX2X1 U1068 ( .B(n1745), .A(n1746), .S(n1809), .Y(n1744) );
  MUX2X1 U1069 ( .B(n1748), .A(n1749), .S(n1831), .Y(n1747) );
  MUX2X1 U1070 ( .B(n1751), .A(n1752), .S(n1831), .Y(n1750) );
  MUX2X1 U1071 ( .B(n1754), .A(n1755), .S(n1831), .Y(n1753) );
  MUX2X1 U1072 ( .B(n1757), .A(n1758), .S(n1831), .Y(n1756) );
  MUX2X1 U1073 ( .B(n1760), .A(n1761), .S(n1809), .Y(n1759) );
  MUX2X1 U1074 ( .B(n1763), .A(n1764), .S(n1831), .Y(n1762) );
  MUX2X1 U1075 ( .B(n1766), .A(n1767), .S(n1831), .Y(n1765) );
  MUX2X1 U1076 ( .B(n1769), .A(n1770), .S(n1831), .Y(n1768) );
  MUX2X1 U1077 ( .B(n1772), .A(n1773), .S(n1831), .Y(n1771) );
  MUX2X1 U1078 ( .B(n1775), .A(n1776), .S(n1809), .Y(n1774) );
  MUX2X1 U1079 ( .B(n1778), .A(n1779), .S(n1831), .Y(n1777) );
  MUX2X1 U1080 ( .B(n1781), .A(n1782), .S(n1831), .Y(n1780) );
  MUX2X1 U1081 ( .B(n1784), .A(n1785), .S(n1831), .Y(n1783) );
  MUX2X1 U1082 ( .B(n1787), .A(n1788), .S(n1831), .Y(n1786) );
  MUX2X1 U1083 ( .B(n1790), .A(n1791), .S(n1809), .Y(n1789) );
  MUX2X1 U1084 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1838), .Y(n1314) );
  MUX2X1 U1085 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1838), .Y(n1313) );
  MUX2X1 U1086 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1838), .Y(n1317) );
  MUX2X1 U1087 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1838), .Y(n1316) );
  MUX2X1 U1088 ( .B(n1315), .A(n1312), .S(n1818), .Y(n1326) );
  MUX2X1 U1089 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1839), .Y(n1320) );
  MUX2X1 U1090 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1839), .Y(n1319) );
  MUX2X1 U1091 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1839), .Y(n1323) );
  MUX2X1 U1092 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1839), .Y(n1322) );
  MUX2X1 U1093 ( .B(n1321), .A(n1318), .S(n1818), .Y(n1325) );
  MUX2X1 U1094 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1839), .Y(n1329) );
  MUX2X1 U1095 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1839), .Y(n1328) );
  MUX2X1 U1096 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1839), .Y(n1332) );
  MUX2X1 U1097 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1839), .Y(n1331) );
  MUX2X1 U1098 ( .B(n1330), .A(n1327), .S(n1818), .Y(n1341) );
  MUX2X1 U1099 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1839), .Y(n1335) );
  MUX2X1 U1100 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1839), .Y(n1334) );
  MUX2X1 U1101 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1839), .Y(n1338) );
  MUX2X1 U1102 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1839), .Y(n1337) );
  MUX2X1 U1103 ( .B(n1336), .A(n1333), .S(n1818), .Y(n1340) );
  MUX2X1 U1104 ( .B(n1339), .A(n1324), .S(n1808), .Y(n1792) );
  MUX2X1 U1105 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1840), .Y(n1344) );
  MUX2X1 U1106 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1840), .Y(n1343) );
  MUX2X1 U1107 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1840), .Y(n1347) );
  MUX2X1 U1108 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1840), .Y(n1346) );
  MUX2X1 U1109 ( .B(n1345), .A(n1342), .S(n1818), .Y(n1356) );
  MUX2X1 U1110 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1840), .Y(n1350) );
  MUX2X1 U1111 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1840), .Y(n1349) );
  MUX2X1 U1112 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1840), .Y(n1353) );
  MUX2X1 U1113 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1840), .Y(n1352) );
  MUX2X1 U1114 ( .B(n1351), .A(n1348), .S(n1818), .Y(n1355) );
  MUX2X1 U1115 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1840), .Y(n1359) );
  MUX2X1 U1116 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1840), .Y(n1358) );
  MUX2X1 U1117 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1840), .Y(n1362) );
  MUX2X1 U1118 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1840), .Y(n1361) );
  MUX2X1 U1119 ( .B(n1360), .A(n1357), .S(n1818), .Y(n1371) );
  MUX2X1 U1120 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1841), .Y(n1365) );
  MUX2X1 U1121 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1841), .Y(n1364) );
  MUX2X1 U1122 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1841), .Y(n1368) );
  MUX2X1 U1123 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1841), .Y(n1367) );
  MUX2X1 U1124 ( .B(n1366), .A(n1363), .S(n1818), .Y(n1370) );
  MUX2X1 U1125 ( .B(n1369), .A(n1354), .S(n1808), .Y(n1793) );
  MUX2X1 U1126 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1841), .Y(n1374) );
  MUX2X1 U1127 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1841), .Y(n1373) );
  MUX2X1 U1128 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1841), .Y(n1377) );
  MUX2X1 U1129 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1841), .Y(n1376) );
  MUX2X1 U1130 ( .B(n1375), .A(n1372), .S(n1818), .Y(n1386) );
  MUX2X1 U1131 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1841), .Y(n1380) );
  MUX2X1 U1132 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1841), .Y(n1379) );
  MUX2X1 U1133 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1841), .Y(n1383) );
  MUX2X1 U1134 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1841), .Y(n1382) );
  MUX2X1 U1135 ( .B(n1381), .A(n1378), .S(n1818), .Y(n1385) );
  MUX2X1 U1136 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1842), .Y(n1389) );
  MUX2X1 U1137 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1842), .Y(n1388) );
  MUX2X1 U1138 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1842), .Y(n1392) );
  MUX2X1 U1139 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1842), .Y(n1391) );
  MUX2X1 U1140 ( .B(n1390), .A(n1387), .S(n1818), .Y(n1401) );
  MUX2X1 U1141 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1842), .Y(n1395) );
  MUX2X1 U1142 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1842), .Y(n1394) );
  MUX2X1 U1143 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1842), .Y(n1398) );
  MUX2X1 U1144 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1842), .Y(n1397) );
  MUX2X1 U1145 ( .B(n1396), .A(n1393), .S(n1818), .Y(n1400) );
  MUX2X1 U1146 ( .B(n1399), .A(n1384), .S(n1808), .Y(n1794) );
  MUX2X1 U1147 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1842), .Y(n1404) );
  MUX2X1 U1148 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1842), .Y(n1403) );
  MUX2X1 U1149 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1842), .Y(n1407) );
  MUX2X1 U1150 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1842), .Y(n1406) );
  MUX2X1 U1151 ( .B(n1405), .A(n1402), .S(n1817), .Y(n1416) );
  MUX2X1 U1152 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1843), .Y(n1410) );
  MUX2X1 U1153 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1843), .Y(n1409) );
  MUX2X1 U1154 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1843), .Y(n1413) );
  MUX2X1 U1155 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1843), .Y(n1412) );
  MUX2X1 U1156 ( .B(n1411), .A(n1408), .S(n1817), .Y(n1415) );
  MUX2X1 U1157 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1843), .Y(n1419) );
  MUX2X1 U1158 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1843), .Y(n1418) );
  MUX2X1 U1159 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1843), .Y(n1422) );
  MUX2X1 U1160 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1843), .Y(n1421) );
  MUX2X1 U1161 ( .B(n1420), .A(n1417), .S(n1817), .Y(n1431) );
  MUX2X1 U1162 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1843), .Y(n1425) );
  MUX2X1 U1163 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1843), .Y(n1424) );
  MUX2X1 U1164 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1843), .Y(n1428) );
  MUX2X1 U1165 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1843), .Y(n1427) );
  MUX2X1 U1166 ( .B(n1426), .A(n1423), .S(n1817), .Y(n1430) );
  MUX2X1 U1167 ( .B(n1429), .A(n1414), .S(n1808), .Y(n1795) );
  MUX2X1 U1168 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1844), .Y(n1434) );
  MUX2X1 U1169 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1844), .Y(n1433) );
  MUX2X1 U1170 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1844), .Y(n1437) );
  MUX2X1 U1171 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1844), .Y(n1436) );
  MUX2X1 U1172 ( .B(n1435), .A(n1432), .S(n1817), .Y(n1446) );
  MUX2X1 U1173 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1844), .Y(n1440) );
  MUX2X1 U1174 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1844), .Y(n1439) );
  MUX2X1 U1175 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1844), .Y(n1443) );
  MUX2X1 U1177 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1844), .Y(n1442) );
  MUX2X1 U1178 ( .B(n1441), .A(n1438), .S(n1817), .Y(n1445) );
  MUX2X1 U1179 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1844), .Y(n1449) );
  MUX2X1 U1180 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1844), .Y(n1448) );
  MUX2X1 U1181 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1844), .Y(n1452) );
  MUX2X1 U1182 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1844), .Y(n1451) );
  MUX2X1 U1183 ( .B(n1450), .A(n1447), .S(n1817), .Y(n1461) );
  MUX2X1 U1184 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1845), .Y(n1455) );
  MUX2X1 U1185 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1845), .Y(n1454) );
  MUX2X1 U1186 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1845), .Y(n1458) );
  MUX2X1 U1187 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1845), .Y(n1457) );
  MUX2X1 U1188 ( .B(n1456), .A(n1453), .S(n1817), .Y(n1460) );
  MUX2X1 U1189 ( .B(n1459), .A(n1444), .S(n1808), .Y(n1796) );
  MUX2X1 U1190 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1845), .Y(n1464) );
  MUX2X1 U1191 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1845), .Y(n1463) );
  MUX2X1 U1192 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1845), .Y(n1467) );
  MUX2X1 U1193 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1845), .Y(n1466) );
  MUX2X1 U1194 ( .B(n1465), .A(n1462), .S(n1817), .Y(n1476) );
  MUX2X1 U1195 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1845), .Y(n1470) );
  MUX2X1 U1196 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1845), .Y(n1469) );
  MUX2X1 U1197 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1845), .Y(n1473) );
  MUX2X1 U1198 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1845), .Y(n1472) );
  MUX2X1 U1199 ( .B(n1471), .A(n1468), .S(n1817), .Y(n1475) );
  MUX2X1 U1200 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1846), .Y(n1479) );
  MUX2X1 U1201 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1846), .Y(n1478) );
  MUX2X1 U1202 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1846), .Y(n1482) );
  MUX2X1 U1203 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1846), .Y(n1481) );
  MUX2X1 U1204 ( .B(n1480), .A(n1477), .S(n1817), .Y(n1491) );
  MUX2X1 U1205 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1846), .Y(n1485) );
  MUX2X1 U1206 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1846), .Y(n1484) );
  MUX2X1 U1207 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1846), .Y(n1488) );
  MUX2X1 U1208 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1846), .Y(n1487) );
  MUX2X1 U1209 ( .B(n1486), .A(n1483), .S(n1817), .Y(n1490) );
  MUX2X1 U1210 ( .B(n1489), .A(n1474), .S(n1808), .Y(n1797) );
  MUX2X1 U1211 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1846), .Y(n1494) );
  MUX2X1 U1212 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1846), .Y(n1493) );
  MUX2X1 U1213 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1846), .Y(n1497) );
  MUX2X1 U1214 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1846), .Y(n1496) );
  MUX2X1 U1215 ( .B(n1495), .A(n1492), .S(n1816), .Y(n1506) );
  MUX2X1 U1216 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1847), .Y(n1500) );
  MUX2X1 U1217 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1847), .Y(n1499) );
  MUX2X1 U1218 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1847), .Y(n1503) );
  MUX2X1 U1219 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1847), .Y(n1502) );
  MUX2X1 U1220 ( .B(n1501), .A(n1498), .S(n1816), .Y(n1505) );
  MUX2X1 U1221 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1847), .Y(n1509) );
  MUX2X1 U1222 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1847), .Y(n1508) );
  MUX2X1 U1223 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1847), .Y(n1512) );
  MUX2X1 U1224 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1847), .Y(n1511) );
  MUX2X1 U1225 ( .B(n1510), .A(n1507), .S(n1816), .Y(n1521) );
  MUX2X1 U1226 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1847), .Y(n1515) );
  MUX2X1 U1227 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1847), .Y(n1514) );
  MUX2X1 U1228 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1847), .Y(n1518) );
  MUX2X1 U1229 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1847), .Y(n1517) );
  MUX2X1 U1230 ( .B(n1516), .A(n1513), .S(n1816), .Y(n1520) );
  MUX2X1 U1231 ( .B(n1519), .A(n1504), .S(n1808), .Y(n1798) );
  MUX2X1 U1232 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1848), .Y(n1524) );
  MUX2X1 U1233 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1848), .Y(n1523) );
  MUX2X1 U1234 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1848), .Y(n1527) );
  MUX2X1 U1235 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1848), .Y(n1526) );
  MUX2X1 U1236 ( .B(n1525), .A(n1522), .S(n1816), .Y(n1536) );
  MUX2X1 U1237 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1848), .Y(n1530) );
  MUX2X1 U1238 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1848), .Y(n1529) );
  MUX2X1 U1239 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1848), .Y(n1533) );
  MUX2X1 U1240 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1848), .Y(n1532) );
  MUX2X1 U1241 ( .B(n1531), .A(n1528), .S(n1816), .Y(n1535) );
  MUX2X1 U1242 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1848), .Y(n1539) );
  MUX2X1 U1243 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1848), .Y(n1538) );
  MUX2X1 U1244 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1848), .Y(n1542) );
  MUX2X1 U1245 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1848), .Y(n1541) );
  MUX2X1 U1246 ( .B(n1540), .A(n1537), .S(n1816), .Y(n1551) );
  MUX2X1 U1247 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1849), .Y(n1545) );
  MUX2X1 U1248 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1849), .Y(n1544) );
  MUX2X1 U1249 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1849), .Y(n1548) );
  MUX2X1 U1250 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1849), .Y(n1547) );
  MUX2X1 U1251 ( .B(n1546), .A(n1543), .S(n1816), .Y(n1550) );
  MUX2X1 U1252 ( .B(n1549), .A(n1534), .S(n1808), .Y(n1799) );
  MUX2X1 U1253 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1849), .Y(n1554) );
  MUX2X1 U1254 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1849), .Y(n1553) );
  MUX2X1 U1255 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1849), .Y(n1557) );
  MUX2X1 U1256 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1849), .Y(n1556) );
  MUX2X1 U1257 ( .B(n1555), .A(n1552), .S(n1816), .Y(n1566) );
  MUX2X1 U1258 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1849), .Y(n1560) );
  MUX2X1 U1259 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1849), .Y(n1559) );
  MUX2X1 U1260 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1849), .Y(n1563) );
  MUX2X1 U1261 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1849), .Y(n1562) );
  MUX2X1 U1262 ( .B(n1561), .A(n1558), .S(n1816), .Y(n1565) );
  MUX2X1 U1263 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1850), .Y(n1569) );
  MUX2X1 U1264 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1850), .Y(n1568) );
  MUX2X1 U1265 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1850), .Y(n1572) );
  MUX2X1 U1266 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1850), .Y(n1571) );
  MUX2X1 U1267 ( .B(n1570), .A(n1567), .S(n1816), .Y(n1581) );
  MUX2X1 U1268 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1850), .Y(n1575) );
  MUX2X1 U1269 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1850), .Y(n1574) );
  MUX2X1 U1270 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1850), .Y(n1578) );
  MUX2X1 U1271 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1850), .Y(n1577) );
  MUX2X1 U1272 ( .B(n1576), .A(n1573), .S(n1816), .Y(n1580) );
  MUX2X1 U1273 ( .B(n1579), .A(n1564), .S(n1808), .Y(n1800) );
  MUX2X1 U1274 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1850), .Y(n1584) );
  MUX2X1 U1275 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1850), .Y(n1583) );
  MUX2X1 U1276 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1850), .Y(n1587) );
  MUX2X1 U1277 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1850), .Y(n1586) );
  MUX2X1 U1278 ( .B(n1585), .A(n1582), .S(n1815), .Y(n1596) );
  MUX2X1 U1279 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1851), .Y(n1590) );
  MUX2X1 U1280 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1851), .Y(n1589) );
  MUX2X1 U1281 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1851), .Y(n1593) );
  MUX2X1 U1282 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1851), .Y(n1592) );
  MUX2X1 U1283 ( .B(n1591), .A(n1588), .S(n1815), .Y(n1595) );
  MUX2X1 U1284 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1851), .Y(n1599) );
  MUX2X1 U1285 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1851), .Y(n1598) );
  MUX2X1 U1286 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1851), .Y(n1602) );
  MUX2X1 U1287 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1851), .Y(n1601) );
  MUX2X1 U1288 ( .B(n1600), .A(n1597), .S(n1815), .Y(n1611) );
  MUX2X1 U1289 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1851), .Y(n1605) );
  MUX2X1 U1290 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1851), .Y(n1604) );
  MUX2X1 U1291 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1851), .Y(n1608) );
  MUX2X1 U1292 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1851), .Y(n1607) );
  MUX2X1 U1293 ( .B(n1606), .A(n1603), .S(n1815), .Y(n1610) );
  MUX2X1 U1294 ( .B(n1609), .A(n1594), .S(n1808), .Y(n1801) );
  MUX2X1 U1295 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1852), .Y(n1614) );
  MUX2X1 U1296 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1852), .Y(n1613) );
  MUX2X1 U1297 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1852), .Y(n1617) );
  MUX2X1 U1298 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1852), .Y(n1616) );
  MUX2X1 U1299 ( .B(n1615), .A(n1612), .S(n1815), .Y(n1626) );
  MUX2X1 U1300 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1852), .Y(n1620) );
  MUX2X1 U1301 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1852), .Y(n1619) );
  MUX2X1 U1302 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1852), .Y(n1623) );
  MUX2X1 U1303 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1852), .Y(n1622) );
  MUX2X1 U1304 ( .B(n1621), .A(n1618), .S(n1815), .Y(n1625) );
  MUX2X1 U1305 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1852), .Y(n1629) );
  MUX2X1 U1306 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1852), .Y(n1628) );
  MUX2X1 U1307 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1852), .Y(n1632) );
  MUX2X1 U1308 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1852), .Y(n1631) );
  MUX2X1 U1309 ( .B(n1630), .A(n1627), .S(n1815), .Y(n1641) );
  MUX2X1 U1310 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1853), .Y(n1635) );
  MUX2X1 U1311 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1853), .Y(n1634) );
  MUX2X1 U1312 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1853), .Y(n1638) );
  MUX2X1 U1313 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1853), .Y(n1637) );
  MUX2X1 U1314 ( .B(n1636), .A(n1633), .S(n1815), .Y(n1640) );
  MUX2X1 U1315 ( .B(n1639), .A(n1624), .S(n1808), .Y(n1802) );
  MUX2X1 U1316 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1853), .Y(n1644) );
  MUX2X1 U1317 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1853), .Y(n1643) );
  MUX2X1 U1318 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1853), .Y(n1647) );
  MUX2X1 U1319 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1853), .Y(n1646) );
  MUX2X1 U1320 ( .B(n1645), .A(n1642), .S(n1815), .Y(n1656) );
  MUX2X1 U1321 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1853), .Y(n1650) );
  MUX2X1 U1322 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1853), .Y(n1649) );
  MUX2X1 U1323 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1853), .Y(n1653) );
  MUX2X1 U1324 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1853), .Y(n1652) );
  MUX2X1 U1325 ( .B(n1651), .A(n1648), .S(n1815), .Y(n1655) );
  MUX2X1 U1326 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1854), .Y(n1659) );
  MUX2X1 U1327 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1854), .Y(n1658) );
  MUX2X1 U1328 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1854), .Y(n1662) );
  MUX2X1 U1329 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1854), .Y(n1661) );
  MUX2X1 U1330 ( .B(n1660), .A(n1657), .S(n1815), .Y(n1671) );
  MUX2X1 U1331 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1854), .Y(n1665) );
  MUX2X1 U1332 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1854), .Y(n1664) );
  MUX2X1 U1333 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1854), .Y(n1668) );
  MUX2X1 U1334 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1854), .Y(n1667) );
  MUX2X1 U1335 ( .B(n1666), .A(n1663), .S(n1815), .Y(n1670) );
  MUX2X1 U1336 ( .B(n1669), .A(n1654), .S(n1808), .Y(n1803) );
  MUX2X1 U1337 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1854), .Y(n1674) );
  MUX2X1 U1338 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1854), .Y(n1673) );
  MUX2X1 U1339 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1854), .Y(n1677) );
  MUX2X1 U1340 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1854), .Y(n1676) );
  MUX2X1 U1341 ( .B(n1675), .A(n1672), .S(n1814), .Y(n1686) );
  MUX2X1 U1342 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1855), .Y(n1680) );
  MUX2X1 U1343 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1855), .Y(n1679) );
  MUX2X1 U1344 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1855), .Y(n1683) );
  MUX2X1 U1345 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1855), .Y(n1682) );
  MUX2X1 U1346 ( .B(n1681), .A(n1678), .S(n1814), .Y(n1685) );
  MUX2X1 U1347 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1855), .Y(n1689) );
  MUX2X1 U1348 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1855), .Y(n1688) );
  MUX2X1 U1349 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1855), .Y(n1692) );
  MUX2X1 U1350 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1855), .Y(n1691) );
  MUX2X1 U1351 ( .B(n1690), .A(n1687), .S(n1814), .Y(n1701) );
  MUX2X1 U1352 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1855), .Y(n1695) );
  MUX2X1 U1353 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1855), .Y(n1694) );
  MUX2X1 U1354 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1855), .Y(n1698) );
  MUX2X1 U1355 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1855), .Y(n1697) );
  MUX2X1 U1356 ( .B(n1696), .A(n1693), .S(n1814), .Y(n1700) );
  MUX2X1 U1357 ( .B(n1699), .A(n1684), .S(n1808), .Y(n1804) );
  MUX2X1 U1358 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1856), .Y(n1704) );
  MUX2X1 U1359 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1856), .Y(n1703) );
  MUX2X1 U1360 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1856), .Y(n1707) );
  MUX2X1 U1361 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1856), .Y(n1706) );
  MUX2X1 U1362 ( .B(n1705), .A(n1702), .S(n1814), .Y(n1716) );
  MUX2X1 U1363 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1856), .Y(n1710) );
  MUX2X1 U1364 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1856), .Y(n1709) );
  MUX2X1 U1365 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1856), .Y(n1713) );
  MUX2X1 U1366 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1856), .Y(n1712) );
  MUX2X1 U1367 ( .B(n1711), .A(n1708), .S(n1814), .Y(n1715) );
  MUX2X1 U1368 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1856), .Y(n1719) );
  MUX2X1 U1369 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1856), .Y(n1718) );
  MUX2X1 U1370 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1856), .Y(n1722) );
  MUX2X1 U1371 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1856), .Y(n1721) );
  MUX2X1 U1372 ( .B(n1720), .A(n1717), .S(n1814), .Y(n1731) );
  MUX2X1 U1373 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1857), .Y(n1725) );
  MUX2X1 U1374 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1857), .Y(n1724) );
  MUX2X1 U1375 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1857), .Y(n1728) );
  MUX2X1 U1376 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1857), .Y(n1727) );
  MUX2X1 U1377 ( .B(n1726), .A(n1723), .S(n1814), .Y(n1730) );
  MUX2X1 U1378 ( .B(n1729), .A(n1714), .S(n1808), .Y(n1805) );
  MUX2X1 U1379 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1857), .Y(n1734) );
  MUX2X1 U1380 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1857), .Y(n1733) );
  MUX2X1 U1381 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1857), .Y(n1737) );
  MUX2X1 U1382 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1857), .Y(n1736) );
  MUX2X1 U1383 ( .B(n1735), .A(n1732), .S(n1814), .Y(n1746) );
  MUX2X1 U1384 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1857), .Y(n1740) );
  MUX2X1 U1385 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1857), .Y(n1739) );
  MUX2X1 U1386 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1857), .Y(n1743) );
  MUX2X1 U1387 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1857), .Y(n1742) );
  MUX2X1 U1388 ( .B(n1741), .A(n1738), .S(n1814), .Y(n1745) );
  MUX2X1 U1389 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1858), .Y(n1749) );
  MUX2X1 U1390 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1858), .Y(n1748) );
  MUX2X1 U1391 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1858), .Y(n1752) );
  MUX2X1 U1392 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1858), .Y(n1751) );
  MUX2X1 U1393 ( .B(n1750), .A(n1747), .S(n1814), .Y(n1761) );
  MUX2X1 U1394 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1858), .Y(n1755) );
  MUX2X1 U1395 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1858), .Y(n1754) );
  MUX2X1 U1396 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1858), .Y(n1758) );
  MUX2X1 U1397 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1858), .Y(n1757) );
  MUX2X1 U1398 ( .B(n1756), .A(n1753), .S(n1814), .Y(n1760) );
  MUX2X1 U1399 ( .B(n1759), .A(n1744), .S(n1808), .Y(n1806) );
  MUX2X1 U1400 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1858), .Y(n1764) );
  MUX2X1 U1401 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1858), .Y(n1763) );
  MUX2X1 U1402 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1858), .Y(n1767) );
  MUX2X1 U1403 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1858), .Y(n1766) );
  MUX2X1 U1404 ( .B(n1765), .A(n1762), .S(n1813), .Y(n1776) );
  MUX2X1 U1405 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1838), .Y(n1770) );
  MUX2X1 U1406 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1858), .Y(n1769) );
  MUX2X1 U1407 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1857), .Y(n1773) );
  MUX2X1 U1408 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1845), .Y(n1772) );
  MUX2X1 U1409 ( .B(n1771), .A(n1768), .S(n1813), .Y(n1775) );
  MUX2X1 U1410 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1839), .Y(n1779) );
  MUX2X1 U1411 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1844), .Y(n1778) );
  MUX2X1 U1412 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1838), .Y(n1782) );
  MUX2X1 U1413 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1857), .Y(n1781) );
  MUX2X1 U1414 ( .B(n1780), .A(n1777), .S(n1813), .Y(n1791) );
  MUX2X1 U1415 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1844), .Y(n1785) );
  MUX2X1 U1416 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1844), .Y(n1784) );
  MUX2X1 U1417 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1838), .Y(n1788) );
  MUX2X1 U1418 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1838), .Y(n1787) );
  MUX2X1 U1419 ( .B(n1786), .A(n1783), .S(n1813), .Y(n1790) );
  MUX2X1 U1420 ( .B(n1789), .A(n1774), .S(n1808), .Y(n1807) );
  INVX8 U1421 ( .A(n1812), .Y(n1814) );
  INVX8 U1422 ( .A(n1812), .Y(n1815) );
  INVX8 U1423 ( .A(n1812), .Y(n1816) );
  INVX8 U1424 ( .A(n1812), .Y(n1817) );
  INVX8 U1425 ( .A(n1812), .Y(n1818) );
  INVX8 U1426 ( .A(n1820), .Y(n1822) );
  INVX8 U1427 ( .A(n1820), .Y(n1823) );
  INVX8 U1428 ( .A(n1820), .Y(n1827) );
  INVX8 U1429 ( .A(n1820), .Y(n1828) );
  INVX8 U1430 ( .A(n1820), .Y(n1830) );
  INVX8 U1431 ( .A(n1820), .Y(n1831) );
  INVX8 U1432 ( .A(n1861), .Y(n1833) );
  INVX8 U1433 ( .A(n1861), .Y(n1834) );
  INVX8 U1434 ( .A(n1861), .Y(n1835) );
  INVX8 U1435 ( .A(n1861), .Y(n1836) );
  INVX8 U1436 ( .A(n1861), .Y(n1837) );
  INVX8 U1437 ( .A(n1837), .Y(n1838) );
  INVX8 U1438 ( .A(n1837), .Y(n1839) );
  INVX8 U1439 ( .A(n1837), .Y(n1840) );
  INVX8 U1440 ( .A(n1836), .Y(n1841) );
  INVX8 U1441 ( .A(n1836), .Y(n1842) );
  INVX8 U1442 ( .A(n1836), .Y(n1843) );
  INVX8 U1443 ( .A(n1837), .Y(n1844) );
  INVX8 U1444 ( .A(n1837), .Y(n1845) );
  INVX8 U1445 ( .A(n1836), .Y(n1846) );
  INVX8 U1446 ( .A(n1835), .Y(n1847) );
  INVX8 U1447 ( .A(n1835), .Y(n1848) );
  INVX8 U1448 ( .A(n1835), .Y(n1849) );
  INVX8 U1449 ( .A(n1834), .Y(n1850) );
  INVX8 U1450 ( .A(n1834), .Y(n1851) );
  INVX8 U1451 ( .A(n1834), .Y(n1852) );
  INVX8 U1452 ( .A(n1833), .Y(n1853) );
  INVX8 U1453 ( .A(n1833), .Y(n1854) );
  INVX8 U1454 ( .A(n1833), .Y(n1855) );
  INVX8 U1455 ( .A(n1832), .Y(n1856) );
  INVX8 U1456 ( .A(n1832), .Y(n1857) );
  INVX8 U1457 ( .A(n1832), .Y(n1858) );
  INVX8 U1458 ( .A(n1859), .Y(n1861) );
  INVX1 U1459 ( .A(N11), .Y(n1961) );
  INVX1 U1460 ( .A(N10), .Y(n1959) );
  INVX8 U1461 ( .A(n1924), .Y(n1921) );
  INVX8 U1462 ( .A(n1924), .Y(n1922) );
  INVX8 U1463 ( .A(n1924), .Y(n1923) );
  INVX8 U1464 ( .A(n623), .Y(n1925) );
  INVX8 U1465 ( .A(n624), .Y(n1927) );
  INVX8 U1466 ( .A(n625), .Y(n1929) );
  INVX8 U1467 ( .A(n626), .Y(n1931) );
  INVX8 U1468 ( .A(n627), .Y(n1933) );
  INVX8 U1469 ( .A(n628), .Y(n1935) );
  INVX8 U1470 ( .A(n629), .Y(n1937) );
  INVX8 U1471 ( .A(n630), .Y(n1939) );
  INVX8 U1472 ( .A(n631), .Y(n1941) );
  INVX8 U1473 ( .A(n632), .Y(n1943) );
  INVX8 U1474 ( .A(n633), .Y(n1945) );
  INVX8 U1475 ( .A(n634), .Y(n1947) );
  INVX8 U1476 ( .A(n635), .Y(n1949) );
  INVX8 U1477 ( .A(n636), .Y(n1951) );
  INVX8 U1478 ( .A(n637), .Y(n1953) );
  INVX8 U1479 ( .A(n638), .Y(n1955) );
  AND2X2 U1480 ( .A(N32), .B(n1233), .Y(\data_out<0> ) );
  AND2X2 U1481 ( .A(N31), .B(n1231), .Y(\data_out<1> ) );
  AND2X2 U1482 ( .A(N30), .B(n1231), .Y(\data_out<2> ) );
  AND2X2 U1483 ( .A(N29), .B(n1234), .Y(\data_out<3> ) );
  AND2X2 U1484 ( .A(N28), .B(n1233), .Y(\data_out<4> ) );
  AND2X2 U1485 ( .A(N27), .B(n1231), .Y(\data_out<5> ) );
  AND2X2 U1486 ( .A(N26), .B(n1233), .Y(\data_out<6> ) );
  AND2X2 U1487 ( .A(N25), .B(n1235), .Y(\data_out<7> ) );
  AND2X2 U1488 ( .A(N24), .B(n1234), .Y(\data_out<8> ) );
  AND2X2 U1489 ( .A(N23), .B(n1235), .Y(\data_out<9> ) );
  AND2X2 U1490 ( .A(N22), .B(n1234), .Y(\data_out<10> ) );
  AND2X2 U1491 ( .A(N21), .B(n1235), .Y(\data_out<11> ) );
  AND2X2 U1492 ( .A(N20), .B(n1231), .Y(\data_out<12> ) );
  AND2X2 U1493 ( .A(N19), .B(n1235), .Y(\data_out<13> ) );
  AND2X2 U1494 ( .A(N18), .B(n1231), .Y(\data_out<14> ) );
  AND2X2 U1495 ( .A(N17), .B(n1233), .Y(\data_out<15> ) );
  OAI21X1 U1496 ( .A(n1863), .B(n1925), .C(n2), .Y(n2700) );
  NAND2X1 U1497 ( .A(\mem<31><1> ), .B(n640), .Y(n1968) );
  OAI21X1 U1498 ( .A(n1928), .B(n1862), .C(n1968), .Y(n2699) );
  NAND2X1 U1499 ( .A(\mem<31><2> ), .B(n640), .Y(n1969) );
  OAI21X1 U1500 ( .A(n1930), .B(n1862), .C(n1969), .Y(n2698) );
  NAND2X1 U1501 ( .A(\mem<31><3> ), .B(n640), .Y(n1970) );
  OAI21X1 U1502 ( .A(n1932), .B(n1862), .C(n1970), .Y(n2697) );
  NAND2X1 U1503 ( .A(\mem<31><4> ), .B(n640), .Y(n1971) );
  OAI21X1 U1504 ( .A(n1934), .B(n1862), .C(n1971), .Y(n2696) );
  NAND2X1 U1505 ( .A(\mem<31><5> ), .B(n640), .Y(n1972) );
  OAI21X1 U1506 ( .A(n1936), .B(n1862), .C(n1972), .Y(n2695) );
  NAND2X1 U1507 ( .A(\mem<31><6> ), .B(n640), .Y(n1973) );
  OAI21X1 U1508 ( .A(n1938), .B(n1862), .C(n1973), .Y(n2694) );
  NAND2X1 U1509 ( .A(\mem<31><7> ), .B(n640), .Y(n1974) );
  OAI21X1 U1510 ( .A(n1940), .B(n1862), .C(n1974), .Y(n2693) );
  NAND2X1 U1511 ( .A(\mem<31><8> ), .B(n640), .Y(n1975) );
  OAI21X1 U1512 ( .A(n1942), .B(n1862), .C(n1975), .Y(n2692) );
  NAND2X1 U1513 ( .A(\mem<31><9> ), .B(n640), .Y(n1976) );
  OAI21X1 U1514 ( .A(n1944), .B(n1863), .C(n1976), .Y(n2691) );
  NAND2X1 U1515 ( .A(\mem<31><10> ), .B(n640), .Y(n1977) );
  OAI21X1 U1516 ( .A(n1946), .B(n1863), .C(n1977), .Y(n2690) );
  NAND2X1 U1517 ( .A(\mem<31><11> ), .B(n640), .Y(n1978) );
  OAI21X1 U1518 ( .A(n1948), .B(n1863), .C(n1978), .Y(n2689) );
  NAND2X1 U1519 ( .A(\mem<31><12> ), .B(n640), .Y(n1979) );
  OAI21X1 U1520 ( .A(n1950), .B(n1863), .C(n1979), .Y(n2688) );
  NAND2X1 U1521 ( .A(\mem<31><13> ), .B(n640), .Y(n1980) );
  OAI21X1 U1522 ( .A(n1952), .B(n1863), .C(n1980), .Y(n2687) );
  NAND2X1 U1523 ( .A(\mem<31><14> ), .B(n640), .Y(n1981) );
  OAI21X1 U1524 ( .A(n1954), .B(n1863), .C(n1981), .Y(n2686) );
  OAI21X1 U1525 ( .A(n1956), .B(n1863), .C(n4), .Y(n2685) );
  OAI21X1 U1526 ( .A(n1864), .B(n1925), .C(n6), .Y(n2684) );
  NAND2X1 U1527 ( .A(\mem<30><1> ), .B(n642), .Y(n1982) );
  OAI21X1 U1528 ( .A(n1864), .B(n1928), .C(n1982), .Y(n2683) );
  NAND2X1 U1529 ( .A(\mem<30><2> ), .B(n642), .Y(n1983) );
  OAI21X1 U1530 ( .A(n1864), .B(n1930), .C(n1983), .Y(n2682) );
  NAND2X1 U1531 ( .A(\mem<30><3> ), .B(n642), .Y(n1984) );
  OAI21X1 U1532 ( .A(n1864), .B(n1932), .C(n1984), .Y(n2681) );
  NAND2X1 U1533 ( .A(\mem<30><4> ), .B(n642), .Y(n1985) );
  OAI21X1 U1534 ( .A(n1864), .B(n1934), .C(n1985), .Y(n2680) );
  NAND2X1 U1535 ( .A(\mem<30><5> ), .B(n642), .Y(n1986) );
  OAI21X1 U1536 ( .A(n1864), .B(n1936), .C(n1986), .Y(n2679) );
  NAND2X1 U1537 ( .A(\mem<30><6> ), .B(n642), .Y(n1987) );
  OAI21X1 U1538 ( .A(n1864), .B(n1938), .C(n1987), .Y(n2678) );
  NAND2X1 U1539 ( .A(\mem<30><7> ), .B(n642), .Y(n1988) );
  OAI21X1 U1540 ( .A(n1864), .B(n1940), .C(n1988), .Y(n2677) );
  NAND2X1 U1541 ( .A(\mem<30><8> ), .B(n642), .Y(n1989) );
  OAI21X1 U1542 ( .A(n1865), .B(n1942), .C(n1989), .Y(n2676) );
  NAND2X1 U1543 ( .A(\mem<30><9> ), .B(n642), .Y(n1990) );
  OAI21X1 U1544 ( .A(n1865), .B(n1944), .C(n1990), .Y(n2675) );
  NAND2X1 U1545 ( .A(\mem<30><10> ), .B(n642), .Y(n1991) );
  OAI21X1 U1546 ( .A(n1865), .B(n1946), .C(n1991), .Y(n2674) );
  NAND2X1 U1547 ( .A(\mem<30><11> ), .B(n642), .Y(n1992) );
  OAI21X1 U1548 ( .A(n1865), .B(n1948), .C(n1992), .Y(n2673) );
  NAND2X1 U1549 ( .A(\mem<30><12> ), .B(n642), .Y(n1993) );
  OAI21X1 U1550 ( .A(n1865), .B(n1950), .C(n1993), .Y(n2672) );
  NAND2X1 U1551 ( .A(\mem<30><13> ), .B(n642), .Y(n1994) );
  OAI21X1 U1552 ( .A(n1865), .B(n1952), .C(n1994), .Y(n2671) );
  NAND2X1 U1553 ( .A(\mem<30><14> ), .B(n642), .Y(n1995) );
  OAI21X1 U1554 ( .A(n1865), .B(n1954), .C(n1995), .Y(n2670) );
  OAI21X1 U1555 ( .A(n1865), .B(n1956), .C(n8), .Y(n2669) );
  NAND3X1 U1556 ( .A(n1958), .B(n1962), .C(n1961), .Y(n1996) );
  NAND2X1 U1557 ( .A(\mem<29><0> ), .B(n645), .Y(n1997) );
  OAI21X1 U1558 ( .A(n1866), .B(n1926), .C(n1997), .Y(n2668) );
  NAND2X1 U1559 ( .A(\mem<29><1> ), .B(n645), .Y(n1998) );
  OAI21X1 U1560 ( .A(n1866), .B(n1928), .C(n1998), .Y(n2667) );
  NAND2X1 U1561 ( .A(\mem<29><2> ), .B(n645), .Y(n1999) );
  OAI21X1 U1562 ( .A(n1866), .B(n1930), .C(n1999), .Y(n2666) );
  NAND2X1 U1563 ( .A(\mem<29><3> ), .B(n645), .Y(n2000) );
  OAI21X1 U1564 ( .A(n1866), .B(n1932), .C(n2000), .Y(n2665) );
  NAND2X1 U1565 ( .A(\mem<29><4> ), .B(n645), .Y(n2001) );
  OAI21X1 U1566 ( .A(n1866), .B(n1934), .C(n2001), .Y(n2664) );
  NAND2X1 U1567 ( .A(\mem<29><5> ), .B(n645), .Y(n2002) );
  OAI21X1 U1568 ( .A(n1866), .B(n1936), .C(n2002), .Y(n2663) );
  NAND2X1 U1569 ( .A(\mem<29><6> ), .B(n645), .Y(n2003) );
  OAI21X1 U1570 ( .A(n1866), .B(n1938), .C(n2003), .Y(n2662) );
  NAND2X1 U1571 ( .A(\mem<29><7> ), .B(n645), .Y(n2004) );
  OAI21X1 U1572 ( .A(n1866), .B(n1940), .C(n2004), .Y(n2661) );
  NAND2X1 U1573 ( .A(\mem<29><8> ), .B(n644), .Y(n2005) );
  OAI21X1 U1574 ( .A(n1867), .B(n1942), .C(n2005), .Y(n2660) );
  NAND2X1 U1575 ( .A(\mem<29><9> ), .B(n644), .Y(n2006) );
  OAI21X1 U1576 ( .A(n1867), .B(n1944), .C(n2006), .Y(n2659) );
  NAND2X1 U1577 ( .A(\mem<29><10> ), .B(n644), .Y(n2007) );
  OAI21X1 U1578 ( .A(n1867), .B(n1946), .C(n2007), .Y(n2658) );
  NAND2X1 U1579 ( .A(\mem<29><11> ), .B(n644), .Y(n2008) );
  OAI21X1 U1580 ( .A(n1867), .B(n1948), .C(n2008), .Y(n2657) );
  NAND2X1 U1581 ( .A(\mem<29><12> ), .B(n644), .Y(n2009) );
  OAI21X1 U1582 ( .A(n1867), .B(n1950), .C(n2009), .Y(n2656) );
  NAND2X1 U1583 ( .A(\mem<29><13> ), .B(n644), .Y(n2010) );
  OAI21X1 U1584 ( .A(n1867), .B(n1952), .C(n2010), .Y(n2655) );
  NAND2X1 U1585 ( .A(\mem<29><14> ), .B(n644), .Y(n2011) );
  OAI21X1 U1586 ( .A(n1867), .B(n1954), .C(n2011), .Y(n2654) );
  OAI21X1 U1587 ( .A(n1867), .B(n1956), .C(n10), .Y(n2653) );
  NAND3X1 U1588 ( .A(n1962), .B(n1961), .C(n1959), .Y(n2012) );
  OAI21X1 U1589 ( .A(n1868), .B(n1925), .C(n12), .Y(n2652) );
  NAND2X1 U1590 ( .A(\mem<28><1> ), .B(n648), .Y(n2013) );
  OAI21X1 U1591 ( .A(n1868), .B(n1928), .C(n2013), .Y(n2651) );
  NAND2X1 U1592 ( .A(\mem<28><2> ), .B(n648), .Y(n2014) );
  OAI21X1 U1593 ( .A(n1868), .B(n1930), .C(n2014), .Y(n2650) );
  NAND2X1 U1594 ( .A(\mem<28><3> ), .B(n648), .Y(n2015) );
  OAI21X1 U1595 ( .A(n1868), .B(n1932), .C(n2015), .Y(n2649) );
  NAND2X1 U1596 ( .A(\mem<28><4> ), .B(n648), .Y(n2016) );
  OAI21X1 U1597 ( .A(n1868), .B(n1934), .C(n2016), .Y(n2648) );
  NAND2X1 U1598 ( .A(\mem<28><5> ), .B(n648), .Y(n2017) );
  OAI21X1 U1599 ( .A(n1868), .B(n1936), .C(n2017), .Y(n2647) );
  NAND2X1 U1600 ( .A(\mem<28><6> ), .B(n648), .Y(n2018) );
  OAI21X1 U1601 ( .A(n1868), .B(n1938), .C(n2018), .Y(n2646) );
  NAND2X1 U1602 ( .A(\mem<28><7> ), .B(n648), .Y(n2019) );
  OAI21X1 U1603 ( .A(n1868), .B(n1940), .C(n2019), .Y(n2645) );
  NAND2X1 U1604 ( .A(\mem<28><8> ), .B(n647), .Y(n2020) );
  OAI21X1 U1605 ( .A(n1869), .B(n1942), .C(n2020), .Y(n2644) );
  NAND2X1 U1606 ( .A(\mem<28><9> ), .B(n647), .Y(n2021) );
  OAI21X1 U1607 ( .A(n1869), .B(n1944), .C(n2021), .Y(n2643) );
  NAND2X1 U1608 ( .A(\mem<28><10> ), .B(n647), .Y(n2022) );
  OAI21X1 U1609 ( .A(n1869), .B(n1946), .C(n2022), .Y(n2642) );
  NAND2X1 U1610 ( .A(\mem<28><11> ), .B(n647), .Y(n2023) );
  OAI21X1 U1611 ( .A(n1869), .B(n1948), .C(n2023), .Y(n2641) );
  NAND2X1 U1612 ( .A(\mem<28><12> ), .B(n647), .Y(n2024) );
  OAI21X1 U1613 ( .A(n1869), .B(n1950), .C(n2024), .Y(n2640) );
  NAND2X1 U1614 ( .A(\mem<28><13> ), .B(n647), .Y(n2025) );
  OAI21X1 U1615 ( .A(n1869), .B(n1952), .C(n2025), .Y(n2639) );
  NAND2X1 U1616 ( .A(\mem<28><14> ), .B(n647), .Y(n2026) );
  OAI21X1 U1617 ( .A(n1869), .B(n1954), .C(n2026), .Y(n2638) );
  OAI21X1 U1618 ( .A(n1869), .B(n1956), .C(n14), .Y(n2637) );
  NAND3X1 U1619 ( .A(n1958), .B(n1960), .C(n1963), .Y(n2027) );
  OAI21X1 U1620 ( .A(n1870), .B(n1925), .C(n16), .Y(n2636) );
  NAND2X1 U1621 ( .A(\mem<27><1> ), .B(n1163), .Y(n2028) );
  OAI21X1 U1622 ( .A(n1870), .B(n1928), .C(n2028), .Y(n2635) );
  NAND2X1 U1623 ( .A(\mem<27><2> ), .B(n1163), .Y(n2029) );
  OAI21X1 U1624 ( .A(n1870), .B(n1930), .C(n2029), .Y(n2634) );
  NAND2X1 U1625 ( .A(\mem<27><3> ), .B(n1163), .Y(n2030) );
  OAI21X1 U1626 ( .A(n1870), .B(n1932), .C(n2030), .Y(n2633) );
  NAND2X1 U1627 ( .A(\mem<27><4> ), .B(n1163), .Y(n2031) );
  OAI21X1 U1628 ( .A(n1870), .B(n1934), .C(n2031), .Y(n2632) );
  NAND2X1 U1629 ( .A(\mem<27><5> ), .B(n1163), .Y(n2032) );
  OAI21X1 U1630 ( .A(n1870), .B(n1936), .C(n2032), .Y(n2631) );
  NAND2X1 U1631 ( .A(\mem<27><6> ), .B(n1163), .Y(n2033) );
  OAI21X1 U1632 ( .A(n1870), .B(n1938), .C(n2033), .Y(n2630) );
  NAND2X1 U1633 ( .A(\mem<27><7> ), .B(n1163), .Y(n2034) );
  OAI21X1 U1634 ( .A(n1870), .B(n1940), .C(n2034), .Y(n2629) );
  NAND2X1 U1635 ( .A(\mem<27><8> ), .B(n650), .Y(n2035) );
  OAI21X1 U1636 ( .A(n1871), .B(n1942), .C(n2035), .Y(n2628) );
  NAND2X1 U1637 ( .A(\mem<27><9> ), .B(n650), .Y(n2036) );
  OAI21X1 U1638 ( .A(n1871), .B(n1944), .C(n2036), .Y(n2627) );
  NAND2X1 U1639 ( .A(\mem<27><10> ), .B(n650), .Y(n2037) );
  OAI21X1 U1640 ( .A(n1871), .B(n1946), .C(n2037), .Y(n2626) );
  NAND2X1 U1641 ( .A(\mem<27><11> ), .B(n650), .Y(n2038) );
  OAI21X1 U1642 ( .A(n1871), .B(n1948), .C(n2038), .Y(n2625) );
  NAND2X1 U1643 ( .A(\mem<27><12> ), .B(n650), .Y(n2039) );
  OAI21X1 U1644 ( .A(n1871), .B(n1950), .C(n2039), .Y(n2624) );
  NAND2X1 U1645 ( .A(\mem<27><13> ), .B(n650), .Y(n2040) );
  OAI21X1 U1646 ( .A(n1871), .B(n1952), .C(n2040), .Y(n2623) );
  NAND2X1 U1647 ( .A(\mem<27><14> ), .B(n650), .Y(n2041) );
  OAI21X1 U1648 ( .A(n1871), .B(n1954), .C(n2041), .Y(n2622) );
  OAI21X1 U1649 ( .A(n1871), .B(n1956), .C(n18), .Y(n2621) );
  NAND3X1 U1650 ( .A(n1963), .B(n1960), .C(n1959), .Y(n2042) );
  NAND2X1 U1651 ( .A(\mem<26><0> ), .B(n1166), .Y(n2043) );
  OAI21X1 U1652 ( .A(n1872), .B(n1926), .C(n2043), .Y(n2620) );
  NAND2X1 U1653 ( .A(\mem<26><1> ), .B(n1166), .Y(n2044) );
  OAI21X1 U1654 ( .A(n1872), .B(n1928), .C(n2044), .Y(n2619) );
  NAND2X1 U1655 ( .A(\mem<26><2> ), .B(n1166), .Y(n2045) );
  OAI21X1 U1656 ( .A(n1872), .B(n1930), .C(n2045), .Y(n2618) );
  NAND2X1 U1657 ( .A(\mem<26><3> ), .B(n1166), .Y(n2046) );
  OAI21X1 U1658 ( .A(n1872), .B(n1932), .C(n2046), .Y(n2617) );
  NAND2X1 U1659 ( .A(\mem<26><4> ), .B(n1166), .Y(n2047) );
  OAI21X1 U1660 ( .A(n1872), .B(n1934), .C(n2047), .Y(n2616) );
  NAND2X1 U1661 ( .A(\mem<26><5> ), .B(n1166), .Y(n2048) );
  OAI21X1 U1662 ( .A(n1872), .B(n1936), .C(n2048), .Y(n2615) );
  NAND2X1 U1663 ( .A(\mem<26><6> ), .B(n1166), .Y(n2049) );
  OAI21X1 U1664 ( .A(n1872), .B(n1938), .C(n2049), .Y(n2614) );
  NAND2X1 U1665 ( .A(\mem<26><7> ), .B(n1166), .Y(n2050) );
  OAI21X1 U1666 ( .A(n1872), .B(n1940), .C(n2050), .Y(n2613) );
  NAND2X1 U1667 ( .A(\mem<26><8> ), .B(n1165), .Y(n2051) );
  OAI21X1 U1668 ( .A(n1873), .B(n1942), .C(n2051), .Y(n2612) );
  NAND2X1 U1669 ( .A(\mem<26><9> ), .B(n1165), .Y(n2052) );
  OAI21X1 U1670 ( .A(n1873), .B(n1944), .C(n2052), .Y(n2611) );
  NAND2X1 U1671 ( .A(\mem<26><10> ), .B(n1165), .Y(n2053) );
  OAI21X1 U1672 ( .A(n1873), .B(n1946), .C(n2053), .Y(n2610) );
  NAND2X1 U1673 ( .A(\mem<26><11> ), .B(n1165), .Y(n2054) );
  OAI21X1 U1674 ( .A(n1873), .B(n1948), .C(n2054), .Y(n2609) );
  NAND2X1 U1675 ( .A(\mem<26><12> ), .B(n1165), .Y(n2055) );
  OAI21X1 U1676 ( .A(n1873), .B(n1950), .C(n2055), .Y(n2608) );
  NAND2X1 U1677 ( .A(\mem<26><13> ), .B(n1165), .Y(n2056) );
  OAI21X1 U1678 ( .A(n1873), .B(n1952), .C(n2056), .Y(n2607) );
  NAND2X1 U1679 ( .A(\mem<26><14> ), .B(n1165), .Y(n2057) );
  OAI21X1 U1680 ( .A(n1873), .B(n1954), .C(n2057), .Y(n2606) );
  OAI21X1 U1681 ( .A(n1873), .B(n1956), .C(n20), .Y(n2605) );
  NAND3X1 U1682 ( .A(n1958), .B(n1963), .C(n1961), .Y(n2058) );
  OAI21X1 U1683 ( .A(n1874), .B(n1925), .C(n22), .Y(n2604) );
  NAND2X1 U1684 ( .A(\mem<25><1> ), .B(n1169), .Y(n2059) );
  OAI21X1 U1685 ( .A(n1874), .B(n1928), .C(n2059), .Y(n2603) );
  NAND2X1 U1686 ( .A(\mem<25><2> ), .B(n1169), .Y(n2060) );
  OAI21X1 U1687 ( .A(n1874), .B(n1930), .C(n2060), .Y(n2602) );
  NAND2X1 U1688 ( .A(\mem<25><3> ), .B(n1169), .Y(n2061) );
  OAI21X1 U1689 ( .A(n1874), .B(n1932), .C(n2061), .Y(n2601) );
  NAND2X1 U1690 ( .A(\mem<25><4> ), .B(n1169), .Y(n2062) );
  OAI21X1 U1691 ( .A(n1874), .B(n1934), .C(n2062), .Y(n2600) );
  NAND2X1 U1692 ( .A(\mem<25><5> ), .B(n1169), .Y(n2063) );
  OAI21X1 U1693 ( .A(n1874), .B(n1936), .C(n2063), .Y(n2599) );
  NAND2X1 U1694 ( .A(\mem<25><6> ), .B(n1169), .Y(n2064) );
  OAI21X1 U1695 ( .A(n1874), .B(n1938), .C(n2064), .Y(n2598) );
  NAND2X1 U1696 ( .A(\mem<25><7> ), .B(n1169), .Y(n2065) );
  OAI21X1 U1697 ( .A(n1874), .B(n1940), .C(n2065), .Y(n2597) );
  NAND2X1 U1698 ( .A(\mem<25><8> ), .B(n1168), .Y(n2066) );
  OAI21X1 U1699 ( .A(n1875), .B(n1942), .C(n2066), .Y(n2596) );
  NAND2X1 U1700 ( .A(\mem<25><9> ), .B(n1168), .Y(n2067) );
  OAI21X1 U1701 ( .A(n1875), .B(n1944), .C(n2067), .Y(n2595) );
  NAND2X1 U1702 ( .A(\mem<25><10> ), .B(n1168), .Y(n2068) );
  OAI21X1 U1703 ( .A(n1875), .B(n1946), .C(n2068), .Y(n2594) );
  NAND2X1 U1704 ( .A(\mem<25><11> ), .B(n1168), .Y(n2069) );
  OAI21X1 U1705 ( .A(n1875), .B(n1948), .C(n2069), .Y(n2593) );
  NAND2X1 U1706 ( .A(\mem<25><12> ), .B(n1168), .Y(n2070) );
  OAI21X1 U1707 ( .A(n1875), .B(n1950), .C(n2070), .Y(n2592) );
  NAND2X1 U1708 ( .A(\mem<25><13> ), .B(n1168), .Y(n2071) );
  OAI21X1 U1709 ( .A(n1875), .B(n1952), .C(n2071), .Y(n2591) );
  NAND2X1 U1710 ( .A(\mem<25><14> ), .B(n1168), .Y(n2072) );
  OAI21X1 U1711 ( .A(n1875), .B(n1954), .C(n2072), .Y(n2590) );
  OAI21X1 U1712 ( .A(n1875), .B(n1956), .C(n24), .Y(n2589) );
  NOR3X1 U1713 ( .A(n1958), .B(n1960), .C(n1962), .Y(n2172) );
  OAI21X1 U1714 ( .A(n1250), .B(n1925), .C(n26), .Y(n2588) );
  NAND2X1 U1715 ( .A(\mem<24><1> ), .B(n1172), .Y(n2073) );
  OAI21X1 U1716 ( .A(n1250), .B(n1928), .C(n2073), .Y(n2587) );
  NAND2X1 U1717 ( .A(\mem<24><2> ), .B(n1172), .Y(n2074) );
  OAI21X1 U1718 ( .A(n1250), .B(n1930), .C(n2074), .Y(n2586) );
  NAND2X1 U1719 ( .A(\mem<24><3> ), .B(n1172), .Y(n2075) );
  OAI21X1 U1720 ( .A(n1250), .B(n1932), .C(n2075), .Y(n2585) );
  NAND2X1 U1721 ( .A(\mem<24><4> ), .B(n1172), .Y(n2076) );
  OAI21X1 U1722 ( .A(n1250), .B(n1934), .C(n2076), .Y(n2584) );
  NAND2X1 U1723 ( .A(\mem<24><5> ), .B(n1172), .Y(n2077) );
  OAI21X1 U1724 ( .A(n1250), .B(n1936), .C(n2077), .Y(n2583) );
  NAND2X1 U1725 ( .A(\mem<24><6> ), .B(n1172), .Y(n2078) );
  OAI21X1 U1726 ( .A(n1250), .B(n1938), .C(n2078), .Y(n2582) );
  NAND2X1 U1727 ( .A(\mem<24><7> ), .B(n1172), .Y(n2079) );
  OAI21X1 U1728 ( .A(n1250), .B(n1940), .C(n2079), .Y(n2581) );
  NAND2X1 U1729 ( .A(\mem<24><8> ), .B(n1171), .Y(n2080) );
  OAI21X1 U1730 ( .A(n1250), .B(n1942), .C(n2080), .Y(n2580) );
  NAND2X1 U1731 ( .A(\mem<24><9> ), .B(n1171), .Y(n2081) );
  OAI21X1 U1732 ( .A(n1250), .B(n1944), .C(n2081), .Y(n2579) );
  NAND2X1 U1733 ( .A(\mem<24><10> ), .B(n1171), .Y(n2082) );
  OAI21X1 U1734 ( .A(n1250), .B(n1946), .C(n2082), .Y(n2578) );
  NAND2X1 U1735 ( .A(\mem<24><11> ), .B(n1171), .Y(n2083) );
  OAI21X1 U1736 ( .A(n1250), .B(n1948), .C(n2083), .Y(n2577) );
  NAND2X1 U1737 ( .A(\mem<24><12> ), .B(n1171), .Y(n2084) );
  OAI21X1 U1738 ( .A(n1250), .B(n1950), .C(n2084), .Y(n2576) );
  NAND2X1 U1739 ( .A(\mem<24><13> ), .B(n1171), .Y(n2085) );
  OAI21X1 U1740 ( .A(n1250), .B(n1952), .C(n2085), .Y(n2575) );
  NAND2X1 U1741 ( .A(\mem<24><14> ), .B(n1171), .Y(n2086) );
  OAI21X1 U1742 ( .A(n1250), .B(n1954), .C(n2086), .Y(n2574) );
  OAI21X1 U1743 ( .A(n1250), .B(n1956), .C(n28), .Y(n2573) );
  OAI21X1 U1744 ( .A(n1876), .B(n1925), .C(n30), .Y(n2572) );
  OAI21X1 U1745 ( .A(n1876), .B(n1927), .C(n32), .Y(n2571) );
  OAI21X1 U1746 ( .A(n1876), .B(n1929), .C(n34), .Y(n2570) );
  OAI21X1 U1747 ( .A(n1876), .B(n1931), .C(n36), .Y(n2569) );
  OAI21X1 U1748 ( .A(n1876), .B(n1933), .C(n38), .Y(n2568) );
  OAI21X1 U1749 ( .A(n1876), .B(n1935), .C(n40), .Y(n2567) );
  OAI21X1 U1750 ( .A(n1876), .B(n1937), .C(n42), .Y(n2566) );
  OAI21X1 U1751 ( .A(n1876), .B(n1939), .C(n44), .Y(n2565) );
  OAI21X1 U1752 ( .A(n1877), .B(n1941), .C(n46), .Y(n2564) );
  OAI21X1 U1753 ( .A(n1877), .B(n1943), .C(n48), .Y(n2563) );
  OAI21X1 U1754 ( .A(n1877), .B(n1945), .C(n50), .Y(n2562) );
  OAI21X1 U1755 ( .A(n1877), .B(n1947), .C(n52), .Y(n2561) );
  OAI21X1 U1756 ( .A(n1877), .B(n1949), .C(n54), .Y(n2560) );
  OAI21X1 U1757 ( .A(n1877), .B(n1951), .C(n56), .Y(n2559) );
  OAI21X1 U1758 ( .A(n1877), .B(n1953), .C(n58), .Y(n2558) );
  OAI21X1 U1759 ( .A(n1877), .B(n1955), .C(n60), .Y(n2557) );
  OAI21X1 U1760 ( .A(n1878), .B(n1925), .C(n62), .Y(n2556) );
  OAI21X1 U1761 ( .A(n1878), .B(n1927), .C(n64), .Y(n2555) );
  OAI21X1 U1762 ( .A(n1878), .B(n1929), .C(n66), .Y(n2554) );
  OAI21X1 U1763 ( .A(n1878), .B(n1931), .C(n68), .Y(n2553) );
  OAI21X1 U1764 ( .A(n1878), .B(n1933), .C(n70), .Y(n2552) );
  OAI21X1 U1765 ( .A(n1878), .B(n1935), .C(n72), .Y(n2551) );
  OAI21X1 U1766 ( .A(n1878), .B(n1937), .C(n74), .Y(n2550) );
  OAI21X1 U1767 ( .A(n1878), .B(n1939), .C(n76), .Y(n2549) );
  OAI21X1 U1768 ( .A(n1879), .B(n1941), .C(n78), .Y(n2548) );
  OAI21X1 U1769 ( .A(n1879), .B(n1943), .C(n80), .Y(n2547) );
  OAI21X1 U1770 ( .A(n1879), .B(n1945), .C(n82), .Y(n2546) );
  OAI21X1 U1771 ( .A(n1879), .B(n1947), .C(n84), .Y(n2545) );
  OAI21X1 U1772 ( .A(n1879), .B(n1949), .C(n86), .Y(n2544) );
  OAI21X1 U1773 ( .A(n1879), .B(n1951), .C(n88), .Y(n2543) );
  OAI21X1 U1774 ( .A(n1879), .B(n1953), .C(n90), .Y(n2542) );
  OAI21X1 U1775 ( .A(n1879), .B(n1955), .C(n92), .Y(n2541) );
  OAI21X1 U1776 ( .A(n1880), .B(n1925), .C(n94), .Y(n2540) );
  OAI21X1 U1777 ( .A(n1880), .B(n1927), .C(n96), .Y(n2539) );
  OAI21X1 U1778 ( .A(n1880), .B(n1929), .C(n98), .Y(n2538) );
  OAI21X1 U1779 ( .A(n1880), .B(n1931), .C(n100), .Y(n2537) );
  OAI21X1 U1780 ( .A(n1880), .B(n1933), .C(n102), .Y(n2536) );
  OAI21X1 U1781 ( .A(n1880), .B(n1935), .C(n104), .Y(n2535) );
  OAI21X1 U1782 ( .A(n1880), .B(n1937), .C(n106), .Y(n2534) );
  OAI21X1 U1783 ( .A(n1880), .B(n1939), .C(n108), .Y(n2533) );
  OAI21X1 U1784 ( .A(n1881), .B(n1941), .C(n110), .Y(n2532) );
  OAI21X1 U1785 ( .A(n1881), .B(n1943), .C(n112), .Y(n2531) );
  OAI21X1 U1786 ( .A(n1881), .B(n1945), .C(n114), .Y(n2530) );
  OAI21X1 U1787 ( .A(n1881), .B(n1947), .C(n116), .Y(n2529) );
  OAI21X1 U1788 ( .A(n1881), .B(n1949), .C(n118), .Y(n2528) );
  OAI21X1 U1789 ( .A(n1881), .B(n1951), .C(n120), .Y(n2527) );
  OAI21X1 U1790 ( .A(n1881), .B(n1953), .C(n122), .Y(n2526) );
  OAI21X1 U1791 ( .A(n1881), .B(n1955), .C(n124), .Y(n2525) );
  NAND2X1 U1792 ( .A(\mem<20><0> ), .B(n615), .Y(n2087) );
  OAI21X1 U1793 ( .A(n1882), .B(n1925), .C(n2087), .Y(n2524) );
  NAND2X1 U1794 ( .A(\mem<20><1> ), .B(n615), .Y(n2088) );
  OAI21X1 U1795 ( .A(n1882), .B(n1927), .C(n2088), .Y(n2523) );
  NAND2X1 U1796 ( .A(\mem<20><2> ), .B(n615), .Y(n2089) );
  OAI21X1 U1797 ( .A(n1882), .B(n1929), .C(n2089), .Y(n2522) );
  NAND2X1 U1798 ( .A(\mem<20><3> ), .B(n615), .Y(n2090) );
  OAI21X1 U1799 ( .A(n1882), .B(n1931), .C(n2090), .Y(n2521) );
  NAND2X1 U1800 ( .A(\mem<20><4> ), .B(n615), .Y(n2091) );
  OAI21X1 U1801 ( .A(n1882), .B(n1933), .C(n2091), .Y(n2520) );
  NAND2X1 U1802 ( .A(\mem<20><5> ), .B(n615), .Y(n2092) );
  OAI21X1 U1803 ( .A(n1882), .B(n1935), .C(n2092), .Y(n2519) );
  NAND2X1 U1804 ( .A(\mem<20><6> ), .B(n615), .Y(n2093) );
  OAI21X1 U1805 ( .A(n1882), .B(n1937), .C(n2093), .Y(n2518) );
  NAND2X1 U1806 ( .A(\mem<20><7> ), .B(n615), .Y(n2094) );
  OAI21X1 U1807 ( .A(n1882), .B(n1939), .C(n2094), .Y(n2517) );
  NAND2X1 U1808 ( .A(\mem<20><8> ), .B(n615), .Y(n2095) );
  OAI21X1 U1809 ( .A(n1883), .B(n1941), .C(n2095), .Y(n2516) );
  NAND2X1 U1810 ( .A(\mem<20><9> ), .B(n615), .Y(n2096) );
  OAI21X1 U1811 ( .A(n1883), .B(n1943), .C(n2096), .Y(n2515) );
  NAND2X1 U1812 ( .A(\mem<20><10> ), .B(n615), .Y(n2097) );
  OAI21X1 U1813 ( .A(n1883), .B(n1945), .C(n2097), .Y(n2514) );
  NAND2X1 U1814 ( .A(\mem<20><11> ), .B(n615), .Y(n2098) );
  OAI21X1 U1815 ( .A(n1883), .B(n1947), .C(n2098), .Y(n2513) );
  NAND2X1 U1816 ( .A(\mem<20><12> ), .B(n615), .Y(n2099) );
  OAI21X1 U1817 ( .A(n1883), .B(n1949), .C(n2099), .Y(n2512) );
  NAND2X1 U1818 ( .A(\mem<20><13> ), .B(n615), .Y(n2100) );
  OAI21X1 U1819 ( .A(n1883), .B(n1951), .C(n2100), .Y(n2511) );
  NAND2X1 U1820 ( .A(\mem<20><14> ), .B(n615), .Y(n2101) );
  OAI21X1 U1821 ( .A(n1883), .B(n1953), .C(n2101), .Y(n2510) );
  NAND2X1 U1822 ( .A(\mem<20><15> ), .B(n615), .Y(n2102) );
  OAI21X1 U1823 ( .A(n1883), .B(n1955), .C(n2102), .Y(n2509) );
  NAND2X1 U1824 ( .A(\mem<19><0> ), .B(n617), .Y(n2103) );
  OAI21X1 U1825 ( .A(n1884), .B(n1925), .C(n2103), .Y(n2508) );
  NAND2X1 U1826 ( .A(\mem<19><1> ), .B(n617), .Y(n2104) );
  OAI21X1 U1827 ( .A(n1884), .B(n1927), .C(n2104), .Y(n2507) );
  NAND2X1 U1828 ( .A(\mem<19><2> ), .B(n617), .Y(n2105) );
  OAI21X1 U1829 ( .A(n1884), .B(n1929), .C(n2105), .Y(n2506) );
  NAND2X1 U1830 ( .A(\mem<19><3> ), .B(n617), .Y(n2106) );
  OAI21X1 U1831 ( .A(n1884), .B(n1931), .C(n2106), .Y(n2505) );
  NAND2X1 U1832 ( .A(\mem<19><4> ), .B(n617), .Y(n2107) );
  OAI21X1 U1833 ( .A(n1884), .B(n1933), .C(n2107), .Y(n2504) );
  NAND2X1 U1834 ( .A(\mem<19><5> ), .B(n617), .Y(n2108) );
  OAI21X1 U1835 ( .A(n1884), .B(n1935), .C(n2108), .Y(n2503) );
  NAND2X1 U1836 ( .A(\mem<19><6> ), .B(n617), .Y(n2109) );
  OAI21X1 U1837 ( .A(n1884), .B(n1937), .C(n2109), .Y(n2502) );
  NAND2X1 U1838 ( .A(\mem<19><7> ), .B(n617), .Y(n2110) );
  OAI21X1 U1839 ( .A(n1884), .B(n1939), .C(n2110), .Y(n2501) );
  NAND2X1 U1840 ( .A(\mem<19><8> ), .B(n617), .Y(n2111) );
  OAI21X1 U1841 ( .A(n1885), .B(n1941), .C(n2111), .Y(n2500) );
  NAND2X1 U1842 ( .A(\mem<19><9> ), .B(n617), .Y(n2112) );
  OAI21X1 U1843 ( .A(n1885), .B(n1943), .C(n2112), .Y(n2499) );
  NAND2X1 U1844 ( .A(\mem<19><10> ), .B(n617), .Y(n2113) );
  OAI21X1 U1845 ( .A(n1885), .B(n1945), .C(n2113), .Y(n2498) );
  NAND2X1 U1846 ( .A(\mem<19><11> ), .B(n617), .Y(n2114) );
  OAI21X1 U1847 ( .A(n1885), .B(n1947), .C(n2114), .Y(n2497) );
  NAND2X1 U1848 ( .A(\mem<19><12> ), .B(n617), .Y(n2115) );
  OAI21X1 U1849 ( .A(n1885), .B(n1949), .C(n2115), .Y(n2496) );
  NAND2X1 U1850 ( .A(\mem<19><13> ), .B(n617), .Y(n2116) );
  OAI21X1 U1851 ( .A(n1885), .B(n1951), .C(n2116), .Y(n2495) );
  NAND2X1 U1852 ( .A(\mem<19><14> ), .B(n617), .Y(n2117) );
  OAI21X1 U1853 ( .A(n1885), .B(n1953), .C(n2117), .Y(n2494) );
  NAND2X1 U1854 ( .A(\mem<19><15> ), .B(n617), .Y(n2118) );
  OAI21X1 U1855 ( .A(n1885), .B(n1955), .C(n2118), .Y(n2493) );
  OAI21X1 U1856 ( .A(n1886), .B(n1925), .C(n126), .Y(n2492) );
  OAI21X1 U1857 ( .A(n1886), .B(n1927), .C(n128), .Y(n2491) );
  OAI21X1 U1858 ( .A(n1886), .B(n1929), .C(n130), .Y(n2490) );
  OAI21X1 U1859 ( .A(n1886), .B(n1931), .C(n132), .Y(n2489) );
  OAI21X1 U1860 ( .A(n1886), .B(n1933), .C(n134), .Y(n2488) );
  OAI21X1 U1861 ( .A(n1886), .B(n1935), .C(n136), .Y(n2487) );
  OAI21X1 U1862 ( .A(n1886), .B(n1937), .C(n138), .Y(n2486) );
  OAI21X1 U1863 ( .A(n1886), .B(n1939), .C(n140), .Y(n2485) );
  OAI21X1 U1864 ( .A(n1887), .B(n1941), .C(n142), .Y(n2484) );
  OAI21X1 U1865 ( .A(n1887), .B(n1943), .C(n144), .Y(n2483) );
  OAI21X1 U1866 ( .A(n1887), .B(n1945), .C(n146), .Y(n2482) );
  OAI21X1 U1867 ( .A(n1887), .B(n1947), .C(n148), .Y(n2481) );
  OAI21X1 U1868 ( .A(n1887), .B(n1949), .C(n150), .Y(n2480) );
  OAI21X1 U1869 ( .A(n1887), .B(n1951), .C(n152), .Y(n2479) );
  OAI21X1 U1870 ( .A(n1887), .B(n1953), .C(n154), .Y(n2478) );
  OAI21X1 U1871 ( .A(n1887), .B(n1955), .C(n156), .Y(n2477) );
  OAI21X1 U1872 ( .A(n1888), .B(n1925), .C(n158), .Y(n2476) );
  OAI21X1 U1873 ( .A(n1888), .B(n1927), .C(n160), .Y(n2475) );
  OAI21X1 U1874 ( .A(n1888), .B(n1929), .C(n162), .Y(n2474) );
  OAI21X1 U1875 ( .A(n1888), .B(n1931), .C(n164), .Y(n2473) );
  OAI21X1 U1876 ( .A(n1888), .B(n1933), .C(n166), .Y(n2472) );
  OAI21X1 U1877 ( .A(n1888), .B(n1935), .C(n168), .Y(n2471) );
  OAI21X1 U1878 ( .A(n1888), .B(n1937), .C(n170), .Y(n2470) );
  OAI21X1 U1879 ( .A(n1888), .B(n1939), .C(n172), .Y(n2469) );
  OAI21X1 U1880 ( .A(n1889), .B(n1941), .C(n174), .Y(n2468) );
  OAI21X1 U1881 ( .A(n1889), .B(n1943), .C(n176), .Y(n2467) );
  OAI21X1 U1882 ( .A(n1889), .B(n1945), .C(n178), .Y(n2466) );
  OAI21X1 U1883 ( .A(n1889), .B(n1947), .C(n180), .Y(n2465) );
  OAI21X1 U1884 ( .A(n1889), .B(n1949), .C(n182), .Y(n2464) );
  OAI21X1 U1885 ( .A(n1889), .B(n1951), .C(n184), .Y(n2463) );
  OAI21X1 U1886 ( .A(n1889), .B(n1953), .C(n186), .Y(n2462) );
  OAI21X1 U1887 ( .A(n1889), .B(n1955), .C(n188), .Y(n2461) );
  OAI21X1 U1888 ( .A(n1890), .B(n1925), .C(n190), .Y(n2460) );
  OAI21X1 U1889 ( .A(n1890), .B(n1927), .C(n192), .Y(n2459) );
  OAI21X1 U1890 ( .A(n1890), .B(n1929), .C(n194), .Y(n2458) );
  OAI21X1 U1891 ( .A(n1890), .B(n1931), .C(n196), .Y(n2457) );
  OAI21X1 U1892 ( .A(n1890), .B(n1933), .C(n198), .Y(n2456) );
  OAI21X1 U1893 ( .A(n1890), .B(n1935), .C(n200), .Y(n2455) );
  OAI21X1 U1894 ( .A(n1890), .B(n1937), .C(n202), .Y(n2454) );
  OAI21X1 U1895 ( .A(n1890), .B(n1939), .C(n204), .Y(n2453) );
  OAI21X1 U1896 ( .A(n1890), .B(n1941), .C(n206), .Y(n2452) );
  OAI21X1 U1897 ( .A(n1890), .B(n1943), .C(n208), .Y(n2451) );
  OAI21X1 U1898 ( .A(n1890), .B(n1945), .C(n210), .Y(n2450) );
  OAI21X1 U1899 ( .A(n1890), .B(n1947), .C(n212), .Y(n2449) );
  OAI21X1 U1900 ( .A(n1890), .B(n1949), .C(n215), .Y(n2448) );
  OAI21X1 U1901 ( .A(n1890), .B(n1951), .C(n217), .Y(n2447) );
  OAI21X1 U1902 ( .A(n1890), .B(n1953), .C(n219), .Y(n2446) );
  OAI21X1 U1903 ( .A(n1890), .B(n1955), .C(n221), .Y(n2445) );
  NAND3X1 U1904 ( .A(n1964), .B(n2701), .C(n1967), .Y(n2119) );
  OAI21X1 U1905 ( .A(n1891), .B(n1925), .C(n223), .Y(n2444) );
  OAI21X1 U1906 ( .A(n1891), .B(n1927), .C(n225), .Y(n2443) );
  OAI21X1 U1907 ( .A(n1891), .B(n1929), .C(n227), .Y(n2442) );
  OAI21X1 U1908 ( .A(n1891), .B(n1931), .C(n229), .Y(n2441) );
  OAI21X1 U1909 ( .A(n1891), .B(n1933), .C(n231), .Y(n2440) );
  OAI21X1 U1910 ( .A(n1891), .B(n1935), .C(n233), .Y(n2439) );
  OAI21X1 U1911 ( .A(n1891), .B(n1937), .C(n235), .Y(n2438) );
  OAI21X1 U1912 ( .A(n1891), .B(n1939), .C(n237), .Y(n2437) );
  OAI21X1 U1913 ( .A(n1892), .B(n1941), .C(n239), .Y(n2436) );
  OAI21X1 U1914 ( .A(n1892), .B(n1943), .C(n241), .Y(n2435) );
  OAI21X1 U1915 ( .A(n1892), .B(n1945), .C(n243), .Y(n2434) );
  OAI21X1 U1916 ( .A(n1892), .B(n1947), .C(n245), .Y(n2433) );
  OAI21X1 U1917 ( .A(n1892), .B(n1949), .C(n247), .Y(n2432) );
  OAI21X1 U1918 ( .A(n1892), .B(n1951), .C(n249), .Y(n2431) );
  OAI21X1 U1919 ( .A(n1892), .B(n1953), .C(n251), .Y(n2430) );
  OAI21X1 U1920 ( .A(n1892), .B(n1955), .C(n253), .Y(n2429) );
  OAI21X1 U1921 ( .A(n1893), .B(n1925), .C(n255), .Y(n2428) );
  OAI21X1 U1922 ( .A(n1893), .B(n1927), .C(n257), .Y(n2427) );
  OAI21X1 U1923 ( .A(n1893), .B(n1929), .C(n259), .Y(n2426) );
  OAI21X1 U1924 ( .A(n1893), .B(n1931), .C(n261), .Y(n2425) );
  OAI21X1 U1925 ( .A(n1893), .B(n1933), .C(n263), .Y(n2424) );
  OAI21X1 U1926 ( .A(n1893), .B(n1935), .C(n265), .Y(n2423) );
  OAI21X1 U1927 ( .A(n1893), .B(n1937), .C(n267), .Y(n2422) );
  OAI21X1 U1928 ( .A(n1893), .B(n1939), .C(n269), .Y(n2421) );
  OAI21X1 U1929 ( .A(n1894), .B(n1941), .C(n271), .Y(n2420) );
  OAI21X1 U1930 ( .A(n1894), .B(n1943), .C(n273), .Y(n2419) );
  OAI21X1 U1931 ( .A(n1894), .B(n1945), .C(n275), .Y(n2418) );
  OAI21X1 U1932 ( .A(n1894), .B(n1947), .C(n277), .Y(n2417) );
  OAI21X1 U1933 ( .A(n1894), .B(n1949), .C(n279), .Y(n2416) );
  OAI21X1 U1934 ( .A(n1894), .B(n1951), .C(n281), .Y(n2415) );
  OAI21X1 U1935 ( .A(n1894), .B(n1953), .C(n283), .Y(n2414) );
  OAI21X1 U1936 ( .A(n1894), .B(n1955), .C(n285), .Y(n2413) );
  OAI21X1 U1937 ( .A(n1895), .B(n1925), .C(n287), .Y(n2412) );
  OAI21X1 U1938 ( .A(n1895), .B(n1927), .C(n289), .Y(n2411) );
  OAI21X1 U1939 ( .A(n1895), .B(n1929), .C(n291), .Y(n2410) );
  OAI21X1 U1940 ( .A(n1895), .B(n1931), .C(n293), .Y(n2409) );
  OAI21X1 U1941 ( .A(n1895), .B(n1933), .C(n295), .Y(n2408) );
  OAI21X1 U1942 ( .A(n1895), .B(n1935), .C(n297), .Y(n2407) );
  OAI21X1 U1943 ( .A(n1895), .B(n1937), .C(n299), .Y(n2406) );
  OAI21X1 U1944 ( .A(n1895), .B(n1939), .C(n301), .Y(n2405) );
  OAI21X1 U1945 ( .A(n1896), .B(n1941), .C(n303), .Y(n2404) );
  OAI21X1 U1946 ( .A(n1896), .B(n1943), .C(n305), .Y(n2403) );
  OAI21X1 U1947 ( .A(n1896), .B(n1945), .C(n307), .Y(n2402) );
  OAI21X1 U1948 ( .A(n1896), .B(n1947), .C(n309), .Y(n2401) );
  OAI21X1 U1949 ( .A(n1896), .B(n1949), .C(n311), .Y(n2400) );
  OAI21X1 U1950 ( .A(n1896), .B(n1951), .C(n313), .Y(n2399) );
  OAI21X1 U1951 ( .A(n1896), .B(n1953), .C(n315), .Y(n2398) );
  OAI21X1 U1952 ( .A(n1896), .B(n1955), .C(n317), .Y(n2397) );
  OAI21X1 U1953 ( .A(n1897), .B(n1925), .C(n319), .Y(n2396) );
  OAI21X1 U1954 ( .A(n1897), .B(n1927), .C(n321), .Y(n2395) );
  OAI21X1 U1955 ( .A(n1897), .B(n1929), .C(n323), .Y(n2394) );
  OAI21X1 U1956 ( .A(n1897), .B(n1931), .C(n325), .Y(n2393) );
  OAI21X1 U1957 ( .A(n1897), .B(n1933), .C(n327), .Y(n2392) );
  OAI21X1 U1958 ( .A(n1897), .B(n1935), .C(n329), .Y(n2391) );
  OAI21X1 U1959 ( .A(n1897), .B(n1937), .C(n331), .Y(n2390) );
  OAI21X1 U1960 ( .A(n1897), .B(n1939), .C(n333), .Y(n2389) );
  OAI21X1 U1961 ( .A(n1898), .B(n1941), .C(n335), .Y(n2388) );
  OAI21X1 U1962 ( .A(n1898), .B(n1943), .C(n337), .Y(n2387) );
  OAI21X1 U1963 ( .A(n1898), .B(n1945), .C(n339), .Y(n2386) );
  OAI21X1 U1964 ( .A(n1898), .B(n1947), .C(n341), .Y(n2385) );
  OAI21X1 U1965 ( .A(n1898), .B(n1949), .C(n343), .Y(n2384) );
  OAI21X1 U1966 ( .A(n1898), .B(n1951), .C(n345), .Y(n2383) );
  OAI21X1 U1967 ( .A(n1898), .B(n1953), .C(n347), .Y(n2382) );
  OAI21X1 U1968 ( .A(n1898), .B(n1955), .C(n349), .Y(n2381) );
  OAI21X1 U1969 ( .A(n1899), .B(n1925), .C(n351), .Y(n2380) );
  OAI21X1 U1970 ( .A(n1899), .B(n1927), .C(n353), .Y(n2379) );
  OAI21X1 U1971 ( .A(n1899), .B(n1929), .C(n355), .Y(n2378) );
  OAI21X1 U1972 ( .A(n1899), .B(n1931), .C(n357), .Y(n2377) );
  OAI21X1 U1973 ( .A(n1899), .B(n1933), .C(n359), .Y(n2376) );
  OAI21X1 U1974 ( .A(n1899), .B(n1935), .C(n361), .Y(n2375) );
  OAI21X1 U1975 ( .A(n1899), .B(n1937), .C(n363), .Y(n2374) );
  OAI21X1 U1976 ( .A(n1899), .B(n1939), .C(n365), .Y(n2373) );
  OAI21X1 U1977 ( .A(n1900), .B(n1941), .C(n367), .Y(n2372) );
  OAI21X1 U1978 ( .A(n1900), .B(n1943), .C(n369), .Y(n2371) );
  OAI21X1 U1979 ( .A(n1900), .B(n1945), .C(n371), .Y(n2370) );
  OAI21X1 U1980 ( .A(n1900), .B(n1947), .C(n373), .Y(n2369) );
  OAI21X1 U1981 ( .A(n1900), .B(n1949), .C(n375), .Y(n2368) );
  OAI21X1 U1982 ( .A(n1900), .B(n1951), .C(n377), .Y(n2367) );
  OAI21X1 U1983 ( .A(n1900), .B(n1953), .C(n379), .Y(n2366) );
  OAI21X1 U1984 ( .A(n1900), .B(n1955), .C(n381), .Y(n2365) );
  OAI21X1 U1985 ( .A(n1901), .B(n1925), .C(n383), .Y(n2364) );
  OAI21X1 U1986 ( .A(n1901), .B(n1927), .C(n385), .Y(n2363) );
  OAI21X1 U1987 ( .A(n1901), .B(n1929), .C(n387), .Y(n2362) );
  OAI21X1 U1988 ( .A(n1901), .B(n1931), .C(n389), .Y(n2361) );
  OAI21X1 U1989 ( .A(n1901), .B(n1933), .C(n391), .Y(n2360) );
  OAI21X1 U1990 ( .A(n1901), .B(n1935), .C(n393), .Y(n2359) );
  OAI21X1 U1991 ( .A(n1901), .B(n1937), .C(n395), .Y(n2358) );
  OAI21X1 U1992 ( .A(n1901), .B(n1939), .C(n397), .Y(n2357) );
  OAI21X1 U1993 ( .A(n1902), .B(n1941), .C(n399), .Y(n2356) );
  OAI21X1 U1994 ( .A(n1902), .B(n1943), .C(n401), .Y(n2355) );
  OAI21X1 U1995 ( .A(n1902), .B(n1945), .C(n403), .Y(n2354) );
  OAI21X1 U1996 ( .A(n1902), .B(n1947), .C(n405), .Y(n2353) );
  OAI21X1 U1997 ( .A(n1902), .B(n1949), .C(n407), .Y(n2352) );
  OAI21X1 U1998 ( .A(n1902), .B(n1951), .C(n409), .Y(n2351) );
  OAI21X1 U1999 ( .A(n1902), .B(n1953), .C(n411), .Y(n2350) );
  OAI21X1 U2000 ( .A(n1902), .B(n1955), .C(n413), .Y(n2349) );
  OAI21X1 U2001 ( .A(n1903), .B(n1925), .C(n415), .Y(n2348) );
  OAI21X1 U2002 ( .A(n1903), .B(n1927), .C(n417), .Y(n2347) );
  OAI21X1 U2003 ( .A(n1903), .B(n1929), .C(n419), .Y(n2346) );
  OAI21X1 U2004 ( .A(n1903), .B(n1931), .C(n421), .Y(n2345) );
  OAI21X1 U2005 ( .A(n1903), .B(n1933), .C(n423), .Y(n2344) );
  OAI21X1 U2006 ( .A(n1903), .B(n1935), .C(n425), .Y(n2343) );
  OAI21X1 U2007 ( .A(n1903), .B(n1937), .C(n427), .Y(n2342) );
  OAI21X1 U2008 ( .A(n1903), .B(n1939), .C(n429), .Y(n2341) );
  OAI21X1 U2009 ( .A(n1904), .B(n1941), .C(n431), .Y(n2340) );
  OAI21X1 U2010 ( .A(n1904), .B(n1943), .C(n433), .Y(n2339) );
  OAI21X1 U2011 ( .A(n1904), .B(n1945), .C(n435), .Y(n2338) );
  OAI21X1 U2012 ( .A(n1904), .B(n1947), .C(n437), .Y(n2337) );
  OAI21X1 U2013 ( .A(n1904), .B(n1949), .C(n439), .Y(n2336) );
  OAI21X1 U2014 ( .A(n1904), .B(n1951), .C(n441), .Y(n2335) );
  OAI21X1 U2015 ( .A(n1904), .B(n1953), .C(n443), .Y(n2334) );
  OAI21X1 U2016 ( .A(n1904), .B(n1955), .C(n445), .Y(n2333) );
  NAND2X1 U2017 ( .A(\mem<8><0> ), .B(n619), .Y(n2121) );
  OAI21X1 U2018 ( .A(n1905), .B(n1925), .C(n2121), .Y(n2332) );
  NAND2X1 U2019 ( .A(\mem<8><1> ), .B(n619), .Y(n2122) );
  OAI21X1 U2020 ( .A(n1905), .B(n1927), .C(n2122), .Y(n2331) );
  NAND2X1 U2021 ( .A(\mem<8><2> ), .B(n619), .Y(n2123) );
  OAI21X1 U2022 ( .A(n1905), .B(n1929), .C(n2123), .Y(n2330) );
  NAND2X1 U2023 ( .A(\mem<8><3> ), .B(n619), .Y(n2124) );
  OAI21X1 U2024 ( .A(n1905), .B(n1931), .C(n2124), .Y(n2329) );
  NAND2X1 U2025 ( .A(\mem<8><4> ), .B(n619), .Y(n2125) );
  OAI21X1 U2026 ( .A(n1905), .B(n1933), .C(n2125), .Y(n2328) );
  NAND2X1 U2027 ( .A(\mem<8><5> ), .B(n619), .Y(n2126) );
  OAI21X1 U2028 ( .A(n1905), .B(n1935), .C(n2126), .Y(n2327) );
  NAND2X1 U2029 ( .A(\mem<8><6> ), .B(n619), .Y(n2127) );
  OAI21X1 U2030 ( .A(n1905), .B(n1937), .C(n2127), .Y(n2326) );
  NAND2X1 U2031 ( .A(\mem<8><7> ), .B(n619), .Y(n2128) );
  OAI21X1 U2032 ( .A(n1905), .B(n1939), .C(n2128), .Y(n2325) );
  NAND2X1 U2033 ( .A(\mem<8><8> ), .B(n619), .Y(n2129) );
  OAI21X1 U2034 ( .A(n1905), .B(n1942), .C(n2129), .Y(n2324) );
  NAND2X1 U2035 ( .A(\mem<8><9> ), .B(n619), .Y(n2130) );
  OAI21X1 U2036 ( .A(n1905), .B(n1944), .C(n2130), .Y(n2323) );
  NAND2X1 U2037 ( .A(\mem<8><10> ), .B(n619), .Y(n2131) );
  OAI21X1 U2038 ( .A(n1905), .B(n1946), .C(n2131), .Y(n2322) );
  NAND2X1 U2039 ( .A(\mem<8><11> ), .B(n619), .Y(n2132) );
  OAI21X1 U2040 ( .A(n1905), .B(n1948), .C(n2132), .Y(n2321) );
  NAND2X1 U2041 ( .A(\mem<8><12> ), .B(n619), .Y(n2133) );
  OAI21X1 U2042 ( .A(n1905), .B(n1950), .C(n2133), .Y(n2320) );
  NAND2X1 U2043 ( .A(\mem<8><13> ), .B(n619), .Y(n2134) );
  OAI21X1 U2044 ( .A(n1905), .B(n1952), .C(n2134), .Y(n2319) );
  NAND2X1 U2045 ( .A(\mem<8><14> ), .B(n619), .Y(n2135) );
  OAI21X1 U2046 ( .A(n1905), .B(n1954), .C(n2135), .Y(n2318) );
  NAND2X1 U2047 ( .A(\mem<8><15> ), .B(n619), .Y(n2136) );
  OAI21X1 U2048 ( .A(n1905), .B(n1956), .C(n2136), .Y(n2317) );
  NAND3X1 U2049 ( .A(n1965), .B(n2701), .C(n1967), .Y(n2137) );
  NAND2X1 U2050 ( .A(\mem<7><0> ), .B(n1211), .Y(n2138) );
  OAI21X1 U2051 ( .A(n1906), .B(n1926), .C(n2138), .Y(n2316) );
  OAI21X1 U2052 ( .A(n1906), .B(n1927), .C(n447), .Y(n2315) );
  OAI21X1 U2053 ( .A(n1906), .B(n1929), .C(n449), .Y(n2314) );
  OAI21X1 U2054 ( .A(n1906), .B(n1931), .C(n451), .Y(n2313) );
  OAI21X1 U2055 ( .A(n1906), .B(n1933), .C(n453), .Y(n2312) );
  OAI21X1 U2056 ( .A(n1906), .B(n1935), .C(n455), .Y(n2311) );
  OAI21X1 U2057 ( .A(n1906), .B(n1937), .C(n457), .Y(n2310) );
  OAI21X1 U2058 ( .A(n1906), .B(n1939), .C(n459), .Y(n2309) );
  OAI21X1 U2059 ( .A(n1907), .B(n1941), .C(n461), .Y(n2308) );
  OAI21X1 U2060 ( .A(n1907), .B(n1943), .C(n463), .Y(n2307) );
  OAI21X1 U2061 ( .A(n1907), .B(n1945), .C(n465), .Y(n2306) );
  OAI21X1 U2062 ( .A(n1907), .B(n1947), .C(n467), .Y(n2305) );
  OAI21X1 U2063 ( .A(n1907), .B(n1949), .C(n469), .Y(n2304) );
  OAI21X1 U2064 ( .A(n1907), .B(n1951), .C(n471), .Y(n2303) );
  OAI21X1 U2065 ( .A(n1907), .B(n1953), .C(n473), .Y(n2302) );
  OAI21X1 U2066 ( .A(n1907), .B(n1955), .C(n475), .Y(n2301) );
  NAND2X1 U2067 ( .A(\mem<6><0> ), .B(n1214), .Y(n2139) );
  OAI21X1 U2068 ( .A(n1908), .B(n1926), .C(n2139), .Y(n2300) );
  OAI21X1 U2069 ( .A(n1908), .B(n1927), .C(n477), .Y(n2299) );
  OAI21X1 U2070 ( .A(n1908), .B(n1929), .C(n479), .Y(n2298) );
  OAI21X1 U2071 ( .A(n1908), .B(n1931), .C(n481), .Y(n2297) );
  OAI21X1 U2072 ( .A(n1908), .B(n1933), .C(n483), .Y(n2296) );
  OAI21X1 U2073 ( .A(n1908), .B(n1935), .C(n485), .Y(n2295) );
  OAI21X1 U2074 ( .A(n1908), .B(n1937), .C(n487), .Y(n2294) );
  OAI21X1 U2075 ( .A(n1908), .B(n1939), .C(n489), .Y(n2293) );
  OAI21X1 U2076 ( .A(n1909), .B(n1941), .C(n491), .Y(n2292) );
  OAI21X1 U2077 ( .A(n1909), .B(n1943), .C(n493), .Y(n2291) );
  OAI21X1 U2078 ( .A(n1909), .B(n1945), .C(n495), .Y(n2290) );
  OAI21X1 U2079 ( .A(n1909), .B(n1947), .C(n497), .Y(n2289) );
  OAI21X1 U2080 ( .A(n1909), .B(n1949), .C(n499), .Y(n2288) );
  OAI21X1 U2081 ( .A(n1909), .B(n1951), .C(n501), .Y(n2287) );
  OAI21X1 U2082 ( .A(n1909), .B(n1953), .C(n503), .Y(n2286) );
  OAI21X1 U2083 ( .A(n1909), .B(n1955), .C(n505), .Y(n2285) );
  NAND2X1 U2084 ( .A(\mem<5><0> ), .B(n1217), .Y(n2141) );
  OAI21X1 U2085 ( .A(n1910), .B(n1926), .C(n2141), .Y(n2284) );
  NAND2X1 U2086 ( .A(\mem<5><1> ), .B(n1217), .Y(n2142) );
  OAI21X1 U2087 ( .A(n1910), .B(n1928), .C(n2142), .Y(n2283) );
  NAND2X1 U2088 ( .A(\mem<5><2> ), .B(n1217), .Y(n2143) );
  OAI21X1 U2089 ( .A(n1910), .B(n1930), .C(n2143), .Y(n2282) );
  NAND2X1 U2090 ( .A(\mem<5><3> ), .B(n1217), .Y(n2144) );
  OAI21X1 U2091 ( .A(n1910), .B(n1932), .C(n2144), .Y(n2281) );
  NAND2X1 U2092 ( .A(\mem<5><4> ), .B(n1217), .Y(n2145) );
  OAI21X1 U2093 ( .A(n1910), .B(n1934), .C(n2145), .Y(n2280) );
  NAND2X1 U2094 ( .A(\mem<5><5> ), .B(n1217), .Y(n2146) );
  OAI21X1 U2095 ( .A(n1910), .B(n1936), .C(n2146), .Y(n2279) );
  NAND2X1 U2096 ( .A(\mem<5><6> ), .B(n1217), .Y(n2147) );
  OAI21X1 U2097 ( .A(n1910), .B(n1938), .C(n2147), .Y(n2278) );
  NAND2X1 U2098 ( .A(\mem<5><7> ), .B(n1217), .Y(n2148) );
  OAI21X1 U2099 ( .A(n1910), .B(n1940), .C(n2148), .Y(n2277) );
  OAI21X1 U2100 ( .A(n1911), .B(n1941), .C(n507), .Y(n2276) );
  OAI21X1 U2101 ( .A(n1911), .B(n1943), .C(n509), .Y(n2275) );
  OAI21X1 U2102 ( .A(n1911), .B(n1945), .C(n511), .Y(n2274) );
  OAI21X1 U2103 ( .A(n1911), .B(n1947), .C(n513), .Y(n2273) );
  OAI21X1 U2104 ( .A(n1911), .B(n1949), .C(n515), .Y(n2272) );
  OAI21X1 U2105 ( .A(n1911), .B(n1951), .C(n517), .Y(n2271) );
  OAI21X1 U2106 ( .A(n1911), .B(n1953), .C(n519), .Y(n2270) );
  OAI21X1 U2107 ( .A(n1911), .B(n1955), .C(n521), .Y(n2269) );
  NAND2X1 U2108 ( .A(\mem<4><0> ), .B(n1220), .Y(n2150) );
  OAI21X1 U2109 ( .A(n1912), .B(n1926), .C(n2150), .Y(n2268) );
  OAI21X1 U2110 ( .A(n1912), .B(n1927), .C(n523), .Y(n2267) );
  OAI21X1 U2111 ( .A(n1912), .B(n1929), .C(n525), .Y(n2266) );
  OAI21X1 U2112 ( .A(n1912), .B(n1931), .C(n527), .Y(n2265) );
  OAI21X1 U2113 ( .A(n1912), .B(n1933), .C(n529), .Y(n2264) );
  OAI21X1 U2114 ( .A(n1912), .B(n1935), .C(n531), .Y(n2263) );
  OAI21X1 U2115 ( .A(n1912), .B(n1937), .C(n533), .Y(n2262) );
  OAI21X1 U2116 ( .A(n1912), .B(n1939), .C(n535), .Y(n2261) );
  OAI21X1 U2117 ( .A(n1913), .B(n1941), .C(n537), .Y(n2260) );
  OAI21X1 U2118 ( .A(n1913), .B(n1943), .C(n539), .Y(n2259) );
  OAI21X1 U2119 ( .A(n1913), .B(n1945), .C(n541), .Y(n2258) );
  OAI21X1 U2120 ( .A(n1913), .B(n1947), .C(n543), .Y(n2257) );
  OAI21X1 U2121 ( .A(n1913), .B(n1949), .C(n545), .Y(n2256) );
  OAI21X1 U2122 ( .A(n1913), .B(n1951), .C(n547), .Y(n2255) );
  OAI21X1 U2123 ( .A(n1913), .B(n1953), .C(n549), .Y(n2254) );
  OAI21X1 U2124 ( .A(n1913), .B(n1955), .C(n551), .Y(n2253) );
  NAND2X1 U2125 ( .A(\mem<3><0> ), .B(n1223), .Y(n2152) );
  OAI21X1 U2126 ( .A(n1914), .B(n1926), .C(n2152), .Y(n2252) );
  OAI21X1 U2127 ( .A(n1914), .B(n1927), .C(n553), .Y(n2251) );
  OAI21X1 U2128 ( .A(n1914), .B(n1929), .C(n555), .Y(n2250) );
  OAI21X1 U2129 ( .A(n1914), .B(n1931), .C(n557), .Y(n2249) );
  OAI21X1 U2130 ( .A(n1914), .B(n1933), .C(n559), .Y(n2248) );
  OAI21X1 U2131 ( .A(n1914), .B(n1935), .C(n561), .Y(n2247) );
  OAI21X1 U2132 ( .A(n1914), .B(n1937), .C(n563), .Y(n2246) );
  OAI21X1 U2133 ( .A(n1914), .B(n1939), .C(n565), .Y(n2245) );
  NAND2X1 U2134 ( .A(\mem<3><8> ), .B(n1222), .Y(n2153) );
  OAI21X1 U2135 ( .A(n1915), .B(n1942), .C(n2153), .Y(n2244) );
  NAND2X1 U2136 ( .A(\mem<3><9> ), .B(n1222), .Y(n2154) );
  OAI21X1 U2137 ( .A(n1915), .B(n1944), .C(n2154), .Y(n2243) );
  NAND2X1 U2138 ( .A(\mem<3><10> ), .B(n1222), .Y(n2155) );
  OAI21X1 U2139 ( .A(n1915), .B(n1946), .C(n2155), .Y(n2242) );
  NAND2X1 U2140 ( .A(\mem<3><11> ), .B(n1222), .Y(n2156) );
  OAI21X1 U2141 ( .A(n1915), .B(n1948), .C(n2156), .Y(n2241) );
  NAND2X1 U2142 ( .A(\mem<3><12> ), .B(n1222), .Y(n2157) );
  OAI21X1 U2143 ( .A(n1915), .B(n1950), .C(n2157), .Y(n2240) );
  NAND2X1 U2144 ( .A(\mem<3><13> ), .B(n1222), .Y(n2158) );
  OAI21X1 U2145 ( .A(n1915), .B(n1952), .C(n2158), .Y(n2239) );
  NAND2X1 U2146 ( .A(\mem<3><14> ), .B(n1222), .Y(n2159) );
  OAI21X1 U2147 ( .A(n1915), .B(n1954), .C(n2159), .Y(n2238) );
  OAI21X1 U2148 ( .A(n1915), .B(n1956), .C(n567), .Y(n2237) );
  NAND2X1 U2149 ( .A(\mem<2><0> ), .B(n1226), .Y(n2161) );
  OAI21X1 U2150 ( .A(n1916), .B(n1926), .C(n2161), .Y(n2236) );
  NAND2X1 U2151 ( .A(\mem<2><1> ), .B(n1226), .Y(n2162) );
  OAI21X1 U2152 ( .A(n1916), .B(n1928), .C(n2162), .Y(n2235) );
  NAND2X1 U2153 ( .A(\mem<2><2> ), .B(n1226), .Y(n2163) );
  OAI21X1 U2154 ( .A(n1916), .B(n1930), .C(n2163), .Y(n2234) );
  NAND2X1 U2155 ( .A(\mem<2><3> ), .B(n1226), .Y(n2164) );
  OAI21X1 U2156 ( .A(n1916), .B(n1932), .C(n2164), .Y(n2233) );
  NAND2X1 U2157 ( .A(\mem<2><4> ), .B(n1226), .Y(n2165) );
  OAI21X1 U2158 ( .A(n1916), .B(n1934), .C(n2165), .Y(n2232) );
  NAND2X1 U2159 ( .A(\mem<2><5> ), .B(n1226), .Y(n2166) );
  OAI21X1 U2160 ( .A(n1916), .B(n1936), .C(n2166), .Y(n2231) );
  NAND2X1 U2161 ( .A(\mem<2><6> ), .B(n1226), .Y(n2167) );
  OAI21X1 U2162 ( .A(n1916), .B(n1938), .C(n2167), .Y(n2230) );
  NAND2X1 U2163 ( .A(\mem<2><7> ), .B(n1226), .Y(n2168) );
  OAI21X1 U2164 ( .A(n1916), .B(n1940), .C(n2168), .Y(n2229) );
  OAI21X1 U2165 ( .A(n1917), .B(n1941), .C(n569), .Y(n2228) );
  OAI21X1 U2166 ( .A(n1917), .B(n1943), .C(n571), .Y(n2227) );
  OAI21X1 U2167 ( .A(n1917), .B(n1945), .C(n573), .Y(n2226) );
  OAI21X1 U2168 ( .A(n1917), .B(n1947), .C(n575), .Y(n2225) );
  OAI21X1 U2169 ( .A(n1917), .B(n1949), .C(n577), .Y(n2224) );
  OAI21X1 U2170 ( .A(n1917), .B(n1951), .C(n579), .Y(n2223) );
  OAI21X1 U2171 ( .A(n1917), .B(n1953), .C(n581), .Y(n2222) );
  OAI21X1 U2172 ( .A(n1917), .B(n1955), .C(n583), .Y(n2221) );
  NAND2X1 U2173 ( .A(\mem<1><0> ), .B(n1229), .Y(n2170) );
  OAI21X1 U2174 ( .A(n1918), .B(n1926), .C(n2170), .Y(n2220) );
  OAI21X1 U2175 ( .A(n1918), .B(n1927), .C(n585), .Y(n2219) );
  OAI21X1 U2176 ( .A(n1918), .B(n1929), .C(n587), .Y(n2218) );
  OAI21X1 U2177 ( .A(n1918), .B(n1931), .C(n589), .Y(n2217) );
  OAI21X1 U2178 ( .A(n1918), .B(n1933), .C(n591), .Y(n2216) );
  OAI21X1 U2179 ( .A(n1918), .B(n1935), .C(n593), .Y(n2215) );
  OAI21X1 U2180 ( .A(n1918), .B(n1937), .C(n595), .Y(n2214) );
  OAI21X1 U2181 ( .A(n1918), .B(n1939), .C(n597), .Y(n2213) );
  OAI21X1 U2182 ( .A(n1919), .B(n1941), .C(n599), .Y(n2212) );
  OAI21X1 U2183 ( .A(n1919), .B(n1943), .C(n601), .Y(n2211) );
  OAI21X1 U2184 ( .A(n1919), .B(n1945), .C(n603), .Y(n2210) );
  OAI21X1 U2185 ( .A(n1919), .B(n1947), .C(n605), .Y(n2209) );
  OAI21X1 U2186 ( .A(n1919), .B(n1949), .C(n607), .Y(n2208) );
  OAI21X1 U2187 ( .A(n1919), .B(n1951), .C(n609), .Y(n2207) );
  OAI21X1 U2188 ( .A(n1919), .B(n1953), .C(n611), .Y(n2206) );
  OAI21X1 U2189 ( .A(n1919), .B(n1955), .C(n613), .Y(n2205) );
  NAND2X1 U2190 ( .A(\mem<0><0> ), .B(n621), .Y(n2173) );
  OAI21X1 U2191 ( .A(n1920), .B(n1926), .C(n2173), .Y(n2204) );
  NAND2X1 U2192 ( .A(\mem<0><1> ), .B(n621), .Y(n2174) );
  OAI21X1 U2193 ( .A(n1920), .B(n1927), .C(n2174), .Y(n2203) );
  NAND2X1 U2194 ( .A(\mem<0><2> ), .B(n621), .Y(n2175) );
  OAI21X1 U2195 ( .A(n1920), .B(n1929), .C(n2175), .Y(n2202) );
  NAND2X1 U2196 ( .A(\mem<0><3> ), .B(n621), .Y(n2176) );
  OAI21X1 U2197 ( .A(n1920), .B(n1931), .C(n2176), .Y(n2201) );
  NAND2X1 U2198 ( .A(\mem<0><4> ), .B(n621), .Y(n2177) );
  OAI21X1 U2199 ( .A(n1920), .B(n1933), .C(n2177), .Y(n2200) );
  NAND2X1 U2200 ( .A(\mem<0><5> ), .B(n621), .Y(n2178) );
  OAI21X1 U2201 ( .A(n1920), .B(n1935), .C(n2178), .Y(n2199) );
  NAND2X1 U2202 ( .A(\mem<0><6> ), .B(n621), .Y(n2179) );
  OAI21X1 U2203 ( .A(n1920), .B(n1937), .C(n2179), .Y(n2198) );
  NAND2X1 U2204 ( .A(\mem<0><7> ), .B(n621), .Y(n2180) );
  OAI21X1 U2205 ( .A(n1920), .B(n1939), .C(n2180), .Y(n2197) );
  NAND2X1 U2206 ( .A(\mem<0><8> ), .B(n621), .Y(n2181) );
  OAI21X1 U2207 ( .A(n1920), .B(n1941), .C(n2181), .Y(n2196) );
  NAND2X1 U2208 ( .A(\mem<0><9> ), .B(n621), .Y(n2182) );
  OAI21X1 U2209 ( .A(n1920), .B(n1943), .C(n2182), .Y(n2195) );
  NAND2X1 U2210 ( .A(\mem<0><10> ), .B(n621), .Y(n2183) );
  OAI21X1 U2211 ( .A(n1920), .B(n1945), .C(n2183), .Y(n2194) );
  NAND2X1 U2212 ( .A(\mem<0><11> ), .B(n621), .Y(n2184) );
  OAI21X1 U2213 ( .A(n1920), .B(n1947), .C(n2184), .Y(n2193) );
  NAND2X1 U2214 ( .A(\mem<0><12> ), .B(n621), .Y(n2185) );
  OAI21X1 U2215 ( .A(n1920), .B(n1949), .C(n2185), .Y(n2192) );
  NAND2X1 U2216 ( .A(\mem<0><13> ), .B(n621), .Y(n2186) );
  OAI21X1 U2217 ( .A(n1920), .B(n1951), .C(n2186), .Y(n2191) );
  NAND2X1 U2218 ( .A(\mem<0><14> ), .B(n621), .Y(n2187) );
  OAI21X1 U2219 ( .A(n1920), .B(n1953), .C(n2187), .Y(n2190) );
  NAND2X1 U2220 ( .A(\mem<0><15> ), .B(n621), .Y(n2188) );
  OAI21X1 U2221 ( .A(n1920), .B(n1955), .C(n2188), .Y(n2189) );
endmodule


module memc_Size16_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2232), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2233), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2234), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2235), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2236), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2237), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2238), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2239), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2240), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2241), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2242), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2243), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2244), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2245), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2246), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2247), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2248), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2249), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2250), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2251), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2252), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2253), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2254), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2255), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2256), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2257), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2258), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2259), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2260), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2261), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2262), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2263), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2264), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2265), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2266), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2267), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2268), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2269), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2270), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2271), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2272), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2273), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2274), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2275), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2276), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2277), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2278), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2279), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2280), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2281), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2282), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2283), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2284), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2285), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2286), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2287), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2288), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2289), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2290), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2291), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2292), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2293), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2294), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2295), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2296), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2297), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2298), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2299), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2300), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2301), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2302), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2303), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2304), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2305), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2306), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2307), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2308), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2309), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2310), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2311), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2312), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2313), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2314), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2315), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2316), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2317), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2318), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2319), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2320), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2321), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2322), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2323), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2324), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2325), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2326), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2327), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2328), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2329), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2330), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2331), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2332), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2333), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2334), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2335), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2336), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2337), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2338), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2339), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2340), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2341), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2342), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2343), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2344), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2345), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2346), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2347), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2348), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2349), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2350), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2351), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2352), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2353), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2354), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2355), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2356), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2357), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2358), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2359), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2360), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2361), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2362), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2363), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2364), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2365), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2366), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2367), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2368), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2369), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2370), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2371), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2372), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2373), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2374), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2375), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2376), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2377), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2378), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2379), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2380), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2381), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2382), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2383), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2384), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2385), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2386), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2387), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2388), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2389), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2390), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2391), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2392), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2393), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2394), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2395), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2396), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2397), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2398), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2399), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2400), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2401), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2402), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2403), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2404), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2405), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2406), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2407), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2408), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2409), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2410), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2411), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2412), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2413), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2414), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2415), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2416), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2417), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2418), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2419), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2420), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2421), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2422), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2423), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2424), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2425), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2426), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2427), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2428), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2429), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2430), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2431), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2432), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2433), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2434), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2435), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2436), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2437), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2438), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2439), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2440), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2441), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2442), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2443), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2444), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2445), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2446), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2447), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2448), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2449), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2450), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2451), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2452), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2453), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2454), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2455), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2456), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2457), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2458), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2459), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2460), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2461), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2462), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2463), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2464), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2465), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2466), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2467), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2468), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2469), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2470), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2471), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2472), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2473), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2474), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2475), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2476), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2477), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2478), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2479), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2480), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2481), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2482), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2483), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2484), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2485), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2486), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2487), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2488), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2489), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2490), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2491), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2492), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2493), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2494), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2495), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2496), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2497), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2498), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2499), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2500), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2501), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2502), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2503), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2504), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2505), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2506), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2507), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2508), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2509), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2510), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2511), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2512), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2513), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2514), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2515), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2516), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2517), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2518), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2519), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2520), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2521), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2522), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2523), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2524), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2525), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2526), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2527), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2528), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2529), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2530), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2531), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2532), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2533), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2534), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2535), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2536), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2537), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2538), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2539), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2540), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2541), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2542), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2543), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2544), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2545), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2546), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2547), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2548), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2549), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2550), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2551), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2552), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2553), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2554), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2555), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2556), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2557), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2558), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2559), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2560), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2561), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2562), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2563), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2564), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2565), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2566), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2567), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2568), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2569), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2570), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2571), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2572), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2573), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2574), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2575), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2576), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2577), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2578), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2579), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2580), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2581), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2582), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2583), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2584), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2585), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2586), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2587), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2588), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2589), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2590), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2591), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2592), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2593), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2594), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2595), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2596), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2597), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2598), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2599), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2600), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2601), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2602), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2603), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2604), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2605), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2606), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2607), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2608), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2609), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2610), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2611), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2612), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2613), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2614), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2615), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2616), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2617), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2618), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2619), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2620), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2621), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2622), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2623), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2624), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2625), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2626), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2627), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2628), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2629), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2630), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2631), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2632), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2633), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2634), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2635), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2636), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2637), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2638), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2639), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2640), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2641), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2642), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2643), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2644), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2645), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2646), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2647), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2648), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2649), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2650), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2651), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2652), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2653), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2654), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2655), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2656), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2657), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2658), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2659), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2660), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2661), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2662), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2663), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2664), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2665), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2666), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2667), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2668), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2669), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2670), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2671), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2672), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2673), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2674), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2675), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2676), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2677), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2678), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2679), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2680), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2681), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2682), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2683), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2684), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2685), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2686), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2687), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2688), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2689), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2690), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2691), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2692), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2693), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2694), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2695), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2696), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2697), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2698), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2699), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2700), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2701), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2702), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2703), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2704), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2705), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2706), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2707), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2708), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2709), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2710), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2711), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2712), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2713), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2714), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2715), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2716), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2717), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2718), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2719), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2720), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2721), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2722), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2723), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2724), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2725), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2726), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2727), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2728), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2729), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2730), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2731), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2732), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2733), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2734), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2735), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2736), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2737), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2738), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2739), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2740), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2741), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2742), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2743), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2744) );
  INVX4 U2 ( .A(n48), .Y(n49) );
  INVX4 U3 ( .A(n46), .Y(n47) );
  INVX4 U4 ( .A(n44), .Y(n45) );
  INVX4 U5 ( .A(n42), .Y(n43) );
  INVX4 U6 ( .A(n40), .Y(n41) );
  INVX4 U7 ( .A(n38), .Y(n39) );
  INVX4 U8 ( .A(n36), .Y(n37) );
  INVX4 U9 ( .A(n34), .Y(n35) );
  INVX4 U10 ( .A(n50), .Y(n51) );
  INVX4 U11 ( .A(n32), .Y(n33) );
  INVX4 U12 ( .A(n30), .Y(n31) );
  INVX4 U13 ( .A(n28), .Y(n29) );
  INVX4 U14 ( .A(n26), .Y(n27) );
  INVX4 U15 ( .A(n24), .Y(n25) );
  INVX4 U16 ( .A(n22), .Y(n23) );
  INVX4 U17 ( .A(n20), .Y(n21) );
  INVX4 U18 ( .A(n18), .Y(n19) );
  INVX4 U19 ( .A(n16), .Y(n17) );
  INVX4 U20 ( .A(n14), .Y(n15) );
  INVX4 U21 ( .A(n12), .Y(n13) );
  INVX4 U22 ( .A(n10), .Y(n11) );
  INVX4 U23 ( .A(n8), .Y(n9) );
  INVX4 U24 ( .A(n6), .Y(n7) );
  INVX4 U25 ( .A(n4), .Y(n5) );
  INVX8 U26 ( .A(n1363), .Y(n1996) );
  INVX2 U27 ( .A(write), .Y(n111) );
  INVX1 U28 ( .A(n2034), .Y(n1883) );
  INVX1 U29 ( .A(n2036), .Y(n1882) );
  INVX1 U30 ( .A(n2036), .Y(n1881) );
  INVX1 U31 ( .A(n2034), .Y(n1884) );
  INVX1 U32 ( .A(n1887), .Y(n1888) );
  INVX2 U33 ( .A(n1887), .Y(n1890) );
  INVX1 U34 ( .A(n1887), .Y(n1892) );
  INVX2 U35 ( .A(n1887), .Y(n1893) );
  INVX2 U36 ( .A(n1887), .Y(n1894) );
  INVX1 U37 ( .A(n1865), .Y(N32) );
  INVX1 U38 ( .A(n1869), .Y(N28) );
  INVX1 U39 ( .A(n1871), .Y(N26) );
  INVX1 U40 ( .A(n1873), .Y(N24) );
  INVX1 U41 ( .A(n1874), .Y(N23) );
  INVX1 U42 ( .A(n1875), .Y(N22) );
  INVX1 U43 ( .A(n1876), .Y(N21) );
  INVX1 U44 ( .A(n1866), .Y(N31) );
  INVX1 U45 ( .A(n1867), .Y(N30) );
  INVX1 U46 ( .A(n1868), .Y(N29) );
  INVX1 U47 ( .A(n1870), .Y(N27) );
  INVX1 U48 ( .A(n1872), .Y(N25) );
  INVX1 U49 ( .A(n1877), .Y(N20) );
  INVX1 U50 ( .A(n1878), .Y(N19) );
  INVX1 U51 ( .A(n1879), .Y(N18) );
  INVX1 U52 ( .A(n1880), .Y(N17) );
  BUFX2 U53 ( .A(n1308), .Y(n1932) );
  BUFX2 U54 ( .A(n1310), .Y(n1934) );
  BUFX2 U55 ( .A(n1312), .Y(n1936) );
  BUFX2 U56 ( .A(n1314), .Y(n1938) );
  BUFX2 U57 ( .A(n1316), .Y(n1940) );
  BUFX2 U58 ( .A(n1318), .Y(n1942) );
  BUFX2 U59 ( .A(n1320), .Y(n1944) );
  BUFX2 U60 ( .A(n1322), .Y(n1947) );
  BUFX2 U61 ( .A(n1324), .Y(n1949) );
  BUFX2 U62 ( .A(n1326), .Y(n1951) );
  BUFX2 U63 ( .A(n1328), .Y(n1953) );
  BUFX2 U64 ( .A(n1330), .Y(n1955) );
  BUFX2 U65 ( .A(n1332), .Y(n1957) );
  BUFX2 U66 ( .A(n1334), .Y(n1959) );
  BUFX2 U67 ( .A(n1336), .Y(n1962) );
  BUFX2 U68 ( .A(n1338), .Y(n1964) );
  BUFX2 U69 ( .A(n1340), .Y(n1966) );
  BUFX2 U70 ( .A(n1342), .Y(n1968) );
  BUFX2 U71 ( .A(n1344), .Y(n1970) );
  BUFX2 U72 ( .A(n1346), .Y(n1972) );
  BUFX2 U73 ( .A(n1348), .Y(n1974) );
  BUFX2 U74 ( .A(n1350), .Y(n1977) );
  BUFX2 U75 ( .A(n1352), .Y(n1979) );
  BUFX2 U76 ( .A(n1354), .Y(n1981) );
  BUFX2 U77 ( .A(n1356), .Y(n1983) );
  BUFX2 U78 ( .A(n1358), .Y(n1985) );
  BUFX2 U79 ( .A(n1360), .Y(n1987) );
  BUFX2 U80 ( .A(n1362), .Y(n1989) );
  INVX1 U81 ( .A(n104), .Y(n2025) );
  INVX4 U82 ( .A(n1898), .Y(n1887) );
  INVX4 U83 ( .A(n2028), .Y(n1927) );
  INVX1 U84 ( .A(n1887), .Y(n1896) );
  INVX1 U85 ( .A(n1887), .Y(n1889) );
  INVX1 U86 ( .A(n1887), .Y(n1897) );
  INVX1 U87 ( .A(n1887), .Y(n1895) );
  INVX1 U88 ( .A(n1887), .Y(n1891) );
  BUFX2 U89 ( .A(n1308), .Y(n1933) );
  INVX1 U90 ( .A(n2036), .Y(n2035) );
  INVX1 U91 ( .A(N14), .Y(n2036) );
  INVX1 U92 ( .A(n1927), .Y(n1928) );
  INVX4 U93 ( .A(n1928), .Y(n1899) );
  BUFX2 U94 ( .A(n1310), .Y(n1935) );
  BUFX2 U95 ( .A(n1312), .Y(n1937) );
  BUFX2 U96 ( .A(n1314), .Y(n1939) );
  BUFX2 U97 ( .A(n1316), .Y(n1941) );
  BUFX2 U98 ( .A(n1318), .Y(n1943) );
  BUFX2 U99 ( .A(n1320), .Y(n1945) );
  INVX1 U100 ( .A(n2034), .Y(n2033) );
  INVX1 U101 ( .A(N13), .Y(n2034) );
  INVX1 U102 ( .A(n1305), .Y(n1976) );
  INVX1 U103 ( .A(n1306), .Y(n1991) );
  INVX1 U104 ( .A(n2030), .Y(n1898) );
  BUFX2 U105 ( .A(n1324), .Y(n1950) );
  BUFX2 U106 ( .A(n1326), .Y(n1952) );
  BUFX2 U107 ( .A(n1328), .Y(n1954) );
  BUFX2 U108 ( .A(n1330), .Y(n1956) );
  BUFX2 U109 ( .A(n1332), .Y(n1958) );
  BUFX2 U110 ( .A(n1334), .Y(n1960) );
  BUFX2 U111 ( .A(n1340), .Y(n1967) );
  BUFX2 U112 ( .A(n1342), .Y(n1969) );
  BUFX2 U113 ( .A(n1344), .Y(n1971) );
  BUFX2 U114 ( .A(n1346), .Y(n1973) );
  BUFX2 U115 ( .A(n1348), .Y(n1975) );
  BUFX2 U116 ( .A(n1354), .Y(n1982) );
  BUFX2 U117 ( .A(n1356), .Y(n1984) );
  BUFX2 U118 ( .A(n1358), .Y(n1986) );
  BUFX2 U119 ( .A(n1360), .Y(n1988) );
  BUFX2 U120 ( .A(n1362), .Y(n1990) );
  BUFX2 U121 ( .A(n1322), .Y(n1948) );
  BUFX2 U122 ( .A(n1336), .Y(n1963) );
  BUFX2 U123 ( .A(n1350), .Y(n1978) );
  INVX1 U124 ( .A(n1303), .Y(n1946) );
  BUFX2 U125 ( .A(n1338), .Y(n1965) );
  BUFX2 U126 ( .A(n1352), .Y(n1980) );
  INVX1 U127 ( .A(n1304), .Y(n1961) );
  AND2X2 U128 ( .A(\mem<30><15> ), .B(n127), .Y(n1) );
  INVX1 U129 ( .A(n1), .Y(n2) );
  AND2X2 U130 ( .A(n111), .B(n2027), .Y(n3) );
  AND2X2 U131 ( .A(n1994), .B(n1321), .Y(n4) );
  AND2X2 U132 ( .A(n1994), .B(n1323), .Y(n6) );
  AND2X2 U133 ( .A(n1994), .B(n1325), .Y(n8) );
  AND2X2 U134 ( .A(n1994), .B(n1327), .Y(n10) );
  AND2X2 U135 ( .A(n1992), .B(n1329), .Y(n12) );
  AND2X2 U136 ( .A(n1992), .B(n1331), .Y(n14) );
  AND2X2 U137 ( .A(n1992), .B(n1333), .Y(n16) );
  AND2X2 U138 ( .A(n1992), .B(n1304), .Y(n18) );
  AND2X2 U139 ( .A(n1992), .B(n1335), .Y(n20) );
  AND2X2 U140 ( .A(n1992), .B(n1337), .Y(n22) );
  AND2X2 U141 ( .A(n1992), .B(n1339), .Y(n24) );
  AND2X2 U142 ( .A(n1992), .B(n1341), .Y(n26) );
  AND2X2 U143 ( .A(n1992), .B(n1343), .Y(n28) );
  AND2X2 U144 ( .A(n1992), .B(n1345), .Y(n30) );
  AND2X2 U145 ( .A(n1992), .B(n1347), .Y(n32) );
  AND2X2 U146 ( .A(n1993), .B(n1305), .Y(n34) );
  AND2X2 U147 ( .A(n1993), .B(n1349), .Y(n36) );
  AND2X2 U148 ( .A(n1993), .B(n1351), .Y(n38) );
  AND2X2 U149 ( .A(n1993), .B(n1353), .Y(n40) );
  AND2X2 U150 ( .A(n1993), .B(n1355), .Y(n42) );
  AND2X2 U151 ( .A(n1993), .B(n1357), .Y(n44) );
  AND2X2 U152 ( .A(n1993), .B(n1359), .Y(n46) );
  AND2X2 U153 ( .A(n1993), .B(n1361), .Y(n48) );
  AND2X2 U154 ( .A(n1992), .B(n1306), .Y(n50) );
  AND2X2 U155 ( .A(n1992), .B(n1307), .Y(n52) );
  AND2X2 U156 ( .A(n1994), .B(n1309), .Y(n53) );
  AND2X2 U157 ( .A(n1993), .B(n1303), .Y(n54) );
  AND2X2 U158 ( .A(n1993), .B(n1311), .Y(n55) );
  AND2X2 U159 ( .A(n1992), .B(n1313), .Y(n56) );
  AND2X2 U160 ( .A(n106), .B(n1315), .Y(n57) );
  AND2X2 U161 ( .A(n106), .B(n1317), .Y(n58) );
  AND2X2 U162 ( .A(n106), .B(n1319), .Y(n59) );
  AND2X2 U163 ( .A(\mem<19><15> ), .B(n13), .Y(n60) );
  INVX1 U164 ( .A(n60), .Y(n61) );
  AND2X2 U165 ( .A(\mem<15><15> ), .B(n21), .Y(n62) );
  INVX1 U166 ( .A(n62), .Y(n63) );
  AND2X2 U167 ( .A(\mem<14><15> ), .B(n23), .Y(n64) );
  INVX1 U168 ( .A(n64), .Y(n65) );
  AND2X2 U169 ( .A(\mem<13><15> ), .B(n25), .Y(n66) );
  INVX1 U170 ( .A(n66), .Y(n67) );
  AND2X2 U171 ( .A(\mem<12><15> ), .B(n27), .Y(n68) );
  INVX1 U172 ( .A(n68), .Y(n69) );
  AND2X2 U173 ( .A(\mem<11><15> ), .B(n29), .Y(n70) );
  INVX1 U174 ( .A(n70), .Y(n71) );
  AND2X2 U175 ( .A(\mem<10><15> ), .B(n31), .Y(n72) );
  INVX1 U176 ( .A(n72), .Y(n73) );
  AND2X2 U177 ( .A(\mem<9><15> ), .B(n33), .Y(n74) );
  INVX1 U178 ( .A(n74), .Y(n75) );
  AND2X2 U179 ( .A(\mem<7><0> ), .B(n37), .Y(n76) );
  INVX1 U180 ( .A(n76), .Y(n77) );
  AND2X2 U181 ( .A(\mem<7><15> ), .B(n37), .Y(n78) );
  INVX1 U182 ( .A(n78), .Y(n79) );
  AND2X2 U183 ( .A(\mem<6><15> ), .B(n39), .Y(n80) );
  INVX1 U184 ( .A(n80), .Y(n81) );
  AND2X2 U185 ( .A(\mem<5><15> ), .B(n41), .Y(n82) );
  INVX1 U186 ( .A(n82), .Y(n83) );
  AND2X2 U187 ( .A(\mem<4><15> ), .B(n43), .Y(n84) );
  INVX1 U188 ( .A(n84), .Y(n85) );
  AND2X2 U189 ( .A(\mem<3><15> ), .B(n45), .Y(n86) );
  INVX1 U190 ( .A(n86), .Y(n87) );
  AND2X2 U191 ( .A(\mem<2><15> ), .B(n47), .Y(n88) );
  INVX1 U192 ( .A(n88), .Y(n89) );
  AND2X2 U193 ( .A(\mem<1><15> ), .B(n49), .Y(n90) );
  INVX1 U194 ( .A(n90), .Y(n91) );
  AND2X2 U195 ( .A(\data_in<1> ), .B(n1994), .Y(n92) );
  AND2X2 U196 ( .A(\data_in<2> ), .B(n1994), .Y(n93) );
  AND2X2 U197 ( .A(\data_in<3> ), .B(n1994), .Y(n94) );
  AND2X2 U198 ( .A(\data_in<4> ), .B(n1994), .Y(n95) );
  AND2X2 U199 ( .A(\data_in<5> ), .B(n1994), .Y(n96) );
  AND2X2 U200 ( .A(\data_in<6> ), .B(n1994), .Y(n97) );
  AND2X2 U201 ( .A(\data_in<7> ), .B(n1994), .Y(n98) );
  AND2X2 U202 ( .A(\data_in<8> ), .B(n1994), .Y(n99) );
  AND2X2 U203 ( .A(\data_in<9> ), .B(n1994), .Y(n100) );
  AND2X2 U204 ( .A(\data_in<10> ), .B(n1994), .Y(n101) );
  AND2X2 U205 ( .A(\data_in<15> ), .B(n1993), .Y(n102) );
  AND2X2 U206 ( .A(\data_in<15> ), .B(n1993), .Y(n103) );
  INVX1 U207 ( .A(n103), .Y(n104) );
  INVX1 U208 ( .A(n103), .Y(n105) );
  AND2X2 U209 ( .A(n2027), .B(write), .Y(n106) );
  AND2X2 U210 ( .A(\data_in<11> ), .B(n1993), .Y(n107) );
  AND2X2 U211 ( .A(\data_in<12> ), .B(n1993), .Y(n108) );
  AND2X2 U212 ( .A(\data_in<13> ), .B(n1993), .Y(n109) );
  AND2X2 U213 ( .A(\data_in<14> ), .B(n1993), .Y(n110) );
  AND2X1 U214 ( .A(N32), .B(n2027), .Y(n112) );
  AND2X2 U215 ( .A(n111), .B(n113), .Y(\data_out<8> ) );
  AND2X1 U216 ( .A(n2027), .B(N24), .Y(n113) );
  AND2X2 U217 ( .A(\mem<29><15> ), .B(n128), .Y(n114) );
  INVX1 U218 ( .A(n114), .Y(n115) );
  AND2X2 U219 ( .A(\mem<28><15> ), .B(n130), .Y(n116) );
  INVX1 U220 ( .A(n116), .Y(n117) );
  AND2X2 U221 ( .A(\mem<27><15> ), .B(n132), .Y(n118) );
  INVX1 U222 ( .A(n118), .Y(n119) );
  AND2X2 U223 ( .A(\mem<26><15> ), .B(n134), .Y(n120) );
  INVX1 U224 ( .A(n120), .Y(n121) );
  AND2X2 U225 ( .A(\mem<25><15> ), .B(n136), .Y(n122) );
  INVX1 U226 ( .A(n122), .Y(n123) );
  INVX1 U227 ( .A(n52), .Y(n124) );
  INVX1 U228 ( .A(n52), .Y(n125) );
  INVX1 U229 ( .A(n53), .Y(n126) );
  INVX1 U230 ( .A(n53), .Y(n127) );
  INVX1 U231 ( .A(n55), .Y(n128) );
  INVX1 U232 ( .A(n55), .Y(n129) );
  INVX1 U233 ( .A(n56), .Y(n130) );
  INVX1 U234 ( .A(n56), .Y(n131) );
  INVX1 U235 ( .A(n57), .Y(n132) );
  INVX1 U236 ( .A(n57), .Y(n133) );
  INVX1 U237 ( .A(n58), .Y(n134) );
  INVX1 U238 ( .A(n58), .Y(n135) );
  INVX1 U239 ( .A(n59), .Y(n136) );
  INVX1 U240 ( .A(n59), .Y(n137) );
  INVX1 U241 ( .A(n54), .Y(n138) );
  INVX1 U242 ( .A(n54), .Y(n139) );
  INVX1 U243 ( .A(n52), .Y(n140) );
  INVX1 U244 ( .A(n52), .Y(n141) );
  INVX1 U245 ( .A(n53), .Y(n142) );
  INVX1 U246 ( .A(n53), .Y(n143) );
  INVX1 U247 ( .A(n55), .Y(n144) );
  INVX1 U248 ( .A(n55), .Y(n145) );
  INVX1 U249 ( .A(n56), .Y(n146) );
  INVX1 U250 ( .A(n56), .Y(n147) );
  INVX1 U251 ( .A(n57), .Y(n148) );
  INVX1 U252 ( .A(n57), .Y(n149) );
  INVX1 U253 ( .A(n58), .Y(n150) );
  INVX1 U254 ( .A(n58), .Y(n151) );
  INVX1 U255 ( .A(n59), .Y(n152) );
  INVX1 U256 ( .A(n59), .Y(n153) );
  INVX1 U257 ( .A(n54), .Y(n154) );
  INVX1 U258 ( .A(n54), .Y(n155) );
  INVX4 U259 ( .A(n1995), .Y(n1994) );
  AND2X1 U260 ( .A(N28), .B(n2027), .Y(n156) );
  INVX1 U261 ( .A(n2027), .Y(n2026) );
  AND2X2 U262 ( .A(\mem<31><1> ), .B(n125), .Y(n157) );
  INVX1 U263 ( .A(n157), .Y(n158) );
  AND2X2 U264 ( .A(\mem<31><2> ), .B(n125), .Y(n159) );
  INVX1 U265 ( .A(n159), .Y(n160) );
  AND2X2 U266 ( .A(\mem<31><3> ), .B(n124), .Y(n161) );
  INVX1 U267 ( .A(n161), .Y(n162) );
  AND2X2 U268 ( .A(\mem<31><4> ), .B(n124), .Y(n163) );
  INVX1 U269 ( .A(n163), .Y(n164) );
  AND2X2 U270 ( .A(\mem<31><5> ), .B(n124), .Y(n165) );
  INVX1 U271 ( .A(n165), .Y(n166) );
  AND2X2 U272 ( .A(\mem<31><6> ), .B(n125), .Y(n167) );
  INVX1 U273 ( .A(n167), .Y(n168) );
  AND2X2 U274 ( .A(\mem<31><7> ), .B(n124), .Y(n169) );
  INVX1 U275 ( .A(n169), .Y(n170) );
  AND2X2 U276 ( .A(\mem<31><8> ), .B(n140), .Y(n171) );
  INVX1 U277 ( .A(n171), .Y(n172) );
  AND2X2 U278 ( .A(\mem<31><9> ), .B(n140), .Y(n173) );
  INVX1 U279 ( .A(n173), .Y(n174) );
  AND2X2 U280 ( .A(\mem<31><10> ), .B(n141), .Y(n175) );
  INVX1 U281 ( .A(n175), .Y(n176) );
  AND2X2 U282 ( .A(\mem<31><11> ), .B(n141), .Y(n177) );
  INVX1 U283 ( .A(n177), .Y(n178) );
  AND2X2 U284 ( .A(\mem<31><12> ), .B(n140), .Y(n179) );
  INVX1 U285 ( .A(n179), .Y(n180) );
  AND2X2 U286 ( .A(\mem<31><13> ), .B(n141), .Y(n181) );
  INVX1 U287 ( .A(n181), .Y(n182) );
  AND2X2 U288 ( .A(\mem<31><14> ), .B(n141), .Y(n183) );
  INVX1 U289 ( .A(n183), .Y(n184) );
  AND2X2 U290 ( .A(\mem<30><1> ), .B(n142), .Y(n185) );
  INVX1 U291 ( .A(n185), .Y(n186) );
  AND2X2 U292 ( .A(\mem<30><2> ), .B(n143), .Y(n187) );
  INVX1 U293 ( .A(n187), .Y(n188) );
  AND2X2 U294 ( .A(\mem<30><3> ), .B(n142), .Y(n189) );
  INVX1 U295 ( .A(n189), .Y(n190) );
  AND2X2 U296 ( .A(\mem<30><4> ), .B(n143), .Y(n191) );
  INVX1 U297 ( .A(n191), .Y(n192) );
  AND2X2 U298 ( .A(\mem<30><5> ), .B(n142), .Y(n193) );
  INVX1 U299 ( .A(n193), .Y(n194) );
  AND2X2 U300 ( .A(\mem<30><6> ), .B(n143), .Y(n195) );
  INVX1 U301 ( .A(n195), .Y(n196) );
  AND2X2 U302 ( .A(\mem<30><7> ), .B(n142), .Y(n197) );
  INVX1 U303 ( .A(n197), .Y(n198) );
  AND2X2 U304 ( .A(\mem<30><8> ), .B(n127), .Y(n199) );
  INVX1 U305 ( .A(n199), .Y(n200) );
  AND2X2 U306 ( .A(\mem<30><9> ), .B(n127), .Y(n201) );
  INVX1 U307 ( .A(n201), .Y(n202) );
  AND2X2 U308 ( .A(\mem<30><10> ), .B(n126), .Y(n203) );
  INVX1 U309 ( .A(n203), .Y(n204) );
  AND2X2 U310 ( .A(\mem<30><11> ), .B(n126), .Y(n205) );
  INVX1 U311 ( .A(n205), .Y(n206) );
  AND2X2 U312 ( .A(\mem<30><12> ), .B(n126), .Y(n207) );
  INVX1 U313 ( .A(n207), .Y(n208) );
  AND2X2 U314 ( .A(\mem<30><13> ), .B(n127), .Y(n209) );
  INVX1 U315 ( .A(n209), .Y(n210) );
  AND2X2 U316 ( .A(\mem<30><14> ), .B(n126), .Y(n211) );
  INVX1 U317 ( .A(n211), .Y(n212) );
  AND2X2 U318 ( .A(\mem<29><1> ), .B(n145), .Y(n213) );
  INVX1 U319 ( .A(n213), .Y(n215) );
  AND2X2 U320 ( .A(\mem<29><2> ), .B(n145), .Y(n216) );
  INVX1 U321 ( .A(n216), .Y(n217) );
  AND2X2 U322 ( .A(\mem<29><3> ), .B(n144), .Y(n218) );
  INVX1 U323 ( .A(n218), .Y(n219) );
  AND2X2 U324 ( .A(\mem<29><4> ), .B(n145), .Y(n220) );
  INVX1 U325 ( .A(n220), .Y(n221) );
  AND2X2 U326 ( .A(\mem<29><5> ), .B(n144), .Y(n222) );
  INVX1 U327 ( .A(n222), .Y(n223) );
  AND2X2 U328 ( .A(\mem<29><6> ), .B(n128), .Y(n224) );
  INVX1 U329 ( .A(n224), .Y(n225) );
  AND2X2 U330 ( .A(\mem<29><7> ), .B(n144), .Y(n226) );
  INVX1 U331 ( .A(n226), .Y(n227) );
  AND2X2 U332 ( .A(\mem<29><8> ), .B(n129), .Y(n228) );
  INVX1 U333 ( .A(n228), .Y(n229) );
  AND2X2 U334 ( .A(\mem<29><9> ), .B(n129), .Y(n230) );
  INVX1 U335 ( .A(n230), .Y(n231) );
  AND2X2 U336 ( .A(\mem<29><10> ), .B(n144), .Y(n232) );
  INVX1 U337 ( .A(n232), .Y(n233) );
  AND2X2 U338 ( .A(\mem<29><11> ), .B(n129), .Y(n234) );
  INVX1 U339 ( .A(n234), .Y(n235) );
  AND2X2 U340 ( .A(\mem<29><12> ), .B(n129), .Y(n236) );
  INVX1 U341 ( .A(n236), .Y(n237) );
  AND2X2 U342 ( .A(\mem<29><13> ), .B(n128), .Y(n238) );
  INVX1 U343 ( .A(n238), .Y(n239) );
  AND2X2 U344 ( .A(\mem<29><14> ), .B(n128), .Y(n240) );
  INVX1 U345 ( .A(n240), .Y(n241) );
  AND2X2 U346 ( .A(\mem<28><1> ), .B(n147), .Y(n242) );
  INVX1 U347 ( .A(n242), .Y(n243) );
  AND2X2 U348 ( .A(\mem<28><2> ), .B(n147), .Y(n244) );
  INVX1 U349 ( .A(n244), .Y(n245) );
  AND2X2 U350 ( .A(\mem<28><3> ), .B(n146), .Y(n246) );
  INVX1 U351 ( .A(n246), .Y(n247) );
  AND2X2 U352 ( .A(\mem<28><4> ), .B(n147), .Y(n248) );
  INVX1 U353 ( .A(n248), .Y(n249) );
  AND2X2 U354 ( .A(\mem<28><5> ), .B(n146), .Y(n250) );
  INVX1 U355 ( .A(n250), .Y(n251) );
  AND2X2 U356 ( .A(\mem<28><6> ), .B(n130), .Y(n252) );
  INVX1 U357 ( .A(n252), .Y(n253) );
  AND2X2 U358 ( .A(\mem<28><7> ), .B(n146), .Y(n254) );
  INVX1 U359 ( .A(n254), .Y(n255) );
  AND2X2 U360 ( .A(\mem<28><8> ), .B(n131), .Y(n256) );
  INVX1 U361 ( .A(n256), .Y(n257) );
  AND2X2 U362 ( .A(\mem<28><9> ), .B(n131), .Y(n258) );
  INVX1 U363 ( .A(n258), .Y(n259) );
  AND2X2 U364 ( .A(\mem<28><10> ), .B(n146), .Y(n260) );
  INVX1 U365 ( .A(n260), .Y(n261) );
  AND2X2 U366 ( .A(\mem<28><11> ), .B(n131), .Y(n262) );
  INVX1 U367 ( .A(n262), .Y(n263) );
  AND2X2 U368 ( .A(\mem<28><12> ), .B(n131), .Y(n264) );
  INVX1 U369 ( .A(n264), .Y(n265) );
  AND2X2 U370 ( .A(\mem<28><13> ), .B(n130), .Y(n266) );
  INVX1 U371 ( .A(n266), .Y(n267) );
  AND2X2 U372 ( .A(\mem<28><14> ), .B(n130), .Y(n268) );
  INVX1 U373 ( .A(n268), .Y(n269) );
  AND2X2 U374 ( .A(\mem<27><1> ), .B(n149), .Y(n270) );
  INVX1 U375 ( .A(n270), .Y(n271) );
  AND2X2 U376 ( .A(\mem<27><2> ), .B(n149), .Y(n272) );
  INVX1 U377 ( .A(n272), .Y(n273) );
  AND2X2 U378 ( .A(\mem<27><3> ), .B(n148), .Y(n274) );
  INVX1 U379 ( .A(n274), .Y(n275) );
  AND2X2 U380 ( .A(\mem<27><4> ), .B(n149), .Y(n276) );
  INVX1 U381 ( .A(n276), .Y(n277) );
  AND2X2 U382 ( .A(\mem<27><5> ), .B(n148), .Y(n278) );
  INVX1 U383 ( .A(n278), .Y(n279) );
  AND2X2 U384 ( .A(\mem<27><6> ), .B(n132), .Y(n280) );
  INVX1 U385 ( .A(n280), .Y(n281) );
  AND2X2 U386 ( .A(\mem<27><7> ), .B(n148), .Y(n282) );
  INVX1 U387 ( .A(n282), .Y(n283) );
  AND2X2 U388 ( .A(\mem<27><8> ), .B(n133), .Y(n284) );
  INVX1 U389 ( .A(n284), .Y(n285) );
  AND2X2 U390 ( .A(\mem<27><9> ), .B(n133), .Y(n286) );
  INVX1 U391 ( .A(n286), .Y(n287) );
  AND2X2 U392 ( .A(\mem<27><10> ), .B(n148), .Y(n288) );
  INVX1 U393 ( .A(n288), .Y(n289) );
  AND2X2 U394 ( .A(\mem<27><11> ), .B(n133), .Y(n290) );
  INVX1 U395 ( .A(n290), .Y(n291) );
  AND2X2 U396 ( .A(\mem<27><12> ), .B(n133), .Y(n292) );
  INVX1 U397 ( .A(n292), .Y(n293) );
  AND2X2 U398 ( .A(\mem<27><13> ), .B(n132), .Y(n294) );
  INVX1 U399 ( .A(n294), .Y(n295) );
  AND2X2 U400 ( .A(\mem<27><14> ), .B(n132), .Y(n296) );
  INVX1 U401 ( .A(n296), .Y(n297) );
  AND2X2 U402 ( .A(\mem<26><1> ), .B(n151), .Y(n298) );
  INVX1 U403 ( .A(n298), .Y(n299) );
  AND2X2 U404 ( .A(\mem<26><2> ), .B(n151), .Y(n300) );
  INVX1 U405 ( .A(n300), .Y(n301) );
  AND2X2 U406 ( .A(\mem<26><3> ), .B(n150), .Y(n302) );
  INVX1 U407 ( .A(n302), .Y(n303) );
  AND2X2 U408 ( .A(\mem<26><4> ), .B(n151), .Y(n304) );
  INVX1 U409 ( .A(n304), .Y(n305) );
  AND2X2 U410 ( .A(\mem<26><5> ), .B(n150), .Y(n306) );
  INVX1 U411 ( .A(n306), .Y(n307) );
  AND2X2 U412 ( .A(\mem<26><6> ), .B(n134), .Y(n308) );
  INVX1 U413 ( .A(n308), .Y(n309) );
  AND2X2 U414 ( .A(\mem<26><7> ), .B(n150), .Y(n310) );
  INVX1 U415 ( .A(n310), .Y(n311) );
  AND2X2 U416 ( .A(\mem<26><8> ), .B(n135), .Y(n312) );
  INVX1 U417 ( .A(n312), .Y(n313) );
  AND2X2 U418 ( .A(\mem<26><9> ), .B(n135), .Y(n314) );
  INVX1 U419 ( .A(n314), .Y(n315) );
  AND2X2 U420 ( .A(\mem<26><10> ), .B(n150), .Y(n316) );
  INVX1 U421 ( .A(n316), .Y(n317) );
  AND2X2 U422 ( .A(\mem<26><11> ), .B(n135), .Y(n318) );
  INVX1 U423 ( .A(n318), .Y(n319) );
  AND2X2 U424 ( .A(\mem<26><12> ), .B(n135), .Y(n320) );
  INVX1 U425 ( .A(n320), .Y(n321) );
  AND2X2 U426 ( .A(\mem<26><13> ), .B(n134), .Y(n322) );
  INVX1 U427 ( .A(n322), .Y(n323) );
  AND2X2 U428 ( .A(\mem<26><14> ), .B(n134), .Y(n324) );
  INVX1 U429 ( .A(n324), .Y(n325) );
  AND2X2 U430 ( .A(\mem<25><1> ), .B(n153), .Y(n326) );
  INVX1 U431 ( .A(n326), .Y(n327) );
  AND2X2 U432 ( .A(\mem<25><2> ), .B(n153), .Y(n328) );
  INVX1 U433 ( .A(n328), .Y(n329) );
  AND2X2 U434 ( .A(\mem<25><3> ), .B(n152), .Y(n330) );
  INVX1 U435 ( .A(n330), .Y(n331) );
  AND2X2 U436 ( .A(\mem<25><4> ), .B(n153), .Y(n332) );
  INVX1 U437 ( .A(n332), .Y(n333) );
  AND2X2 U438 ( .A(\mem<25><5> ), .B(n152), .Y(n334) );
  INVX1 U439 ( .A(n334), .Y(n335) );
  AND2X2 U440 ( .A(\mem<25><6> ), .B(n136), .Y(n336) );
  INVX1 U441 ( .A(n336), .Y(n337) );
  AND2X2 U442 ( .A(\mem<25><7> ), .B(n152), .Y(n338) );
  INVX1 U443 ( .A(n338), .Y(n339) );
  AND2X2 U444 ( .A(\mem<25><8> ), .B(n137), .Y(n340) );
  INVX1 U445 ( .A(n340), .Y(n341) );
  AND2X2 U446 ( .A(\mem<25><9> ), .B(n137), .Y(n342) );
  INVX1 U447 ( .A(n342), .Y(n343) );
  AND2X2 U448 ( .A(\mem<25><10> ), .B(n152), .Y(n344) );
  INVX1 U449 ( .A(n344), .Y(n345) );
  AND2X2 U450 ( .A(\mem<25><11> ), .B(n137), .Y(n346) );
  INVX1 U451 ( .A(n346), .Y(n347) );
  AND2X2 U452 ( .A(\mem<25><12> ), .B(n137), .Y(n348) );
  INVX1 U453 ( .A(n348), .Y(n349) );
  AND2X2 U454 ( .A(\mem<25><13> ), .B(n136), .Y(n350) );
  INVX1 U455 ( .A(n350), .Y(n351) );
  AND2X2 U456 ( .A(\mem<25><14> ), .B(n136), .Y(n352) );
  INVX1 U457 ( .A(n352), .Y(n353) );
  AND2X2 U458 ( .A(\mem<24><1> ), .B(n155), .Y(n354) );
  INVX1 U459 ( .A(n354), .Y(n355) );
  AND2X2 U460 ( .A(\mem<24><2> ), .B(n154), .Y(n356) );
  INVX1 U461 ( .A(n356), .Y(n357) );
  AND2X2 U462 ( .A(\mem<24><3> ), .B(n154), .Y(n358) );
  INVX1 U463 ( .A(n358), .Y(n359) );
  AND2X2 U464 ( .A(\mem<24><4> ), .B(n154), .Y(n360) );
  INVX1 U465 ( .A(n360), .Y(n361) );
  AND2X2 U466 ( .A(\mem<24><5> ), .B(n155), .Y(n362) );
  INVX1 U467 ( .A(n362), .Y(n363) );
  AND2X2 U468 ( .A(\mem<24><6> ), .B(n155), .Y(n364) );
  INVX1 U469 ( .A(n364), .Y(n365) );
  AND2X2 U470 ( .A(\mem<24><7> ), .B(n155), .Y(n366) );
  INVX1 U471 ( .A(n366), .Y(n367) );
  AND2X2 U472 ( .A(\mem<24><8> ), .B(n138), .Y(n368) );
  INVX1 U473 ( .A(n368), .Y(n369) );
  AND2X2 U474 ( .A(\mem<24><9> ), .B(n139), .Y(n370) );
  INVX1 U475 ( .A(n370), .Y(n371) );
  AND2X2 U476 ( .A(\mem<24><10> ), .B(n139), .Y(n372) );
  INVX1 U477 ( .A(n372), .Y(n373) );
  AND2X2 U478 ( .A(\mem<24><11> ), .B(n138), .Y(n374) );
  INVX1 U479 ( .A(n374), .Y(n375) );
  AND2X2 U480 ( .A(\mem<24><12> ), .B(n138), .Y(n376) );
  INVX1 U481 ( .A(n376), .Y(n377) );
  AND2X2 U482 ( .A(\mem<24><13> ), .B(n139), .Y(n378) );
  INVX1 U483 ( .A(n378), .Y(n379) );
  AND2X2 U484 ( .A(\mem<24><14> ), .B(n138), .Y(n380) );
  INVX1 U485 ( .A(n380), .Y(n381) );
  AND2X2 U486 ( .A(\mem<9><8> ), .B(n33), .Y(n382) );
  INVX1 U487 ( .A(n382), .Y(n383) );
  AND2X2 U488 ( .A(\mem<9><9> ), .B(n33), .Y(n384) );
  INVX1 U489 ( .A(n384), .Y(n385) );
  INVX1 U490 ( .A(n2029), .Y(n2028) );
  AND2X1 U491 ( .A(n2031), .B(n1891), .Y(n386) );
  INVX1 U492 ( .A(n2032), .Y(n2031) );
  AND2X1 U493 ( .A(n2744), .B(n2035), .Y(n387) );
  AND2X2 U494 ( .A(\mem<19><8> ), .B(n13), .Y(n388) );
  INVX1 U495 ( .A(n388), .Y(n389) );
  AND2X2 U496 ( .A(\mem<19><9> ), .B(n13), .Y(n390) );
  INVX1 U497 ( .A(n390), .Y(n391) );
  AND2X2 U498 ( .A(\mem<19><10> ), .B(n13), .Y(n392) );
  INVX1 U499 ( .A(n392), .Y(n393) );
  AND2X2 U500 ( .A(\mem<19><11> ), .B(n13), .Y(n394) );
  INVX1 U501 ( .A(n394), .Y(n395) );
  AND2X2 U502 ( .A(\mem<19><12> ), .B(n13), .Y(n396) );
  INVX1 U503 ( .A(n396), .Y(n397) );
  AND2X2 U504 ( .A(\mem<19><13> ), .B(n13), .Y(n398) );
  INVX1 U505 ( .A(n398), .Y(n399) );
  AND2X2 U506 ( .A(\mem<19><14> ), .B(n13), .Y(n400) );
  INVX1 U507 ( .A(n400), .Y(n401) );
  AND2X2 U508 ( .A(\mem<18><8> ), .B(n15), .Y(n402) );
  INVX1 U509 ( .A(n402), .Y(n403) );
  AND2X2 U510 ( .A(\mem<18><9> ), .B(n15), .Y(n404) );
  INVX1 U511 ( .A(n404), .Y(n405) );
  AND2X2 U512 ( .A(\mem<18><10> ), .B(n15), .Y(n406) );
  INVX1 U513 ( .A(n406), .Y(n407) );
  AND2X2 U514 ( .A(\mem<18><11> ), .B(n15), .Y(n408) );
  INVX1 U515 ( .A(n408), .Y(n409) );
  AND2X2 U516 ( .A(\mem<18><12> ), .B(n15), .Y(n410) );
  INVX1 U517 ( .A(n410), .Y(n411) );
  AND2X2 U518 ( .A(\mem<18><13> ), .B(n15), .Y(n412) );
  INVX1 U519 ( .A(n412), .Y(n413) );
  AND2X2 U520 ( .A(\mem<18><14> ), .B(n15), .Y(n414) );
  INVX1 U521 ( .A(n414), .Y(n415) );
  AND2X2 U522 ( .A(\mem<18><15> ), .B(n15), .Y(n416) );
  INVX1 U523 ( .A(n416), .Y(n417) );
  AND2X2 U524 ( .A(\mem<17><8> ), .B(n17), .Y(n418) );
  INVX1 U525 ( .A(n418), .Y(n419) );
  AND2X2 U526 ( .A(\mem<17><9> ), .B(n17), .Y(n420) );
  INVX1 U527 ( .A(n420), .Y(n421) );
  AND2X2 U528 ( .A(\mem<17><10> ), .B(n17), .Y(n422) );
  INVX1 U529 ( .A(n422), .Y(n423) );
  AND2X2 U530 ( .A(\mem<17><11> ), .B(n17), .Y(n424) );
  INVX1 U531 ( .A(n424), .Y(n425) );
  AND2X2 U532 ( .A(\mem<17><12> ), .B(n17), .Y(n426) );
  INVX1 U533 ( .A(n426), .Y(n427) );
  AND2X2 U534 ( .A(\mem<17><13> ), .B(n17), .Y(n428) );
  INVX1 U535 ( .A(n428), .Y(n429) );
  AND2X2 U536 ( .A(\mem<17><14> ), .B(n17), .Y(n430) );
  INVX1 U537 ( .A(n430), .Y(n431) );
  AND2X2 U538 ( .A(\mem<17><15> ), .B(n17), .Y(n432) );
  INVX1 U539 ( .A(n432), .Y(n433) );
  AND2X2 U540 ( .A(\mem<16><8> ), .B(n19), .Y(n434) );
  INVX1 U541 ( .A(n434), .Y(n435) );
  AND2X2 U542 ( .A(\mem<16><9> ), .B(n19), .Y(n436) );
  INVX1 U543 ( .A(n436), .Y(n437) );
  AND2X2 U544 ( .A(\mem<16><10> ), .B(n19), .Y(n438) );
  INVX1 U545 ( .A(n438), .Y(n439) );
  AND2X2 U546 ( .A(\mem<16><11> ), .B(n19), .Y(n440) );
  INVX1 U547 ( .A(n440), .Y(n441) );
  AND2X2 U548 ( .A(\mem<16><12> ), .B(n19), .Y(n442) );
  INVX1 U549 ( .A(n442), .Y(n443) );
  AND2X2 U550 ( .A(\mem<16><13> ), .B(n19), .Y(n444) );
  INVX1 U551 ( .A(n444), .Y(n445) );
  AND2X2 U552 ( .A(\mem<16><14> ), .B(n19), .Y(n446) );
  INVX1 U553 ( .A(n446), .Y(n447) );
  AND2X2 U554 ( .A(\mem<15><8> ), .B(n21), .Y(n448) );
  INVX1 U555 ( .A(n448), .Y(n449) );
  AND2X2 U556 ( .A(\mem<15><9> ), .B(n21), .Y(n450) );
  INVX1 U557 ( .A(n450), .Y(n451) );
  AND2X2 U558 ( .A(\mem<15><10> ), .B(n21), .Y(n452) );
  INVX1 U559 ( .A(n452), .Y(n453) );
  AND2X2 U560 ( .A(\mem<15><11> ), .B(n21), .Y(n454) );
  INVX1 U561 ( .A(n454), .Y(n455) );
  AND2X2 U562 ( .A(\mem<15><12> ), .B(n21), .Y(n456) );
  INVX1 U563 ( .A(n456), .Y(n457) );
  AND2X2 U564 ( .A(\mem<15><13> ), .B(n21), .Y(n458) );
  INVX1 U565 ( .A(n458), .Y(n459) );
  AND2X2 U566 ( .A(\mem<15><14> ), .B(n21), .Y(n460) );
  INVX1 U567 ( .A(n460), .Y(n461) );
  AND2X2 U568 ( .A(\mem<14><8> ), .B(n23), .Y(n462) );
  INVX1 U569 ( .A(n462), .Y(n463) );
  AND2X2 U570 ( .A(\mem<14><9> ), .B(n23), .Y(n464) );
  INVX1 U571 ( .A(n464), .Y(n465) );
  AND2X2 U572 ( .A(\mem<14><10> ), .B(n23), .Y(n466) );
  INVX1 U573 ( .A(n466), .Y(n467) );
  AND2X2 U574 ( .A(\mem<14><11> ), .B(n23), .Y(n468) );
  INVX1 U575 ( .A(n468), .Y(n469) );
  AND2X2 U576 ( .A(\mem<14><12> ), .B(n23), .Y(n470) );
  INVX1 U577 ( .A(n470), .Y(n471) );
  AND2X2 U578 ( .A(\mem<14><13> ), .B(n23), .Y(n472) );
  INVX1 U579 ( .A(n472), .Y(n473) );
  AND2X2 U580 ( .A(\mem<14><14> ), .B(n23), .Y(n474) );
  INVX1 U581 ( .A(n474), .Y(n475) );
  AND2X2 U582 ( .A(\mem<13><8> ), .B(n25), .Y(n476) );
  INVX1 U583 ( .A(n476), .Y(n477) );
  AND2X2 U584 ( .A(\mem<13><9> ), .B(n25), .Y(n478) );
  INVX1 U585 ( .A(n478), .Y(n479) );
  AND2X2 U586 ( .A(\mem<13><10> ), .B(n25), .Y(n480) );
  INVX1 U587 ( .A(n480), .Y(n481) );
  AND2X2 U588 ( .A(\mem<13><11> ), .B(n25), .Y(n482) );
  INVX1 U589 ( .A(n482), .Y(n483) );
  AND2X2 U590 ( .A(\mem<13><12> ), .B(n25), .Y(n484) );
  INVX1 U591 ( .A(n484), .Y(n485) );
  AND2X2 U592 ( .A(\mem<13><13> ), .B(n25), .Y(n486) );
  INVX1 U593 ( .A(n486), .Y(n487) );
  AND2X2 U594 ( .A(\mem<13><14> ), .B(n25), .Y(n488) );
  INVX1 U595 ( .A(n488), .Y(n489) );
  AND2X2 U596 ( .A(\mem<12><8> ), .B(n27), .Y(n490) );
  INVX1 U597 ( .A(n490), .Y(n491) );
  AND2X2 U598 ( .A(\mem<12><9> ), .B(n27), .Y(n492) );
  INVX1 U599 ( .A(n492), .Y(n493) );
  AND2X2 U600 ( .A(\mem<12><10> ), .B(n27), .Y(n494) );
  INVX1 U601 ( .A(n494), .Y(n495) );
  AND2X2 U602 ( .A(\mem<12><11> ), .B(n27), .Y(n496) );
  INVX1 U603 ( .A(n496), .Y(n497) );
  AND2X2 U604 ( .A(\mem<12><12> ), .B(n27), .Y(n498) );
  INVX1 U605 ( .A(n498), .Y(n499) );
  AND2X2 U606 ( .A(\mem<12><13> ), .B(n27), .Y(n500) );
  INVX1 U607 ( .A(n500), .Y(n501) );
  AND2X2 U608 ( .A(\mem<12><14> ), .B(n27), .Y(n502) );
  INVX1 U609 ( .A(n502), .Y(n503) );
  AND2X2 U610 ( .A(\mem<11><8> ), .B(n29), .Y(n504) );
  INVX1 U611 ( .A(n504), .Y(n505) );
  AND2X2 U612 ( .A(\mem<11><9> ), .B(n29), .Y(n506) );
  INVX1 U613 ( .A(n506), .Y(n507) );
  AND2X2 U614 ( .A(\mem<11><10> ), .B(n29), .Y(n508) );
  INVX1 U615 ( .A(n508), .Y(n509) );
  AND2X2 U616 ( .A(\mem<11><11> ), .B(n29), .Y(n510) );
  INVX1 U617 ( .A(n510), .Y(n511) );
  AND2X2 U618 ( .A(\mem<11><12> ), .B(n29), .Y(n512) );
  INVX1 U619 ( .A(n512), .Y(n513) );
  AND2X2 U620 ( .A(\mem<11><13> ), .B(n29), .Y(n514) );
  INVX1 U621 ( .A(n514), .Y(n515) );
  AND2X2 U622 ( .A(\mem<11><14> ), .B(n29), .Y(n516) );
  INVX1 U623 ( .A(n516), .Y(n517) );
  AND2X2 U624 ( .A(\mem<10><8> ), .B(n31), .Y(n518) );
  INVX1 U625 ( .A(n518), .Y(n519) );
  AND2X2 U626 ( .A(\mem<10><9> ), .B(n31), .Y(n520) );
  INVX1 U627 ( .A(n520), .Y(n521) );
  AND2X2 U628 ( .A(\mem<10><10> ), .B(n31), .Y(n522) );
  INVX1 U629 ( .A(n522), .Y(n523) );
  AND2X2 U630 ( .A(\mem<10><11> ), .B(n31), .Y(n524) );
  INVX1 U631 ( .A(n524), .Y(n525) );
  AND2X2 U632 ( .A(\mem<10><12> ), .B(n31), .Y(n526) );
  INVX1 U633 ( .A(n526), .Y(n527) );
  AND2X2 U634 ( .A(\mem<10><13> ), .B(n31), .Y(n528) );
  INVX1 U635 ( .A(n528), .Y(n529) );
  AND2X2 U636 ( .A(\mem<10><14> ), .B(n31), .Y(n530) );
  INVX1 U637 ( .A(n530), .Y(n531) );
  AND2X2 U638 ( .A(\mem<9><10> ), .B(n33), .Y(n532) );
  INVX1 U639 ( .A(n532), .Y(n533) );
  AND2X2 U640 ( .A(\mem<9><11> ), .B(n33), .Y(n534) );
  INVX1 U641 ( .A(n534), .Y(n535) );
  AND2X2 U642 ( .A(\mem<9><12> ), .B(n33), .Y(n536) );
  INVX1 U643 ( .A(n536), .Y(n537) );
  AND2X2 U644 ( .A(\mem<9><13> ), .B(n33), .Y(n538) );
  INVX1 U645 ( .A(n538), .Y(n539) );
  AND2X2 U646 ( .A(\mem<9><14> ), .B(n33), .Y(n540) );
  INVX1 U647 ( .A(n540), .Y(n541) );
  AND2X2 U648 ( .A(\mem<8><1> ), .B(n35), .Y(n542) );
  INVX1 U649 ( .A(n542), .Y(n543) );
  AND2X2 U650 ( .A(\mem<8><2> ), .B(n35), .Y(n544) );
  INVX1 U651 ( .A(n544), .Y(n545) );
  AND2X2 U652 ( .A(\mem<8><3> ), .B(n35), .Y(n546) );
  INVX1 U653 ( .A(n546), .Y(n547) );
  AND2X2 U654 ( .A(\mem<8><4> ), .B(n35), .Y(n548) );
  INVX1 U655 ( .A(n548), .Y(n549) );
  AND2X2 U656 ( .A(\mem<8><5> ), .B(n35), .Y(n550) );
  INVX1 U657 ( .A(n550), .Y(n551) );
  AND2X2 U658 ( .A(\mem<8><6> ), .B(n35), .Y(n552) );
  INVX1 U659 ( .A(n552), .Y(n553) );
  AND2X2 U660 ( .A(\mem<8><7> ), .B(n35), .Y(n554) );
  INVX1 U661 ( .A(n554), .Y(n555) );
  AND2X2 U662 ( .A(\mem<8><8> ), .B(n35), .Y(n556) );
  INVX1 U663 ( .A(n556), .Y(n557) );
  AND2X2 U664 ( .A(\mem<8><9> ), .B(n35), .Y(n558) );
  INVX1 U665 ( .A(n558), .Y(n559) );
  AND2X2 U666 ( .A(\mem<8><10> ), .B(n35), .Y(n560) );
  INVX1 U667 ( .A(n560), .Y(n561) );
  AND2X2 U668 ( .A(\mem<8><11> ), .B(n35), .Y(n562) );
  INVX1 U669 ( .A(n562), .Y(n563) );
  AND2X2 U670 ( .A(\mem<8><12> ), .B(n35), .Y(n564) );
  INVX1 U671 ( .A(n564), .Y(n565) );
  AND2X2 U672 ( .A(\mem<8><13> ), .B(n35), .Y(n566) );
  INVX1 U673 ( .A(n566), .Y(n567) );
  AND2X2 U674 ( .A(\mem<8><14> ), .B(n35), .Y(n568) );
  INVX1 U675 ( .A(n568), .Y(n569) );
  AND2X2 U676 ( .A(\mem<7><1> ), .B(n37), .Y(n570) );
  INVX1 U677 ( .A(n570), .Y(n571) );
  AND2X2 U678 ( .A(\mem<7><2> ), .B(n37), .Y(n572) );
  INVX1 U679 ( .A(n572), .Y(n573) );
  AND2X2 U680 ( .A(\mem<7><3> ), .B(n37), .Y(n574) );
  INVX1 U681 ( .A(n574), .Y(n575) );
  AND2X2 U682 ( .A(\mem<7><4> ), .B(n37), .Y(n576) );
  INVX1 U683 ( .A(n576), .Y(n577) );
  AND2X2 U684 ( .A(\mem<7><5> ), .B(n37), .Y(n578) );
  INVX1 U685 ( .A(n578), .Y(n579) );
  AND2X2 U686 ( .A(\mem<7><6> ), .B(n37), .Y(n580) );
  INVX1 U687 ( .A(n580), .Y(n581) );
  AND2X2 U688 ( .A(\mem<7><7> ), .B(n37), .Y(n582) );
  INVX1 U689 ( .A(n582), .Y(n583) );
  AND2X2 U690 ( .A(\mem<7><8> ), .B(n37), .Y(n584) );
  INVX1 U691 ( .A(n584), .Y(n585) );
  AND2X2 U692 ( .A(\mem<7><9> ), .B(n37), .Y(n586) );
  INVX1 U693 ( .A(n586), .Y(n587) );
  AND2X2 U694 ( .A(\mem<7><10> ), .B(n37), .Y(n588) );
  INVX1 U695 ( .A(n588), .Y(n589) );
  AND2X2 U696 ( .A(\mem<7><11> ), .B(n37), .Y(n590) );
  INVX1 U697 ( .A(n590), .Y(n591) );
  AND2X2 U698 ( .A(\mem<7><12> ), .B(n37), .Y(n592) );
  INVX1 U699 ( .A(n592), .Y(n593) );
  AND2X2 U700 ( .A(\mem<7><13> ), .B(n37), .Y(n594) );
  INVX1 U701 ( .A(n594), .Y(n595) );
  AND2X2 U702 ( .A(\mem<7><14> ), .B(n37), .Y(n596) );
  INVX1 U703 ( .A(n596), .Y(n597) );
  AND2X2 U704 ( .A(\mem<6><1> ), .B(n39), .Y(n598) );
  INVX1 U705 ( .A(n598), .Y(n599) );
  AND2X2 U706 ( .A(\mem<6><2> ), .B(n39), .Y(n600) );
  INVX1 U707 ( .A(n600), .Y(n601) );
  AND2X2 U708 ( .A(\mem<6><3> ), .B(n39), .Y(n602) );
  INVX1 U709 ( .A(n602), .Y(n603) );
  AND2X2 U710 ( .A(\mem<6><4> ), .B(n39), .Y(n604) );
  INVX1 U711 ( .A(n604), .Y(n605) );
  AND2X2 U712 ( .A(\mem<6><5> ), .B(n39), .Y(n606) );
  INVX1 U713 ( .A(n606), .Y(n607) );
  AND2X2 U714 ( .A(\mem<6><6> ), .B(n39), .Y(n608) );
  INVX1 U715 ( .A(n608), .Y(n609) );
  AND2X2 U716 ( .A(\mem<6><7> ), .B(n39), .Y(n610) );
  INVX1 U717 ( .A(n610), .Y(n611) );
  AND2X2 U718 ( .A(\mem<6><8> ), .B(n39), .Y(n612) );
  INVX1 U719 ( .A(n612), .Y(n613) );
  AND2X2 U720 ( .A(\mem<6><9> ), .B(n39), .Y(n614) );
  INVX1 U721 ( .A(n614), .Y(n615) );
  AND2X2 U722 ( .A(\mem<6><10> ), .B(n39), .Y(n616) );
  INVX1 U723 ( .A(n616), .Y(n617) );
  AND2X2 U724 ( .A(\mem<6><11> ), .B(n39), .Y(n618) );
  INVX1 U725 ( .A(n618), .Y(n619) );
  AND2X2 U726 ( .A(\mem<6><12> ), .B(n39), .Y(n620) );
  INVX1 U727 ( .A(n620), .Y(n621) );
  AND2X2 U728 ( .A(\mem<6><13> ), .B(n39), .Y(n622) );
  INVX1 U729 ( .A(n622), .Y(n623) );
  AND2X2 U730 ( .A(\mem<6><14> ), .B(n39), .Y(n624) );
  INVX1 U731 ( .A(n624), .Y(n625) );
  AND2X2 U732 ( .A(\mem<5><1> ), .B(n41), .Y(n626) );
  INVX1 U733 ( .A(n626), .Y(n627) );
  AND2X2 U734 ( .A(\mem<5><2> ), .B(n41), .Y(n628) );
  INVX1 U735 ( .A(n628), .Y(n629) );
  AND2X2 U736 ( .A(\mem<5><3> ), .B(n41), .Y(n630) );
  INVX1 U737 ( .A(n630), .Y(n631) );
  AND2X2 U738 ( .A(\mem<5><4> ), .B(n41), .Y(n632) );
  INVX1 U739 ( .A(n632), .Y(n633) );
  AND2X2 U740 ( .A(\mem<5><5> ), .B(n41), .Y(n634) );
  INVX1 U741 ( .A(n634), .Y(n635) );
  AND2X2 U742 ( .A(\mem<5><6> ), .B(n41), .Y(n636) );
  INVX1 U743 ( .A(n636), .Y(n637) );
  AND2X2 U744 ( .A(\mem<5><7> ), .B(n41), .Y(n638) );
  INVX1 U745 ( .A(n638), .Y(n639) );
  AND2X2 U746 ( .A(\mem<5><8> ), .B(n41), .Y(n640) );
  INVX1 U747 ( .A(n640), .Y(n641) );
  AND2X2 U748 ( .A(\mem<5><9> ), .B(n41), .Y(n642) );
  INVX1 U749 ( .A(n642), .Y(n643) );
  AND2X2 U750 ( .A(\mem<5><10> ), .B(n41), .Y(n644) );
  INVX1 U751 ( .A(n644), .Y(n645) );
  AND2X2 U752 ( .A(\mem<5><11> ), .B(n41), .Y(n646) );
  INVX1 U753 ( .A(n646), .Y(n647) );
  AND2X2 U754 ( .A(\mem<5><12> ), .B(n41), .Y(n648) );
  INVX1 U755 ( .A(n648), .Y(n649) );
  AND2X2 U756 ( .A(\mem<5><13> ), .B(n41), .Y(n650) );
  INVX1 U757 ( .A(n650), .Y(n1163) );
  AND2X2 U758 ( .A(\mem<5><14> ), .B(n41), .Y(n1164) );
  INVX1 U759 ( .A(n1164), .Y(n1165) );
  AND2X2 U760 ( .A(\mem<4><1> ), .B(n43), .Y(n1166) );
  INVX1 U761 ( .A(n1166), .Y(n1167) );
  AND2X2 U762 ( .A(\mem<4><2> ), .B(n43), .Y(n1168) );
  INVX1 U763 ( .A(n1168), .Y(n1169) );
  AND2X2 U764 ( .A(\mem<4><3> ), .B(n43), .Y(n1170) );
  INVX1 U765 ( .A(n1170), .Y(n1171) );
  AND2X2 U766 ( .A(\mem<4><4> ), .B(n43), .Y(n1172) );
  INVX1 U767 ( .A(n1172), .Y(n1173) );
  AND2X2 U768 ( .A(\mem<4><5> ), .B(n43), .Y(n1174) );
  INVX1 U769 ( .A(n1174), .Y(n1175) );
  AND2X2 U770 ( .A(\mem<4><6> ), .B(n43), .Y(n1176) );
  INVX1 U771 ( .A(n1176), .Y(n1177) );
  AND2X2 U772 ( .A(\mem<4><7> ), .B(n43), .Y(n1178) );
  INVX1 U773 ( .A(n1178), .Y(n1179) );
  AND2X2 U774 ( .A(\mem<4><8> ), .B(n43), .Y(n1180) );
  INVX1 U775 ( .A(n1180), .Y(n1181) );
  AND2X2 U776 ( .A(\mem<4><9> ), .B(n43), .Y(n1182) );
  INVX1 U777 ( .A(n1182), .Y(n1183) );
  AND2X2 U778 ( .A(\mem<4><10> ), .B(n43), .Y(n1184) );
  INVX1 U779 ( .A(n1184), .Y(n1185) );
  AND2X2 U780 ( .A(\mem<4><11> ), .B(n43), .Y(n1186) );
  INVX1 U781 ( .A(n1186), .Y(n1187) );
  AND2X2 U782 ( .A(\mem<4><12> ), .B(n43), .Y(n1188) );
  INVX1 U783 ( .A(n1188), .Y(n1189) );
  AND2X2 U784 ( .A(\mem<4><13> ), .B(n43), .Y(n1190) );
  INVX1 U785 ( .A(n1190), .Y(n1191) );
  AND2X2 U786 ( .A(\mem<4><14> ), .B(n43), .Y(n1192) );
  INVX1 U787 ( .A(n1192), .Y(n1193) );
  AND2X2 U788 ( .A(\mem<3><1> ), .B(n45), .Y(n1194) );
  INVX1 U789 ( .A(n1194), .Y(n1195) );
  AND2X2 U790 ( .A(\mem<3><2> ), .B(n45), .Y(n1196) );
  INVX1 U791 ( .A(n1196), .Y(n1197) );
  AND2X2 U792 ( .A(\mem<3><3> ), .B(n45), .Y(n1198) );
  INVX1 U793 ( .A(n1198), .Y(n1199) );
  AND2X2 U794 ( .A(\mem<3><4> ), .B(n45), .Y(n1200) );
  INVX1 U795 ( .A(n1200), .Y(n1201) );
  AND2X2 U796 ( .A(\mem<3><5> ), .B(n45), .Y(n1202) );
  INVX1 U797 ( .A(n1202), .Y(n1203) );
  AND2X2 U798 ( .A(\mem<3><6> ), .B(n45), .Y(n1204) );
  INVX1 U799 ( .A(n1204), .Y(n1205) );
  AND2X2 U800 ( .A(\mem<3><7> ), .B(n45), .Y(n1206) );
  INVX1 U801 ( .A(n1206), .Y(n1207) );
  AND2X2 U802 ( .A(\mem<3><8> ), .B(n45), .Y(n1208) );
  INVX1 U803 ( .A(n1208), .Y(n1209) );
  AND2X2 U804 ( .A(\mem<3><9> ), .B(n45), .Y(n1210) );
  INVX1 U805 ( .A(n1210), .Y(n1211) );
  AND2X2 U806 ( .A(\mem<3><10> ), .B(n45), .Y(n1212) );
  INVX1 U807 ( .A(n1212), .Y(n1213) );
  AND2X2 U808 ( .A(\mem<3><11> ), .B(n45), .Y(n1214) );
  INVX1 U809 ( .A(n1214), .Y(n1215) );
  AND2X2 U810 ( .A(\mem<3><12> ), .B(n45), .Y(n1216) );
  INVX1 U811 ( .A(n1216), .Y(n1217) );
  AND2X2 U812 ( .A(\mem<3><13> ), .B(n45), .Y(n1218) );
  INVX1 U813 ( .A(n1218), .Y(n1219) );
  AND2X2 U814 ( .A(\mem<3><14> ), .B(n45), .Y(n1220) );
  INVX1 U815 ( .A(n1220), .Y(n1221) );
  AND2X2 U816 ( .A(\mem<2><1> ), .B(n47), .Y(n1222) );
  INVX1 U817 ( .A(n1222), .Y(n1223) );
  AND2X2 U818 ( .A(\mem<2><2> ), .B(n47), .Y(n1224) );
  INVX1 U819 ( .A(n1224), .Y(n1225) );
  AND2X2 U820 ( .A(\mem<2><3> ), .B(n47), .Y(n1226) );
  INVX1 U821 ( .A(n1226), .Y(n1227) );
  AND2X2 U822 ( .A(\mem<2><4> ), .B(n47), .Y(n1228) );
  INVX1 U823 ( .A(n1228), .Y(n1229) );
  AND2X2 U824 ( .A(\mem<2><5> ), .B(n47), .Y(n1230) );
  INVX1 U825 ( .A(n1230), .Y(n1231) );
  AND2X2 U826 ( .A(\mem<2><6> ), .B(n47), .Y(n1232) );
  INVX1 U827 ( .A(n1232), .Y(n1233) );
  AND2X2 U828 ( .A(\mem<2><7> ), .B(n47), .Y(n1234) );
  INVX1 U829 ( .A(n1234), .Y(n1235) );
  AND2X2 U830 ( .A(\mem<2><8> ), .B(n47), .Y(n1236) );
  INVX1 U831 ( .A(n1236), .Y(n1237) );
  AND2X2 U832 ( .A(\mem<2><9> ), .B(n47), .Y(n1238) );
  INVX1 U833 ( .A(n1238), .Y(n1239) );
  AND2X2 U834 ( .A(\mem<2><10> ), .B(n47), .Y(n1240) );
  INVX1 U835 ( .A(n1240), .Y(n1241) );
  AND2X2 U836 ( .A(\mem<2><11> ), .B(n47), .Y(n1242) );
  INVX1 U837 ( .A(n1242), .Y(n1243) );
  AND2X2 U838 ( .A(\mem<2><12> ), .B(n47), .Y(n1244) );
  INVX1 U839 ( .A(n1244), .Y(n1245) );
  AND2X2 U840 ( .A(\mem<2><13> ), .B(n47), .Y(n1246) );
  INVX1 U841 ( .A(n1246), .Y(n1247) );
  AND2X2 U842 ( .A(\mem<2><14> ), .B(n47), .Y(n1248) );
  INVX1 U843 ( .A(n1248), .Y(n1249) );
  AND2X2 U844 ( .A(\mem<1><1> ), .B(n49), .Y(n1250) );
  INVX1 U845 ( .A(n1250), .Y(n1251) );
  AND2X2 U846 ( .A(\mem<1><2> ), .B(n49), .Y(n1252) );
  INVX1 U847 ( .A(n1252), .Y(n1253) );
  AND2X2 U848 ( .A(\mem<1><3> ), .B(n49), .Y(n1254) );
  INVX1 U849 ( .A(n1254), .Y(n1255) );
  AND2X2 U850 ( .A(\mem<1><4> ), .B(n49), .Y(n1256) );
  INVX1 U851 ( .A(n1256), .Y(n1257) );
  AND2X2 U852 ( .A(\mem<1><5> ), .B(n49), .Y(n1258) );
  INVX1 U853 ( .A(n1258), .Y(n1259) );
  AND2X2 U854 ( .A(\mem<1><6> ), .B(n49), .Y(n1260) );
  INVX1 U855 ( .A(n1260), .Y(n1261) );
  AND2X2 U856 ( .A(\mem<1><7> ), .B(n49), .Y(n1262) );
  INVX1 U857 ( .A(n1262), .Y(n1263) );
  AND2X2 U858 ( .A(\mem<1><8> ), .B(n49), .Y(n1264) );
  INVX1 U859 ( .A(n1264), .Y(n1265) );
  AND2X2 U860 ( .A(\mem<1><9> ), .B(n49), .Y(n1266) );
  INVX1 U861 ( .A(n1266), .Y(n1267) );
  AND2X2 U862 ( .A(\mem<1><10> ), .B(n49), .Y(n1268) );
  INVX1 U863 ( .A(n1268), .Y(n1269) );
  AND2X2 U864 ( .A(\mem<1><11> ), .B(n49), .Y(n1270) );
  INVX1 U865 ( .A(n1270), .Y(n1271) );
  AND2X2 U866 ( .A(\mem<1><12> ), .B(n49), .Y(n1272) );
  INVX1 U867 ( .A(n1272), .Y(n1273) );
  AND2X2 U868 ( .A(\mem<1><13> ), .B(n49), .Y(n1274) );
  INVX1 U869 ( .A(n1274), .Y(n1275) );
  AND2X2 U870 ( .A(\mem<1><14> ), .B(n49), .Y(n1276) );
  INVX1 U871 ( .A(n1276), .Y(n1277) );
  AND2X2 U872 ( .A(\mem<0><8> ), .B(n51), .Y(n1278) );
  INVX1 U873 ( .A(n1278), .Y(n1279) );
  AND2X2 U874 ( .A(\mem<0><9> ), .B(n51), .Y(n1280) );
  INVX1 U875 ( .A(n1280), .Y(n1281) );
  AND2X2 U876 ( .A(\mem<0><10> ), .B(n51), .Y(n1282) );
  INVX1 U877 ( .A(n1282), .Y(n1283) );
  AND2X2 U878 ( .A(\mem<0><11> ), .B(n51), .Y(n1284) );
  INVX1 U879 ( .A(n1284), .Y(n1285) );
  AND2X2 U880 ( .A(\mem<0><12> ), .B(n51), .Y(n1286) );
  INVX1 U881 ( .A(n1286), .Y(n1287) );
  AND2X2 U882 ( .A(\mem<0><13> ), .B(n51), .Y(n1288) );
  INVX1 U883 ( .A(n1288), .Y(n1289) );
  AND2X2 U884 ( .A(\mem<0><14> ), .B(n51), .Y(n1290) );
  INVX1 U885 ( .A(n1290), .Y(n1291) );
  BUFX2 U886 ( .A(n2040), .Y(n1292) );
  INVX1 U887 ( .A(n1292), .Y(n2211) );
  BUFX2 U888 ( .A(n2042), .Y(n1293) );
  INVX1 U889 ( .A(n1293), .Y(n2213) );
  BUFX2 U890 ( .A(n2044), .Y(n1294) );
  INVX1 U891 ( .A(n1294), .Y(n2215) );
  BUFX2 U892 ( .A(n2046), .Y(n1295) );
  INVX1 U893 ( .A(n1295), .Y(n2217) );
  BUFX2 U894 ( .A(n2048), .Y(n1296) );
  INVX1 U895 ( .A(n1296), .Y(n2219) );
  BUFX2 U896 ( .A(n2149), .Y(n1297) );
  INVX1 U897 ( .A(n1297), .Y(n2206) );
  BUFX2 U898 ( .A(n2209), .Y(n1298) );
  INVX1 U899 ( .A(n1298), .Y(n2221) );
  AND2X1 U900 ( .A(n2028), .B(n386), .Y(n1299) );
  AND2X1 U901 ( .A(n2033), .B(n387), .Y(n1300) );
  INVX4 U902 ( .A(n93), .Y(n2000) );
  INVX4 U903 ( .A(n94), .Y(n2002) );
  INVX4 U904 ( .A(n95), .Y(n2004) );
  INVX4 U905 ( .A(n96), .Y(n2006) );
  INVX4 U906 ( .A(n97), .Y(n2008) );
  INVX4 U907 ( .A(n98), .Y(n2010) );
  INVX4 U908 ( .A(n99), .Y(n2012) );
  INVX4 U909 ( .A(n100), .Y(n2014) );
  INVX4 U910 ( .A(n101), .Y(n2016) );
  AND2X1 U911 ( .A(n2029), .B(n386), .Y(n1301) );
  AND2X1 U912 ( .A(n2034), .B(n387), .Y(n1302) );
  INVX4 U913 ( .A(n92), .Y(n1998) );
  AND2X1 U914 ( .A(n1300), .B(n2222), .Y(n1303) );
  AND2X1 U915 ( .A(n2222), .B(n1302), .Y(n1304) );
  AND2X1 U916 ( .A(n2222), .B(n2206), .Y(n1305) );
  AND2X1 U917 ( .A(n2222), .B(n2221), .Y(n1306) );
  AND2X1 U918 ( .A(n1299), .B(n1300), .Y(n1307) );
  INVX1 U919 ( .A(n1307), .Y(n1308) );
  AND2X1 U920 ( .A(n1300), .B(n1301), .Y(n1309) );
  INVX1 U921 ( .A(n1309), .Y(n1310) );
  AND2X1 U922 ( .A(n1300), .B(n2211), .Y(n1311) );
  INVX1 U923 ( .A(n1311), .Y(n1312) );
  AND2X1 U924 ( .A(n1300), .B(n2213), .Y(n1313) );
  INVX1 U925 ( .A(n1313), .Y(n1314) );
  AND2X1 U926 ( .A(n1300), .B(n2215), .Y(n1315) );
  INVX1 U927 ( .A(n1315), .Y(n1316) );
  AND2X1 U928 ( .A(n1300), .B(n2217), .Y(n1317) );
  INVX1 U929 ( .A(n1317), .Y(n1318) );
  AND2X1 U930 ( .A(n1300), .B(n2219), .Y(n1319) );
  INVX1 U931 ( .A(n1319), .Y(n1320) );
  AND2X1 U932 ( .A(n1299), .B(n1302), .Y(n1321) );
  INVX1 U933 ( .A(n1321), .Y(n1322) );
  AND2X1 U934 ( .A(n1301), .B(n1302), .Y(n1323) );
  INVX1 U935 ( .A(n1323), .Y(n1324) );
  AND2X1 U936 ( .A(n2211), .B(n1302), .Y(n1325) );
  INVX1 U937 ( .A(n1325), .Y(n1326) );
  AND2X1 U938 ( .A(n2213), .B(n1302), .Y(n1327) );
  INVX1 U939 ( .A(n1327), .Y(n1328) );
  AND2X1 U940 ( .A(n2215), .B(n1302), .Y(n1329) );
  INVX1 U941 ( .A(n1329), .Y(n1330) );
  AND2X1 U942 ( .A(n2217), .B(n1302), .Y(n1331) );
  INVX1 U943 ( .A(n1331), .Y(n1332) );
  AND2X1 U944 ( .A(n2219), .B(n1302), .Y(n1333) );
  INVX1 U945 ( .A(n1333), .Y(n1334) );
  AND2X1 U946 ( .A(n1299), .B(n2206), .Y(n1335) );
  INVX1 U947 ( .A(n1335), .Y(n1336) );
  AND2X1 U948 ( .A(n1301), .B(n2206), .Y(n1337) );
  INVX1 U949 ( .A(n1337), .Y(n1338) );
  AND2X1 U950 ( .A(n2211), .B(n2206), .Y(n1339) );
  INVX1 U951 ( .A(n1339), .Y(n1340) );
  AND2X1 U952 ( .A(n2213), .B(n2206), .Y(n1341) );
  INVX1 U953 ( .A(n1341), .Y(n1342) );
  AND2X1 U954 ( .A(n2215), .B(n2206), .Y(n1343) );
  INVX1 U955 ( .A(n1343), .Y(n1344) );
  AND2X1 U956 ( .A(n2217), .B(n2206), .Y(n1345) );
  INVX1 U957 ( .A(n1345), .Y(n1346) );
  AND2X1 U958 ( .A(n2219), .B(n2206), .Y(n1347) );
  INVX1 U959 ( .A(n1347), .Y(n1348) );
  AND2X1 U960 ( .A(n1299), .B(n2221), .Y(n1349) );
  INVX1 U961 ( .A(n1349), .Y(n1350) );
  AND2X1 U962 ( .A(n1301), .B(n2221), .Y(n1351) );
  INVX1 U963 ( .A(n1351), .Y(n1352) );
  AND2X1 U964 ( .A(n2211), .B(n2221), .Y(n1353) );
  INVX1 U965 ( .A(n1353), .Y(n1354) );
  AND2X1 U966 ( .A(n2213), .B(n2221), .Y(n1355) );
  INVX1 U967 ( .A(n1355), .Y(n1356) );
  AND2X1 U968 ( .A(n2215), .B(n2221), .Y(n1357) );
  INVX1 U969 ( .A(n1357), .Y(n1358) );
  AND2X1 U970 ( .A(n2217), .B(n2221), .Y(n1359) );
  INVX1 U971 ( .A(n1359), .Y(n1360) );
  AND2X1 U972 ( .A(n2219), .B(n2221), .Y(n1361) );
  INVX1 U973 ( .A(n1361), .Y(n1362) );
  AND2X2 U974 ( .A(n106), .B(\data_in<0> ), .Y(n1363) );
  INVX1 U975 ( .A(n2025), .Y(n1364) );
  INVX1 U976 ( .A(n102), .Y(n1365) );
  INVX1 U977 ( .A(n102), .Y(n1366) );
  INVX1 U978 ( .A(n102), .Y(n1367) );
  INVX1 U979 ( .A(n102), .Y(n1368) );
  INVX1 U980 ( .A(n102), .Y(n1369) );
  INVX1 U981 ( .A(n102), .Y(n1370) );
  INVX1 U982 ( .A(n105), .Y(n1371) );
  INVX1 U983 ( .A(n1371), .Y(n1372) );
  INVX1 U984 ( .A(n1371), .Y(n1373) );
  INVX1 U985 ( .A(n1371), .Y(n1374) );
  INVX1 U986 ( .A(n105), .Y(n1375) );
  INVX1 U987 ( .A(n2025), .Y(n1376) );
  INVX1 U988 ( .A(n2025), .Y(n1377) );
  INVX1 U989 ( .A(n1375), .Y(n1378) );
  INVX1 U990 ( .A(n1375), .Y(n1379) );
  INVX1 U991 ( .A(n1375), .Y(n1380) );
  INVX1 U992 ( .A(n1384), .Y(n1381) );
  AND2X1 U993 ( .A(N22), .B(n2027), .Y(n1382) );
  AND2X2 U994 ( .A(n111), .B(n2027), .Y(n1383) );
  INVX1 U995 ( .A(rst), .Y(n2027) );
  INVX1 U996 ( .A(N12), .Y(n2032) );
  OR2X2 U997 ( .A(write), .B(n2026), .Y(n1384) );
  MUX2X1 U998 ( .B(n1386), .A(n1387), .S(n1888), .Y(n1385) );
  MUX2X1 U999 ( .B(n1389), .A(n1390), .S(n1888), .Y(n1388) );
  MUX2X1 U1000 ( .B(n1392), .A(n1393), .S(n1888), .Y(n1391) );
  MUX2X1 U1001 ( .B(n1395), .A(n1396), .S(n1888), .Y(n1394) );
  MUX2X1 U1002 ( .B(n1398), .A(n1399), .S(n1884), .Y(n1397) );
  MUX2X1 U1003 ( .B(n1401), .A(n1402), .S(n1888), .Y(n1400) );
  MUX2X1 U1004 ( .B(n1404), .A(n1405), .S(n1888), .Y(n1403) );
  MUX2X1 U1005 ( .B(n1407), .A(n1408), .S(n1888), .Y(n1406) );
  MUX2X1 U1006 ( .B(n1410), .A(n1411), .S(n1888), .Y(n1409) );
  MUX2X1 U1007 ( .B(n1413), .A(n1414), .S(n1884), .Y(n1412) );
  MUX2X1 U1008 ( .B(n1416), .A(n1417), .S(n1897), .Y(n1415) );
  MUX2X1 U1009 ( .B(n1419), .A(n1420), .S(n1890), .Y(n1418) );
  MUX2X1 U1010 ( .B(n1422), .A(n1423), .S(n1889), .Y(n1421) );
  MUX2X1 U1011 ( .B(n1425), .A(n1426), .S(n1890), .Y(n1424) );
  MUX2X1 U1012 ( .B(n1428), .A(n1429), .S(n1884), .Y(n1427) );
  MUX2X1 U1013 ( .B(n1431), .A(n1432), .S(n1890), .Y(n1430) );
  MUX2X1 U1014 ( .B(n1434), .A(n1435), .S(n1890), .Y(n1433) );
  MUX2X1 U1015 ( .B(n1437), .A(n1438), .S(n1890), .Y(n1436) );
  MUX2X1 U1016 ( .B(n1440), .A(n1441), .S(n1890), .Y(n1439) );
  MUX2X1 U1017 ( .B(n1443), .A(n1444), .S(n1884), .Y(n1442) );
  MUX2X1 U1018 ( .B(n1446), .A(n1447), .S(n1890), .Y(n1445) );
  MUX2X1 U1019 ( .B(n1449), .A(n1450), .S(n1890), .Y(n1448) );
  MUX2X1 U1020 ( .B(n1452), .A(n1453), .S(n1896), .Y(n1451) );
  MUX2X1 U1021 ( .B(n1455), .A(n1456), .S(n1890), .Y(n1454) );
  MUX2X1 U1022 ( .B(n1458), .A(n1459), .S(n1884), .Y(n1457) );
  MUX2X1 U1023 ( .B(n1461), .A(n1462), .S(n1889), .Y(n1460) );
  MUX2X1 U1024 ( .B(n1464), .A(n1465), .S(n1889), .Y(n1463) );
  MUX2X1 U1025 ( .B(n1467), .A(n1468), .S(n1889), .Y(n1466) );
  MUX2X1 U1026 ( .B(n1470), .A(n1471), .S(n1889), .Y(n1469) );
  MUX2X1 U1027 ( .B(n1473), .A(n1474), .S(n1884), .Y(n1472) );
  MUX2X1 U1028 ( .B(n1476), .A(n1477), .S(n1889), .Y(n1475) );
  MUX2X1 U1029 ( .B(n1479), .A(n1480), .S(n1889), .Y(n1478) );
  MUX2X1 U1030 ( .B(n1482), .A(n1483), .S(n1889), .Y(n1481) );
  MUX2X1 U1031 ( .B(n1485), .A(n1486), .S(n1889), .Y(n1484) );
  MUX2X1 U1032 ( .B(n1488), .A(n1489), .S(n1884), .Y(n1487) );
  MUX2X1 U1033 ( .B(n1491), .A(n1492), .S(n1889), .Y(n1490) );
  MUX2X1 U1034 ( .B(n1494), .A(n1495), .S(n1889), .Y(n1493) );
  MUX2X1 U1035 ( .B(n1497), .A(n1498), .S(n1889), .Y(n1496) );
  MUX2X1 U1036 ( .B(n1500), .A(n1501), .S(n1889), .Y(n1499) );
  MUX2X1 U1037 ( .B(n1503), .A(n1504), .S(n1884), .Y(n1502) );
  MUX2X1 U1038 ( .B(n1506), .A(n1507), .S(n1890), .Y(n1505) );
  MUX2X1 U1039 ( .B(n1509), .A(n1510), .S(n1890), .Y(n1508) );
  MUX2X1 U1040 ( .B(n1512), .A(n1513), .S(n1890), .Y(n1511) );
  MUX2X1 U1041 ( .B(n1515), .A(n1516), .S(n1890), .Y(n1514) );
  MUX2X1 U1042 ( .B(n1518), .A(n1519), .S(n1884), .Y(n1517) );
  MUX2X1 U1043 ( .B(n1521), .A(n1522), .S(n1890), .Y(n1520) );
  MUX2X1 U1044 ( .B(n1524), .A(n1525), .S(n1890), .Y(n1523) );
  MUX2X1 U1045 ( .B(n1527), .A(n1528), .S(n1890), .Y(n1526) );
  MUX2X1 U1046 ( .B(n1530), .A(n1531), .S(n1890), .Y(n1529) );
  MUX2X1 U1047 ( .B(n1533), .A(n1534), .S(n1884), .Y(n1532) );
  MUX2X1 U1048 ( .B(n1536), .A(n1537), .S(n1890), .Y(n1535) );
  MUX2X1 U1049 ( .B(n1539), .A(n1540), .S(n1890), .Y(n1538) );
  MUX2X1 U1050 ( .B(n1542), .A(n1543), .S(n1890), .Y(n1541) );
  MUX2X1 U1051 ( .B(n1545), .A(n1546), .S(n1890), .Y(n1544) );
  MUX2X1 U1052 ( .B(n1548), .A(n1549), .S(n1884), .Y(n1547) );
  MUX2X1 U1053 ( .B(n1551), .A(n1552), .S(n1891), .Y(n1550) );
  MUX2X1 U1054 ( .B(n1554), .A(n1555), .S(n1891), .Y(n1553) );
  MUX2X1 U1055 ( .B(n1557), .A(n1558), .S(n1891), .Y(n1556) );
  MUX2X1 U1056 ( .B(n1560), .A(n1561), .S(n1891), .Y(n1559) );
  MUX2X1 U1057 ( .B(n1563), .A(n1564), .S(n1884), .Y(n1562) );
  MUX2X1 U1058 ( .B(n1566), .A(n1567), .S(n1891), .Y(n1565) );
  MUX2X1 U1059 ( .B(n1569), .A(n1570), .S(n1891), .Y(n1568) );
  MUX2X1 U1060 ( .B(n1572), .A(n1573), .S(n1891), .Y(n1571) );
  MUX2X1 U1061 ( .B(n1575), .A(n1576), .S(n1891), .Y(n1574) );
  MUX2X1 U1062 ( .B(n1578), .A(n1579), .S(n1883), .Y(n1577) );
  MUX2X1 U1063 ( .B(n1581), .A(n1582), .S(n1891), .Y(n1580) );
  MUX2X1 U1064 ( .B(n1584), .A(n1585), .S(n1891), .Y(n1583) );
  MUX2X1 U1065 ( .B(n1587), .A(n1588), .S(n1891), .Y(n1586) );
  MUX2X1 U1066 ( .B(n1590), .A(n1591), .S(n1891), .Y(n1589) );
  MUX2X1 U1067 ( .B(n1593), .A(n1594), .S(n1883), .Y(n1592) );
  MUX2X1 U1068 ( .B(n1596), .A(n1597), .S(n1892), .Y(n1595) );
  MUX2X1 U1069 ( .B(n1599), .A(n1600), .S(n1892), .Y(n1598) );
  MUX2X1 U1070 ( .B(n1602), .A(n1603), .S(n1892), .Y(n1601) );
  MUX2X1 U1071 ( .B(n1605), .A(n1606), .S(n1892), .Y(n1604) );
  MUX2X1 U1072 ( .B(n1608), .A(n1609), .S(n1883), .Y(n1607) );
  MUX2X1 U1073 ( .B(n1611), .A(n1612), .S(n1892), .Y(n1610) );
  MUX2X1 U1074 ( .B(n1614), .A(n1615), .S(n1892), .Y(n1613) );
  MUX2X1 U1075 ( .B(n1617), .A(n1618), .S(n1892), .Y(n1616) );
  MUX2X1 U1076 ( .B(n1620), .A(n1621), .S(n1892), .Y(n1619) );
  MUX2X1 U1077 ( .B(n1623), .A(n1624), .S(n1883), .Y(n1622) );
  MUX2X1 U1078 ( .B(n1626), .A(n1627), .S(n1892), .Y(n1625) );
  MUX2X1 U1079 ( .B(n1629), .A(n1630), .S(n1892), .Y(n1628) );
  MUX2X1 U1080 ( .B(n1632), .A(n1633), .S(n1892), .Y(n1631) );
  MUX2X1 U1081 ( .B(n1635), .A(n1636), .S(n1892), .Y(n1634) );
  MUX2X1 U1082 ( .B(n1638), .A(n1639), .S(n1883), .Y(n1637) );
  MUX2X1 U1083 ( .B(n1641), .A(n1642), .S(n1893), .Y(n1640) );
  MUX2X1 U1084 ( .B(n1644), .A(n1645), .S(n1893), .Y(n1643) );
  MUX2X1 U1085 ( .B(n1647), .A(n1648), .S(n1893), .Y(n1646) );
  MUX2X1 U1086 ( .B(n1650), .A(n1651), .S(n1893), .Y(n1649) );
  MUX2X1 U1087 ( .B(n1653), .A(n1654), .S(n1883), .Y(n1652) );
  MUX2X1 U1088 ( .B(n1656), .A(n1657), .S(n1893), .Y(n1655) );
  MUX2X1 U1089 ( .B(n1659), .A(n1660), .S(n1893), .Y(n1658) );
  MUX2X1 U1090 ( .B(n1662), .A(n1663), .S(n1893), .Y(n1661) );
  MUX2X1 U1091 ( .B(n1665), .A(n1666), .S(n1893), .Y(n1664) );
  MUX2X1 U1092 ( .B(n1668), .A(n1669), .S(n1883), .Y(n1667) );
  MUX2X1 U1093 ( .B(n1671), .A(n1672), .S(n1893), .Y(n1670) );
  MUX2X1 U1094 ( .B(n1674), .A(n1675), .S(n1893), .Y(n1673) );
  MUX2X1 U1095 ( .B(n1677), .A(n1678), .S(n1893), .Y(n1676) );
  MUX2X1 U1096 ( .B(n1680), .A(n1681), .S(n1893), .Y(n1679) );
  MUX2X1 U1097 ( .B(n1683), .A(n1684), .S(n1883), .Y(n1682) );
  MUX2X1 U1098 ( .B(n1686), .A(n1687), .S(n1894), .Y(n1685) );
  MUX2X1 U1099 ( .B(n1689), .A(n1690), .S(n1894), .Y(n1688) );
  MUX2X1 U1100 ( .B(n1692), .A(n1693), .S(n1894), .Y(n1691) );
  MUX2X1 U1101 ( .B(n1695), .A(n1696), .S(n1894), .Y(n1694) );
  MUX2X1 U1102 ( .B(n1698), .A(n1699), .S(n1883), .Y(n1697) );
  MUX2X1 U1103 ( .B(n1701), .A(n1702), .S(n1894), .Y(n1700) );
  MUX2X1 U1104 ( .B(n1704), .A(n1705), .S(n1894), .Y(n1703) );
  MUX2X1 U1105 ( .B(n1707), .A(n1708), .S(n1894), .Y(n1706) );
  MUX2X1 U1106 ( .B(n1710), .A(n1711), .S(n1894), .Y(n1709) );
  MUX2X1 U1107 ( .B(n1713), .A(n1714), .S(n1883), .Y(n1712) );
  MUX2X1 U1108 ( .B(n1716), .A(n1717), .S(n1894), .Y(n1715) );
  MUX2X1 U1109 ( .B(n1719), .A(n1720), .S(n1894), .Y(n1718) );
  MUX2X1 U1110 ( .B(n1722), .A(n1723), .S(n1894), .Y(n1721) );
  MUX2X1 U1111 ( .B(n1725), .A(n1726), .S(n1894), .Y(n1724) );
  MUX2X1 U1112 ( .B(n1728), .A(n1729), .S(n1883), .Y(n1727) );
  MUX2X1 U1113 ( .B(n1731), .A(n1732), .S(n1895), .Y(n1730) );
  MUX2X1 U1114 ( .B(n1734), .A(n1735), .S(n1895), .Y(n1733) );
  MUX2X1 U1115 ( .B(n1737), .A(n1738), .S(n1895), .Y(n1736) );
  MUX2X1 U1116 ( .B(n1740), .A(n1741), .S(n1895), .Y(n1739) );
  MUX2X1 U1117 ( .B(n1743), .A(n1744), .S(n1883), .Y(n1742) );
  MUX2X1 U1118 ( .B(n1746), .A(n1747), .S(n1895), .Y(n1745) );
  MUX2X1 U1119 ( .B(n1749), .A(n1750), .S(n1895), .Y(n1748) );
  MUX2X1 U1120 ( .B(n1752), .A(n1753), .S(n1895), .Y(n1751) );
  MUX2X1 U1121 ( .B(n1755), .A(n1756), .S(n1895), .Y(n1754) );
  MUX2X1 U1122 ( .B(n1758), .A(n1759), .S(n1884), .Y(n1757) );
  MUX2X1 U1123 ( .B(n1761), .A(n1762), .S(n1895), .Y(n1760) );
  MUX2X1 U1124 ( .B(n1764), .A(n1765), .S(n1895), .Y(n1763) );
  MUX2X1 U1125 ( .B(n1767), .A(n1768), .S(n1895), .Y(n1766) );
  MUX2X1 U1126 ( .B(n1770), .A(n1771), .S(n1895), .Y(n1769) );
  MUX2X1 U1127 ( .B(n1773), .A(n1774), .S(n1884), .Y(n1772) );
  MUX2X1 U1128 ( .B(n1776), .A(n1777), .S(n1896), .Y(n1775) );
  MUX2X1 U1129 ( .B(n1779), .A(n1780), .S(n1896), .Y(n1778) );
  MUX2X1 U1130 ( .B(n1782), .A(n1783), .S(n1896), .Y(n1781) );
  MUX2X1 U1131 ( .B(n1785), .A(n1786), .S(n1896), .Y(n1784) );
  MUX2X1 U1132 ( .B(n1788), .A(n1789), .S(n1884), .Y(n1787) );
  MUX2X1 U1133 ( .B(n1791), .A(n1792), .S(n1896), .Y(n1790) );
  MUX2X1 U1134 ( .B(n1794), .A(n1795), .S(n1896), .Y(n1793) );
  MUX2X1 U1135 ( .B(n1797), .A(n1798), .S(n1896), .Y(n1796) );
  MUX2X1 U1136 ( .B(n1800), .A(n1801), .S(n1896), .Y(n1799) );
  MUX2X1 U1137 ( .B(n1803), .A(n1804), .S(n2033), .Y(n1802) );
  MUX2X1 U1138 ( .B(n1806), .A(n1807), .S(n1896), .Y(n1805) );
  MUX2X1 U1139 ( .B(n1809), .A(n1810), .S(n1896), .Y(n1808) );
  MUX2X1 U1140 ( .B(n1812), .A(n1813), .S(n1896), .Y(n1811) );
  MUX2X1 U1141 ( .B(n1815), .A(n1816), .S(n1896), .Y(n1814) );
  MUX2X1 U1142 ( .B(n1818), .A(n1819), .S(n1884), .Y(n1817) );
  MUX2X1 U1143 ( .B(n1821), .A(n1822), .S(n1897), .Y(n1820) );
  MUX2X1 U1144 ( .B(n1824), .A(n1825), .S(n1897), .Y(n1823) );
  MUX2X1 U1145 ( .B(n1827), .A(n1828), .S(n1897), .Y(n1826) );
  MUX2X1 U1146 ( .B(n1830), .A(n1831), .S(n1897), .Y(n1829) );
  MUX2X1 U1147 ( .B(n1833), .A(n1834), .S(n2033), .Y(n1832) );
  MUX2X1 U1148 ( .B(n1836), .A(n1837), .S(n1897), .Y(n1835) );
  MUX2X1 U1149 ( .B(n1839), .A(n1840), .S(n1897), .Y(n1838) );
  MUX2X1 U1150 ( .B(n1842), .A(n1843), .S(n1897), .Y(n1841) );
  MUX2X1 U1151 ( .B(n1845), .A(n1846), .S(n1897), .Y(n1844) );
  MUX2X1 U1152 ( .B(n1848), .A(n1849), .S(n2033), .Y(n1847) );
  MUX2X1 U1153 ( .B(n1851), .A(n1852), .S(n1897), .Y(n1850) );
  MUX2X1 U1154 ( .B(n1854), .A(n1855), .S(n1897), .Y(n1853) );
  MUX2X1 U1155 ( .B(n1857), .A(n1858), .S(n1897), .Y(n1856) );
  MUX2X1 U1156 ( .B(n1860), .A(n1861), .S(n1897), .Y(n1859) );
  MUX2X1 U1157 ( .B(n1863), .A(n1864), .S(n2033), .Y(n1862) );
  MUX2X1 U1158 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1905), .Y(n1387) );
  MUX2X1 U1159 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1905), .Y(n1386) );
  MUX2X1 U1160 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1905), .Y(n1390) );
  MUX2X1 U1161 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1905), .Y(n1389) );
  MUX2X1 U1162 ( .B(n1388), .A(n1385), .S(n1886), .Y(n1399) );
  MUX2X1 U1163 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1906), .Y(n1393) );
  MUX2X1 U1164 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1906), .Y(n1392) );
  MUX2X1 U1165 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1906), .Y(n1396) );
  MUX2X1 U1166 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1906), .Y(n1395) );
  MUX2X1 U1167 ( .B(n1394), .A(n1391), .S(n1886), .Y(n1398) );
  MUX2X1 U1168 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1906), .Y(n1402) );
  MUX2X1 U1169 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1906), .Y(n1401) );
  MUX2X1 U1170 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1906), .Y(n1405) );
  MUX2X1 U1171 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1906), .Y(n1404) );
  MUX2X1 U1172 ( .B(n1403), .A(n1400), .S(n1886), .Y(n1414) );
  MUX2X1 U1173 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1906), .Y(n1408) );
  MUX2X1 U1174 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1906), .Y(n1407) );
  MUX2X1 U1175 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1906), .Y(n1411) );
  MUX2X1 U1177 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1906), .Y(n1410) );
  MUX2X1 U1178 ( .B(n1409), .A(n1406), .S(n1886), .Y(n1413) );
  MUX2X1 U1179 ( .B(n1412), .A(n1397), .S(n1882), .Y(n1865) );
  MUX2X1 U1180 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1907), .Y(n1417) );
  MUX2X1 U1181 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1907), .Y(n1416) );
  MUX2X1 U1182 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1907), .Y(n1420) );
  MUX2X1 U1183 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1907), .Y(n1419) );
  MUX2X1 U1184 ( .B(n1418), .A(n1415), .S(n1886), .Y(n1429) );
  MUX2X1 U1185 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1907), .Y(n1423) );
  MUX2X1 U1186 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1907), .Y(n1422) );
  MUX2X1 U1187 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1907), .Y(n1426) );
  MUX2X1 U1188 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1907), .Y(n1425) );
  MUX2X1 U1189 ( .B(n1424), .A(n1421), .S(n1886), .Y(n1428) );
  MUX2X1 U1190 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1907), .Y(n1432) );
  MUX2X1 U1191 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1907), .Y(n1431) );
  MUX2X1 U1192 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1907), .Y(n1435) );
  MUX2X1 U1193 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1907), .Y(n1434) );
  MUX2X1 U1194 ( .B(n1433), .A(n1430), .S(n1886), .Y(n1444) );
  MUX2X1 U1195 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1908), .Y(n1438) );
  MUX2X1 U1196 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1908), .Y(n1437) );
  MUX2X1 U1197 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1908), .Y(n1441) );
  MUX2X1 U1198 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1908), .Y(n1440) );
  MUX2X1 U1199 ( .B(n1439), .A(n1436), .S(n1886), .Y(n1443) );
  MUX2X1 U1200 ( .B(n1442), .A(n1427), .S(n1882), .Y(n1866) );
  MUX2X1 U1201 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1908), .Y(n1447) );
  MUX2X1 U1202 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1908), .Y(n1446) );
  MUX2X1 U1203 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1908), .Y(n1450) );
  MUX2X1 U1204 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1908), .Y(n1449) );
  MUX2X1 U1205 ( .B(n1448), .A(n1445), .S(n1886), .Y(n1459) );
  MUX2X1 U1206 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1908), .Y(n1453) );
  MUX2X1 U1207 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1908), .Y(n1452) );
  MUX2X1 U1208 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1908), .Y(n1456) );
  MUX2X1 U1209 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1908), .Y(n1455) );
  MUX2X1 U1210 ( .B(n1454), .A(n1451), .S(n1886), .Y(n1458) );
  MUX2X1 U1211 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1909), .Y(n1462) );
  MUX2X1 U1212 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1909), .Y(n1461) );
  MUX2X1 U1213 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1909), .Y(n1465) );
  MUX2X1 U1214 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1909), .Y(n1464) );
  MUX2X1 U1215 ( .B(n1463), .A(n1460), .S(n1886), .Y(n1474) );
  MUX2X1 U1216 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1909), .Y(n1468) );
  MUX2X1 U1217 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1909), .Y(n1467) );
  MUX2X1 U1218 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1909), .Y(n1471) );
  MUX2X1 U1219 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1909), .Y(n1470) );
  MUX2X1 U1220 ( .B(n1469), .A(n1466), .S(n1886), .Y(n1473) );
  MUX2X1 U1221 ( .B(n1472), .A(n1457), .S(n1882), .Y(n1867) );
  MUX2X1 U1222 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1909), .Y(n1477) );
  MUX2X1 U1223 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1909), .Y(n1476) );
  MUX2X1 U1224 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1909), .Y(n1480) );
  MUX2X1 U1225 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1909), .Y(n1479) );
  MUX2X1 U1226 ( .B(n1478), .A(n1475), .S(n1885), .Y(n1489) );
  MUX2X1 U1227 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1910), .Y(n1483) );
  MUX2X1 U1228 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1910), .Y(n1482) );
  MUX2X1 U1229 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1910), .Y(n1486) );
  MUX2X1 U1230 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1910), .Y(n1485) );
  MUX2X1 U1231 ( .B(n1484), .A(n1481), .S(n1885), .Y(n1488) );
  MUX2X1 U1232 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1910), .Y(n1492) );
  MUX2X1 U1233 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1910), .Y(n1491) );
  MUX2X1 U1234 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1910), .Y(n1495) );
  MUX2X1 U1235 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1910), .Y(n1494) );
  MUX2X1 U1236 ( .B(n1493), .A(n1490), .S(n1885), .Y(n1504) );
  MUX2X1 U1237 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1910), .Y(n1498) );
  MUX2X1 U1238 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1910), .Y(n1497) );
  MUX2X1 U1239 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1910), .Y(n1501) );
  MUX2X1 U1240 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1910), .Y(n1500) );
  MUX2X1 U1241 ( .B(n1499), .A(n1496), .S(n1885), .Y(n1503) );
  MUX2X1 U1242 ( .B(n1502), .A(n1487), .S(n1882), .Y(n1868) );
  MUX2X1 U1243 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1911), .Y(n1507) );
  MUX2X1 U1244 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1911), .Y(n1506) );
  MUX2X1 U1245 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1911), .Y(n1510) );
  MUX2X1 U1246 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1911), .Y(n1509) );
  MUX2X1 U1247 ( .B(n1508), .A(n1505), .S(n1885), .Y(n1519) );
  MUX2X1 U1248 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1911), .Y(n1513) );
  MUX2X1 U1249 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1911), .Y(n1512) );
  MUX2X1 U1250 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1911), .Y(n1516) );
  MUX2X1 U1251 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1911), .Y(n1515) );
  MUX2X1 U1252 ( .B(n1514), .A(n1511), .S(n1885), .Y(n1518) );
  MUX2X1 U1253 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1911), .Y(n1522) );
  MUX2X1 U1254 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1911), .Y(n1521) );
  MUX2X1 U1255 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1911), .Y(n1525) );
  MUX2X1 U1256 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1911), .Y(n1524) );
  MUX2X1 U1257 ( .B(n1523), .A(n1520), .S(n1885), .Y(n1534) );
  MUX2X1 U1258 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1912), .Y(n1528) );
  MUX2X1 U1259 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1912), .Y(n1527) );
  MUX2X1 U1260 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1912), .Y(n1531) );
  MUX2X1 U1261 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1912), .Y(n1530) );
  MUX2X1 U1262 ( .B(n1529), .A(n1526), .S(n1885), .Y(n1533) );
  MUX2X1 U1263 ( .B(n1532), .A(n1517), .S(n1882), .Y(n1869) );
  MUX2X1 U1264 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1912), .Y(n1537) );
  MUX2X1 U1265 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1912), .Y(n1536) );
  MUX2X1 U1266 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1912), .Y(n1540) );
  MUX2X1 U1267 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1912), .Y(n1539) );
  MUX2X1 U1268 ( .B(n1538), .A(n1535), .S(n1885), .Y(n1549) );
  MUX2X1 U1269 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1912), .Y(n1543) );
  MUX2X1 U1270 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1912), .Y(n1542) );
  MUX2X1 U1271 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1912), .Y(n1546) );
  MUX2X1 U1272 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1912), .Y(n1545) );
  MUX2X1 U1273 ( .B(n1544), .A(n1541), .S(n1885), .Y(n1548) );
  MUX2X1 U1274 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1913), .Y(n1552) );
  MUX2X1 U1275 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1913), .Y(n1551) );
  MUX2X1 U1276 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1913), .Y(n1555) );
  MUX2X1 U1277 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1913), .Y(n1554) );
  MUX2X1 U1278 ( .B(n1553), .A(n1550), .S(n1885), .Y(n1564) );
  MUX2X1 U1279 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1913), .Y(n1558) );
  MUX2X1 U1280 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1913), .Y(n1557) );
  MUX2X1 U1281 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1913), .Y(n1561) );
  MUX2X1 U1282 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1913), .Y(n1560) );
  MUX2X1 U1283 ( .B(n1559), .A(n1556), .S(n1885), .Y(n1563) );
  MUX2X1 U1284 ( .B(n1562), .A(n1547), .S(n1882), .Y(n1870) );
  MUX2X1 U1285 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1913), .Y(n1567) );
  MUX2X1 U1286 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1913), .Y(n1566) );
  MUX2X1 U1287 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1913), .Y(n1570) );
  MUX2X1 U1288 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1913), .Y(n1569) );
  MUX2X1 U1289 ( .B(n1568), .A(n1565), .S(n1886), .Y(n1579) );
  MUX2X1 U1290 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1914), .Y(n1573) );
  MUX2X1 U1291 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1914), .Y(n1572) );
  MUX2X1 U1292 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1914), .Y(n1576) );
  MUX2X1 U1293 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1914), .Y(n1575) );
  MUX2X1 U1294 ( .B(n1574), .A(n1571), .S(n1886), .Y(n1578) );
  MUX2X1 U1295 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1914), .Y(n1582) );
  MUX2X1 U1296 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1914), .Y(n1581) );
  MUX2X1 U1297 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1914), .Y(n1585) );
  MUX2X1 U1298 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1914), .Y(n1584) );
  MUX2X1 U1299 ( .B(n1583), .A(n1580), .S(n1886), .Y(n1594) );
  MUX2X1 U1300 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1914), .Y(n1588) );
  MUX2X1 U1301 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1914), .Y(n1587) );
  MUX2X1 U1302 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1914), .Y(n1591) );
  MUX2X1 U1303 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1914), .Y(n1590) );
  MUX2X1 U1304 ( .B(n1589), .A(n1586), .S(n1886), .Y(n1593) );
  MUX2X1 U1305 ( .B(n1592), .A(n1577), .S(n1882), .Y(n1871) );
  MUX2X1 U1306 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1915), .Y(n1597) );
  MUX2X1 U1307 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1915), .Y(n1596) );
  MUX2X1 U1308 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1915), .Y(n1600) );
  MUX2X1 U1309 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1915), .Y(n1599) );
  MUX2X1 U1310 ( .B(n1598), .A(n1595), .S(n1885), .Y(n1609) );
  MUX2X1 U1311 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1915), .Y(n1603) );
  MUX2X1 U1312 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1915), .Y(n1602) );
  MUX2X1 U1313 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1915), .Y(n1606) );
  MUX2X1 U1314 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1915), .Y(n1605) );
  MUX2X1 U1315 ( .B(n1604), .A(n1601), .S(n1885), .Y(n1608) );
  MUX2X1 U1316 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1915), .Y(n1612) );
  MUX2X1 U1317 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1915), .Y(n1611) );
  MUX2X1 U1318 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1915), .Y(n1615) );
  MUX2X1 U1319 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1915), .Y(n1614) );
  MUX2X1 U1320 ( .B(n1613), .A(n1610), .S(n1885), .Y(n1624) );
  MUX2X1 U1321 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1916), .Y(n1618) );
  MUX2X1 U1322 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1916), .Y(n1617) );
  MUX2X1 U1323 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1916), .Y(n1621) );
  MUX2X1 U1324 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1916), .Y(n1620) );
  MUX2X1 U1325 ( .B(n1619), .A(n1616), .S(n1885), .Y(n1623) );
  MUX2X1 U1326 ( .B(n1622), .A(n1607), .S(n1882), .Y(n1872) );
  MUX2X1 U1327 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1916), .Y(n1627) );
  MUX2X1 U1328 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1916), .Y(n1626) );
  MUX2X1 U1329 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1916), .Y(n1630) );
  MUX2X1 U1330 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1916), .Y(n1629) );
  MUX2X1 U1331 ( .B(n1628), .A(n1625), .S(n1886), .Y(n1639) );
  MUX2X1 U1332 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1916), .Y(n1633) );
  MUX2X1 U1333 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1916), .Y(n1632) );
  MUX2X1 U1334 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1916), .Y(n1636) );
  MUX2X1 U1335 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1916), .Y(n1635) );
  MUX2X1 U1336 ( .B(n1634), .A(n1631), .S(n1886), .Y(n1638) );
  MUX2X1 U1337 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1917), .Y(n1642) );
  MUX2X1 U1338 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1917), .Y(n1641) );
  MUX2X1 U1339 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1917), .Y(n1645) );
  MUX2X1 U1340 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1917), .Y(n1644) );
  MUX2X1 U1341 ( .B(n1643), .A(n1640), .S(n1885), .Y(n1654) );
  MUX2X1 U1342 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1917), .Y(n1648) );
  MUX2X1 U1343 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1917), .Y(n1647) );
  MUX2X1 U1344 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1917), .Y(n1651) );
  MUX2X1 U1345 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1917), .Y(n1650) );
  MUX2X1 U1346 ( .B(n1649), .A(n1646), .S(n1886), .Y(n1653) );
  MUX2X1 U1347 ( .B(n1652), .A(n1637), .S(n1882), .Y(n1873) );
  MUX2X1 U1348 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1917), .Y(n1657) );
  MUX2X1 U1349 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1917), .Y(n1656) );
  MUX2X1 U1350 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1917), .Y(n1660) );
  MUX2X1 U1351 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1917), .Y(n1659) );
  MUX2X1 U1352 ( .B(n1658), .A(n1655), .S(n1885), .Y(n1669) );
  MUX2X1 U1353 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1918), .Y(n1663) );
  MUX2X1 U1354 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1918), .Y(n1662) );
  MUX2X1 U1355 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1918), .Y(n1666) );
  MUX2X1 U1356 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1918), .Y(n1665) );
  MUX2X1 U1357 ( .B(n1664), .A(n1661), .S(n1885), .Y(n1668) );
  MUX2X1 U1358 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1918), .Y(n1672) );
  MUX2X1 U1359 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1918), .Y(n1671) );
  MUX2X1 U1360 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1918), .Y(n1675) );
  MUX2X1 U1361 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1918), .Y(n1674) );
  MUX2X1 U1362 ( .B(n1673), .A(n1670), .S(n1885), .Y(n1684) );
  MUX2X1 U1363 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1918), .Y(n1678) );
  MUX2X1 U1364 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1918), .Y(n1677) );
  MUX2X1 U1365 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1918), .Y(n1681) );
  MUX2X1 U1366 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1918), .Y(n1680) );
  MUX2X1 U1367 ( .B(n1679), .A(n1676), .S(n1885), .Y(n1683) );
  MUX2X1 U1368 ( .B(n1682), .A(n1667), .S(n1882), .Y(n1874) );
  MUX2X1 U1369 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1919), .Y(n1687) );
  MUX2X1 U1370 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1919), .Y(n1686) );
  MUX2X1 U1371 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1919), .Y(n1690) );
  MUX2X1 U1372 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1919), .Y(n1689) );
  MUX2X1 U1373 ( .B(n1688), .A(n1685), .S(n1885), .Y(n1699) );
  MUX2X1 U1374 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1919), .Y(n1693) );
  MUX2X1 U1375 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1919), .Y(n1692) );
  MUX2X1 U1376 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1919), .Y(n1696) );
  MUX2X1 U1377 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1919), .Y(n1695) );
  MUX2X1 U1378 ( .B(n1694), .A(n1691), .S(n1885), .Y(n1698) );
  MUX2X1 U1379 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1919), .Y(n1702) );
  MUX2X1 U1380 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1919), .Y(n1701) );
  MUX2X1 U1381 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1919), .Y(n1705) );
  MUX2X1 U1382 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1919), .Y(n1704) );
  MUX2X1 U1383 ( .B(n1703), .A(n1700), .S(n1885), .Y(n1714) );
  MUX2X1 U1384 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1920), .Y(n1708) );
  MUX2X1 U1385 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1920), .Y(n1707) );
  MUX2X1 U1386 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1920), .Y(n1711) );
  MUX2X1 U1387 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1920), .Y(n1710) );
  MUX2X1 U1388 ( .B(n1709), .A(n1706), .S(n1885), .Y(n1713) );
  MUX2X1 U1389 ( .B(n1712), .A(n1697), .S(n1882), .Y(n1875) );
  MUX2X1 U1390 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1920), .Y(n1717) );
  MUX2X1 U1391 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1920), .Y(n1716) );
  MUX2X1 U1392 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1920), .Y(n1720) );
  MUX2X1 U1393 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1920), .Y(n1719) );
  MUX2X1 U1394 ( .B(n1718), .A(n1715), .S(n1885), .Y(n1729) );
  MUX2X1 U1395 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1920), .Y(n1723) );
  MUX2X1 U1396 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1920), .Y(n1722) );
  MUX2X1 U1397 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1920), .Y(n1726) );
  MUX2X1 U1398 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1920), .Y(n1725) );
  MUX2X1 U1399 ( .B(n1724), .A(n1721), .S(n1885), .Y(n1728) );
  MUX2X1 U1400 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1921), .Y(n1732) );
  MUX2X1 U1401 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1921), .Y(n1731) );
  MUX2X1 U1402 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1921), .Y(n1735) );
  MUX2X1 U1403 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1921), .Y(n1734) );
  MUX2X1 U1404 ( .B(n1733), .A(n1730), .S(n1885), .Y(n1744) );
  MUX2X1 U1405 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1921), .Y(n1738) );
  MUX2X1 U1406 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1921), .Y(n1737) );
  MUX2X1 U1407 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1921), .Y(n1741) );
  MUX2X1 U1408 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1921), .Y(n1740) );
  MUX2X1 U1409 ( .B(n1739), .A(n1736), .S(n1885), .Y(n1743) );
  MUX2X1 U1410 ( .B(n1742), .A(n1727), .S(n1882), .Y(n1876) );
  MUX2X1 U1411 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1921), .Y(n1747) );
  MUX2X1 U1412 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1921), .Y(n1746) );
  MUX2X1 U1413 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1921), .Y(n1750) );
  MUX2X1 U1414 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1921), .Y(n1749) );
  MUX2X1 U1415 ( .B(n1748), .A(n1745), .S(n1886), .Y(n1759) );
  MUX2X1 U1416 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1922), .Y(n1753) );
  MUX2X1 U1417 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1922), .Y(n1752) );
  MUX2X1 U1418 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1922), .Y(n1756) );
  MUX2X1 U1419 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1922), .Y(n1755) );
  MUX2X1 U1420 ( .B(n1754), .A(n1751), .S(n2031), .Y(n1758) );
  MUX2X1 U1421 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1922), .Y(n1762) );
  MUX2X1 U1422 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1922), .Y(n1761) );
  MUX2X1 U1423 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1922), .Y(n1765) );
  MUX2X1 U1424 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1922), .Y(n1764) );
  MUX2X1 U1425 ( .B(n1763), .A(n1760), .S(n1886), .Y(n1774) );
  MUX2X1 U1426 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1922), .Y(n1768) );
  MUX2X1 U1427 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1922), .Y(n1767) );
  MUX2X1 U1428 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1922), .Y(n1771) );
  MUX2X1 U1429 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1922), .Y(n1770) );
  MUX2X1 U1430 ( .B(n1769), .A(n1766), .S(n1886), .Y(n1773) );
  MUX2X1 U1431 ( .B(n1772), .A(n1757), .S(n1881), .Y(n1877) );
  MUX2X1 U1432 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1923), .Y(n1777) );
  MUX2X1 U1433 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1923), .Y(n1776) );
  MUX2X1 U1434 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1923), .Y(n1780) );
  MUX2X1 U1435 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1923), .Y(n1779) );
  MUX2X1 U1436 ( .B(n1778), .A(n1775), .S(n1886), .Y(n1789) );
  MUX2X1 U1437 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1923), .Y(n1783) );
  MUX2X1 U1438 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1923), .Y(n1782) );
  MUX2X1 U1439 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1923), .Y(n1786) );
  MUX2X1 U1440 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1923), .Y(n1785) );
  MUX2X1 U1441 ( .B(n1784), .A(n1781), .S(n1886), .Y(n1788) );
  MUX2X1 U1442 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1923), .Y(n1792) );
  MUX2X1 U1443 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1923), .Y(n1791) );
  MUX2X1 U1444 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1923), .Y(n1795) );
  MUX2X1 U1445 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1923), .Y(n1794) );
  MUX2X1 U1446 ( .B(n1793), .A(n1790), .S(n2031), .Y(n1804) );
  MUX2X1 U1447 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1924), .Y(n1798) );
  MUX2X1 U1448 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1924), .Y(n1797) );
  MUX2X1 U1449 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1924), .Y(n1801) );
  MUX2X1 U1450 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1924), .Y(n1800) );
  MUX2X1 U1451 ( .B(n1799), .A(n1796), .S(n1886), .Y(n1803) );
  MUX2X1 U1452 ( .B(n1802), .A(n1787), .S(n1881), .Y(n1878) );
  MUX2X1 U1453 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1924), .Y(n1807) );
  MUX2X1 U1454 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1924), .Y(n1806) );
  MUX2X1 U1455 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1924), .Y(n1810) );
  MUX2X1 U1456 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1924), .Y(n1809) );
  MUX2X1 U1457 ( .B(n1808), .A(n1805), .S(n1886), .Y(n1819) );
  MUX2X1 U1458 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1924), .Y(n1813) );
  MUX2X1 U1459 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1924), .Y(n1812) );
  MUX2X1 U1460 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1924), .Y(n1816) );
  MUX2X1 U1461 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1924), .Y(n1815) );
  MUX2X1 U1462 ( .B(n1814), .A(n1811), .S(n1886), .Y(n1818) );
  MUX2X1 U1463 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1925), .Y(n1822) );
  MUX2X1 U1464 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1925), .Y(n1821) );
  MUX2X1 U1465 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1925), .Y(n1825) );
  MUX2X1 U1466 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1925), .Y(n1824) );
  MUX2X1 U1467 ( .B(n1823), .A(n1820), .S(n2031), .Y(n1834) );
  MUX2X1 U1468 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1925), .Y(n1828) );
  MUX2X1 U1469 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1925), .Y(n1827) );
  MUX2X1 U1470 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1925), .Y(n1831) );
  MUX2X1 U1471 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1925), .Y(n1830) );
  MUX2X1 U1472 ( .B(n1829), .A(n1826), .S(n1886), .Y(n1833) );
  MUX2X1 U1473 ( .B(n1832), .A(n1817), .S(n1881), .Y(n1879) );
  MUX2X1 U1474 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1925), .Y(n1837) );
  MUX2X1 U1475 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1925), .Y(n1836) );
  MUX2X1 U1476 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1925), .Y(n1840) );
  MUX2X1 U1477 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1925), .Y(n1839) );
  MUX2X1 U1478 ( .B(n1838), .A(n1835), .S(n1886), .Y(n1849) );
  MUX2X1 U1479 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1926), .Y(n1843) );
  MUX2X1 U1480 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1926), .Y(n1842) );
  MUX2X1 U1481 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1926), .Y(n1846) );
  MUX2X1 U1482 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1926), .Y(n1845) );
  MUX2X1 U1483 ( .B(n1844), .A(n1841), .S(n1886), .Y(n1848) );
  MUX2X1 U1484 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1926), .Y(n1852) );
  MUX2X1 U1485 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1926), .Y(n1851) );
  MUX2X1 U1486 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1926), .Y(n1855) );
  MUX2X1 U1487 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1926), .Y(n1854) );
  MUX2X1 U1488 ( .B(n1853), .A(n1850), .S(n2031), .Y(n1864) );
  MUX2X1 U1489 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1926), .Y(n1858) );
  MUX2X1 U1490 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1926), .Y(n1857) );
  MUX2X1 U1491 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1926), .Y(n1861) );
  MUX2X1 U1492 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1926), .Y(n1860) );
  MUX2X1 U1493 ( .B(n1859), .A(n1856), .S(n2031), .Y(n1863) );
  MUX2X1 U1494 ( .B(n1862), .A(n1847), .S(n1881), .Y(n1880) );
  INVX8 U1495 ( .A(n2032), .Y(n1885) );
  INVX8 U1496 ( .A(n2032), .Y(n1886) );
  INVX8 U1497 ( .A(n1929), .Y(n1900) );
  INVX8 U1498 ( .A(n1929), .Y(n1901) );
  INVX8 U1499 ( .A(n1930), .Y(n1902) );
  INVX8 U1500 ( .A(n1930), .Y(n1903) );
  INVX8 U1501 ( .A(n1930), .Y(n1904) );
  INVX8 U1502 ( .A(n1904), .Y(n1905) );
  INVX8 U1503 ( .A(n1904), .Y(n1906) );
  INVX8 U1504 ( .A(n1904), .Y(n1907) );
  INVX8 U1505 ( .A(n1903), .Y(n1908) );
  INVX8 U1506 ( .A(n1903), .Y(n1909) );
  INVX8 U1507 ( .A(n1903), .Y(n1910) );
  INVX8 U1508 ( .A(n1902), .Y(n1911) );
  INVX8 U1509 ( .A(n1902), .Y(n1912) );
  INVX8 U1510 ( .A(n1902), .Y(n1913) );
  INVX8 U1511 ( .A(n1901), .Y(n1914) );
  INVX8 U1512 ( .A(n1901), .Y(n1915) );
  INVX8 U1513 ( .A(n1901), .Y(n1916) );
  INVX8 U1514 ( .A(n1927), .Y(n1917) );
  INVX8 U1515 ( .A(n1903), .Y(n1918) );
  INVX8 U1516 ( .A(n1927), .Y(n1919) );
  INVX8 U1517 ( .A(n1900), .Y(n1920) );
  INVX8 U1518 ( .A(n1900), .Y(n1921) );
  INVX8 U1519 ( .A(n1900), .Y(n1922) );
  INVX8 U1520 ( .A(n1899), .Y(n1923) );
  INVX8 U1521 ( .A(n1899), .Y(n1924) );
  INVX8 U1522 ( .A(n1899), .Y(n1925) );
  INVX8 U1523 ( .A(n1899), .Y(n1926) );
  INVX8 U1524 ( .A(n1927), .Y(n1929) );
  INVX8 U1525 ( .A(n1927), .Y(n1930) );
  INVX1 U1526 ( .A(n1384), .Y(n1931) );
  AND2X2 U1527 ( .A(N20), .B(n3), .Y(\data_out<12> ) );
  INVX1 U1528 ( .A(N11), .Y(n2030) );
  INVX1 U1529 ( .A(N10), .Y(n2029) );
  INVX8 U1530 ( .A(n1995), .Y(n1992) );
  INVX8 U1531 ( .A(n1995), .Y(n1993) );
  INVX8 U1532 ( .A(n106), .Y(n1995) );
  INVX8 U1533 ( .A(n92), .Y(n1997) );
  INVX8 U1534 ( .A(n93), .Y(n1999) );
  INVX8 U1535 ( .A(n94), .Y(n2001) );
  INVX8 U1536 ( .A(n95), .Y(n2003) );
  INVX8 U1537 ( .A(n96), .Y(n2005) );
  INVX8 U1538 ( .A(n97), .Y(n2007) );
  INVX8 U1539 ( .A(n98), .Y(n2009) );
  INVX8 U1540 ( .A(n99), .Y(n2011) );
  INVX8 U1541 ( .A(n100), .Y(n2013) );
  INVX8 U1542 ( .A(n101), .Y(n2015) );
  INVX8 U1543 ( .A(n107), .Y(n2017) );
  INVX8 U1544 ( .A(n107), .Y(n2018) );
  INVX8 U1545 ( .A(n108), .Y(n2019) );
  INVX8 U1546 ( .A(n108), .Y(n2020) );
  INVX8 U1547 ( .A(n109), .Y(n2021) );
  INVX8 U1548 ( .A(n109), .Y(n2022) );
  INVX8 U1549 ( .A(n110), .Y(n2023) );
  INVX8 U1550 ( .A(n110), .Y(n2024) );
  AND2X2 U1551 ( .A(n111), .B(n112), .Y(\data_out<0> ) );
  AND2X2 U1552 ( .A(N31), .B(n1383), .Y(\data_out<1> ) );
  AND2X2 U1553 ( .A(N30), .B(n3), .Y(\data_out<2> ) );
  AND2X2 U1554 ( .A(n1383), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U1555 ( .A(n111), .B(n156), .Y(\data_out<4> ) );
  AND2X2 U1556 ( .A(n1383), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U1557 ( .A(n1383), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U1558 ( .A(n1381), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U1559 ( .A(N23), .B(n3), .Y(\data_out<9> ) );
  AND2X2 U1560 ( .A(n111), .B(n1382), .Y(\data_out<10> ) );
  AND2X2 U1561 ( .A(n1383), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U1562 ( .A(n1931), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U1563 ( .A(n1931), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U1564 ( .A(n1381), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U1565 ( .A(\mem<31><0> ), .B(n125), .Y(n2037) );
  OAI21X1 U1566 ( .A(n1933), .B(n1996), .C(n2037), .Y(n2743) );
  OAI21X1 U1567 ( .A(n1998), .B(n1932), .C(n158), .Y(n2742) );
  OAI21X1 U1568 ( .A(n2000), .B(n1932), .C(n160), .Y(n2741) );
  OAI21X1 U1569 ( .A(n2002), .B(n1932), .C(n162), .Y(n2740) );
  OAI21X1 U1570 ( .A(n2004), .B(n1932), .C(n164), .Y(n2739) );
  OAI21X1 U1571 ( .A(n2006), .B(n1932), .C(n166), .Y(n2738) );
  OAI21X1 U1572 ( .A(n2008), .B(n1932), .C(n168), .Y(n2737) );
  OAI21X1 U1573 ( .A(n2010), .B(n1932), .C(n170), .Y(n2736) );
  OAI21X1 U1574 ( .A(n2012), .B(n1932), .C(n172), .Y(n2735) );
  OAI21X1 U1575 ( .A(n2014), .B(n1933), .C(n174), .Y(n2734) );
  OAI21X1 U1576 ( .A(n2016), .B(n1933), .C(n176), .Y(n2733) );
  OAI21X1 U1577 ( .A(n2018), .B(n1933), .C(n178), .Y(n2732) );
  OAI21X1 U1578 ( .A(n2020), .B(n1933), .C(n180), .Y(n2731) );
  OAI21X1 U1579 ( .A(n2022), .B(n1933), .C(n182), .Y(n2730) );
  OAI21X1 U1580 ( .A(n2024), .B(n1933), .C(n184), .Y(n2729) );
  NAND2X1 U1581 ( .A(\mem<31><15> ), .B(n140), .Y(n2038) );
  OAI21X1 U1582 ( .A(n1366), .B(n1933), .C(n2038), .Y(n2728) );
  NAND2X1 U1583 ( .A(\mem<30><0> ), .B(n143), .Y(n2039) );
  OAI21X1 U1584 ( .A(n1934), .B(n1996), .C(n2039), .Y(n2727) );
  OAI21X1 U1585 ( .A(n1934), .B(n1998), .C(n186), .Y(n2726) );
  OAI21X1 U1586 ( .A(n1934), .B(n2000), .C(n188), .Y(n2725) );
  OAI21X1 U1587 ( .A(n1934), .B(n2002), .C(n190), .Y(n2724) );
  OAI21X1 U1588 ( .A(n1934), .B(n2004), .C(n192), .Y(n2723) );
  OAI21X1 U1589 ( .A(n1934), .B(n2006), .C(n194), .Y(n2722) );
  OAI21X1 U1590 ( .A(n1934), .B(n2008), .C(n196), .Y(n2721) );
  OAI21X1 U1591 ( .A(n1934), .B(n2010), .C(n198), .Y(n2720) );
  OAI21X1 U1592 ( .A(n1935), .B(n2012), .C(n200), .Y(n2719) );
  OAI21X1 U1593 ( .A(n1935), .B(n2014), .C(n202), .Y(n2718) );
  OAI21X1 U1594 ( .A(n1935), .B(n2016), .C(n204), .Y(n2717) );
  OAI21X1 U1595 ( .A(n1935), .B(n2017), .C(n206), .Y(n2716) );
  OAI21X1 U1596 ( .A(n1935), .B(n2019), .C(n208), .Y(n2715) );
  OAI21X1 U1597 ( .A(n1935), .B(n2021), .C(n210), .Y(n2714) );
  OAI21X1 U1598 ( .A(n1935), .B(n2023), .C(n212), .Y(n2713) );
  OAI21X1 U1599 ( .A(n1935), .B(n1372), .C(n2), .Y(n2712) );
  NAND3X1 U1600 ( .A(n2028), .B(n2031), .C(n2030), .Y(n2040) );
  NAND2X1 U1601 ( .A(\mem<29><0> ), .B(n145), .Y(n2041) );
  OAI21X1 U1602 ( .A(n1936), .B(n1996), .C(n2041), .Y(n2711) );
  OAI21X1 U1603 ( .A(n1936), .B(n1998), .C(n215), .Y(n2710) );
  OAI21X1 U1604 ( .A(n1936), .B(n2000), .C(n217), .Y(n2709) );
  OAI21X1 U1605 ( .A(n1936), .B(n2002), .C(n219), .Y(n2708) );
  OAI21X1 U1606 ( .A(n1936), .B(n2004), .C(n221), .Y(n2707) );
  OAI21X1 U1607 ( .A(n1936), .B(n2006), .C(n223), .Y(n2706) );
  OAI21X1 U1608 ( .A(n1936), .B(n2008), .C(n225), .Y(n2705) );
  OAI21X1 U1609 ( .A(n1936), .B(n2010), .C(n227), .Y(n2704) );
  OAI21X1 U1610 ( .A(n1937), .B(n2012), .C(n229), .Y(n2703) );
  OAI21X1 U1611 ( .A(n1937), .B(n2014), .C(n231), .Y(n2702) );
  OAI21X1 U1612 ( .A(n1937), .B(n2016), .C(n233), .Y(n2701) );
  OAI21X1 U1613 ( .A(n1937), .B(n2018), .C(n235), .Y(n2700) );
  OAI21X1 U1614 ( .A(n1937), .B(n2020), .C(n237), .Y(n2699) );
  OAI21X1 U1615 ( .A(n1937), .B(n2022), .C(n239), .Y(n2698) );
  OAI21X1 U1616 ( .A(n1937), .B(n2024), .C(n241), .Y(n2697) );
  OAI21X1 U1617 ( .A(n1937), .B(n1373), .C(n115), .Y(n2696) );
  NAND3X1 U1618 ( .A(n2031), .B(n2030), .C(n2029), .Y(n2042) );
  NAND2X1 U1619 ( .A(\mem<28><0> ), .B(n147), .Y(n2043) );
  OAI21X1 U1620 ( .A(n1938), .B(n1996), .C(n2043), .Y(n2695) );
  OAI21X1 U1621 ( .A(n1938), .B(n1998), .C(n243), .Y(n2694) );
  OAI21X1 U1622 ( .A(n1938), .B(n2000), .C(n245), .Y(n2693) );
  OAI21X1 U1623 ( .A(n1938), .B(n2002), .C(n247), .Y(n2692) );
  OAI21X1 U1624 ( .A(n1938), .B(n2004), .C(n249), .Y(n2691) );
  OAI21X1 U1625 ( .A(n1938), .B(n2006), .C(n251), .Y(n2690) );
  OAI21X1 U1626 ( .A(n1938), .B(n2008), .C(n253), .Y(n2689) );
  OAI21X1 U1627 ( .A(n1938), .B(n2010), .C(n255), .Y(n2688) );
  OAI21X1 U1628 ( .A(n1939), .B(n2012), .C(n257), .Y(n2687) );
  OAI21X1 U1629 ( .A(n1939), .B(n2014), .C(n259), .Y(n2686) );
  OAI21X1 U1630 ( .A(n1939), .B(n2016), .C(n261), .Y(n2685) );
  OAI21X1 U1631 ( .A(n1939), .B(n2017), .C(n263), .Y(n2684) );
  OAI21X1 U1632 ( .A(n1939), .B(n2019), .C(n265), .Y(n2683) );
  OAI21X1 U1633 ( .A(n1939), .B(n2021), .C(n267), .Y(n2682) );
  OAI21X1 U1634 ( .A(n1939), .B(n2023), .C(n269), .Y(n2681) );
  OAI21X1 U1635 ( .A(n1939), .B(n1374), .C(n117), .Y(n2680) );
  NAND3X1 U1636 ( .A(n2028), .B(n1895), .C(n2032), .Y(n2044) );
  NAND2X1 U1637 ( .A(\mem<27><0> ), .B(n149), .Y(n2045) );
  OAI21X1 U1638 ( .A(n1940), .B(n1996), .C(n2045), .Y(n2679) );
  OAI21X1 U1639 ( .A(n1940), .B(n1998), .C(n271), .Y(n2678) );
  OAI21X1 U1640 ( .A(n1940), .B(n2000), .C(n273), .Y(n2677) );
  OAI21X1 U1641 ( .A(n1940), .B(n2002), .C(n275), .Y(n2676) );
  OAI21X1 U1642 ( .A(n1940), .B(n2004), .C(n277), .Y(n2675) );
  OAI21X1 U1643 ( .A(n1940), .B(n2006), .C(n279), .Y(n2674) );
  OAI21X1 U1644 ( .A(n1940), .B(n2008), .C(n281), .Y(n2673) );
  OAI21X1 U1645 ( .A(n1940), .B(n2010), .C(n283), .Y(n2672) );
  OAI21X1 U1646 ( .A(n1941), .B(n2012), .C(n285), .Y(n2671) );
  OAI21X1 U1647 ( .A(n1941), .B(n2014), .C(n287), .Y(n2670) );
  OAI21X1 U1648 ( .A(n1941), .B(n2016), .C(n289), .Y(n2669) );
  OAI21X1 U1649 ( .A(n1941), .B(n2018), .C(n291), .Y(n2668) );
  OAI21X1 U1650 ( .A(n1941), .B(n2020), .C(n293), .Y(n2667) );
  OAI21X1 U1651 ( .A(n1941), .B(n2022), .C(n295), .Y(n2666) );
  OAI21X1 U1652 ( .A(n1941), .B(n2024), .C(n297), .Y(n2665) );
  OAI21X1 U1653 ( .A(n1941), .B(n1380), .C(n119), .Y(n2664) );
  NAND3X1 U1654 ( .A(n2032), .B(n1891), .C(n2029), .Y(n2046) );
  NAND2X1 U1655 ( .A(\mem<26><0> ), .B(n151), .Y(n2047) );
  OAI21X1 U1656 ( .A(n1942), .B(n1996), .C(n2047), .Y(n2663) );
  OAI21X1 U1657 ( .A(n1942), .B(n1998), .C(n299), .Y(n2662) );
  OAI21X1 U1658 ( .A(n1942), .B(n2000), .C(n301), .Y(n2661) );
  OAI21X1 U1659 ( .A(n1942), .B(n2002), .C(n303), .Y(n2660) );
  OAI21X1 U1660 ( .A(n1942), .B(n2004), .C(n305), .Y(n2659) );
  OAI21X1 U1661 ( .A(n1942), .B(n2006), .C(n307), .Y(n2658) );
  OAI21X1 U1662 ( .A(n1942), .B(n2008), .C(n309), .Y(n2657) );
  OAI21X1 U1663 ( .A(n1942), .B(n2010), .C(n311), .Y(n2656) );
  OAI21X1 U1664 ( .A(n1943), .B(n2012), .C(n313), .Y(n2655) );
  OAI21X1 U1665 ( .A(n1943), .B(n2014), .C(n315), .Y(n2654) );
  OAI21X1 U1666 ( .A(n1943), .B(n2016), .C(n317), .Y(n2653) );
  OAI21X1 U1667 ( .A(n1943), .B(n2017), .C(n319), .Y(n2652) );
  OAI21X1 U1668 ( .A(n1943), .B(n2019), .C(n321), .Y(n2651) );
  OAI21X1 U1669 ( .A(n1943), .B(n2021), .C(n323), .Y(n2650) );
  OAI21X1 U1670 ( .A(n1943), .B(n2023), .C(n325), .Y(n2649) );
  OAI21X1 U1671 ( .A(n1943), .B(n1367), .C(n121), .Y(n2648) );
  NAND3X1 U1672 ( .A(n2028), .B(n2032), .C(n2030), .Y(n2048) );
  NAND2X1 U1673 ( .A(\mem<25><0> ), .B(n153), .Y(n2049) );
  OAI21X1 U1674 ( .A(n1944), .B(n1996), .C(n2049), .Y(n2647) );
  OAI21X1 U1675 ( .A(n1944), .B(n1998), .C(n327), .Y(n2646) );
  OAI21X1 U1676 ( .A(n1944), .B(n2000), .C(n329), .Y(n2645) );
  OAI21X1 U1677 ( .A(n1944), .B(n2002), .C(n331), .Y(n2644) );
  OAI21X1 U1678 ( .A(n1944), .B(n2004), .C(n333), .Y(n2643) );
  OAI21X1 U1679 ( .A(n1944), .B(n2006), .C(n335), .Y(n2642) );
  OAI21X1 U1680 ( .A(n1944), .B(n2008), .C(n337), .Y(n2641) );
  OAI21X1 U1681 ( .A(n1944), .B(n2010), .C(n339), .Y(n2640) );
  OAI21X1 U1682 ( .A(n1945), .B(n2012), .C(n341), .Y(n2639) );
  OAI21X1 U1683 ( .A(n1945), .B(n2014), .C(n343), .Y(n2638) );
  OAI21X1 U1684 ( .A(n1945), .B(n2016), .C(n345), .Y(n2637) );
  OAI21X1 U1685 ( .A(n1945), .B(n2018), .C(n347), .Y(n2636) );
  OAI21X1 U1686 ( .A(n1945), .B(n2020), .C(n349), .Y(n2635) );
  OAI21X1 U1687 ( .A(n1945), .B(n2022), .C(n351), .Y(n2634) );
  OAI21X1 U1688 ( .A(n1945), .B(n2024), .C(n353), .Y(n2633) );
  OAI21X1 U1689 ( .A(n1945), .B(n1366), .C(n123), .Y(n2632) );
  NOR3X1 U1690 ( .A(n2028), .B(n1895), .C(n2031), .Y(n2222) );
  NAND2X1 U1691 ( .A(\mem<24><0> ), .B(n154), .Y(n2050) );
  OAI21X1 U1692 ( .A(n1946), .B(n1996), .C(n2050), .Y(n2631) );
  OAI21X1 U1693 ( .A(n1946), .B(n1998), .C(n355), .Y(n2630) );
  OAI21X1 U1694 ( .A(n1946), .B(n2000), .C(n357), .Y(n2629) );
  OAI21X1 U1695 ( .A(n1946), .B(n2002), .C(n359), .Y(n2628) );
  OAI21X1 U1696 ( .A(n1946), .B(n2004), .C(n361), .Y(n2627) );
  OAI21X1 U1697 ( .A(n1946), .B(n2006), .C(n363), .Y(n2626) );
  OAI21X1 U1698 ( .A(n1946), .B(n2008), .C(n365), .Y(n2625) );
  OAI21X1 U1699 ( .A(n1946), .B(n2010), .C(n367), .Y(n2624) );
  OAI21X1 U1700 ( .A(n1946), .B(n2012), .C(n369), .Y(n2623) );
  OAI21X1 U1701 ( .A(n1946), .B(n2014), .C(n371), .Y(n2622) );
  OAI21X1 U1702 ( .A(n1946), .B(n2016), .C(n373), .Y(n2621) );
  OAI21X1 U1703 ( .A(n1946), .B(n2017), .C(n375), .Y(n2620) );
  OAI21X1 U1704 ( .A(n1946), .B(n2019), .C(n377), .Y(n2619) );
  OAI21X1 U1705 ( .A(n1946), .B(n2021), .C(n379), .Y(n2618) );
  OAI21X1 U1706 ( .A(n1946), .B(n2023), .C(n381), .Y(n2617) );
  NAND2X1 U1707 ( .A(\mem<24><15> ), .B(n139), .Y(n2051) );
  OAI21X1 U1708 ( .A(n1946), .B(n1365), .C(n2051), .Y(n2616) );
  NAND2X1 U1709 ( .A(\mem<23><0> ), .B(n5), .Y(n2052) );
  OAI21X1 U1710 ( .A(n1947), .B(n1996), .C(n2052), .Y(n2615) );
  NAND2X1 U1711 ( .A(\mem<23><1> ), .B(n5), .Y(n2053) );
  OAI21X1 U1712 ( .A(n1947), .B(n1997), .C(n2053), .Y(n2614) );
  NAND2X1 U1713 ( .A(\mem<23><2> ), .B(n5), .Y(n2054) );
  OAI21X1 U1714 ( .A(n1947), .B(n1999), .C(n2054), .Y(n2613) );
  NAND2X1 U1715 ( .A(\mem<23><3> ), .B(n5), .Y(n2055) );
  OAI21X1 U1716 ( .A(n1947), .B(n2001), .C(n2055), .Y(n2612) );
  NAND2X1 U1717 ( .A(\mem<23><4> ), .B(n5), .Y(n2056) );
  OAI21X1 U1718 ( .A(n1947), .B(n2003), .C(n2056), .Y(n2611) );
  NAND2X1 U1719 ( .A(\mem<23><5> ), .B(n5), .Y(n2057) );
  OAI21X1 U1720 ( .A(n1947), .B(n2005), .C(n2057), .Y(n2610) );
  NAND2X1 U1721 ( .A(\mem<23><6> ), .B(n5), .Y(n2058) );
  OAI21X1 U1722 ( .A(n1947), .B(n2007), .C(n2058), .Y(n2609) );
  NAND2X1 U1723 ( .A(\mem<23><7> ), .B(n5), .Y(n2059) );
  OAI21X1 U1724 ( .A(n1947), .B(n2009), .C(n2059), .Y(n2608) );
  NAND2X1 U1725 ( .A(\mem<23><8> ), .B(n5), .Y(n2060) );
  OAI21X1 U1726 ( .A(n1948), .B(n2011), .C(n2060), .Y(n2607) );
  NAND2X1 U1727 ( .A(\mem<23><9> ), .B(n5), .Y(n2061) );
  OAI21X1 U1728 ( .A(n1948), .B(n2013), .C(n2061), .Y(n2606) );
  NAND2X1 U1729 ( .A(\mem<23><10> ), .B(n5), .Y(n2062) );
  OAI21X1 U1730 ( .A(n1948), .B(n2015), .C(n2062), .Y(n2605) );
  NAND2X1 U1731 ( .A(\mem<23><11> ), .B(n5), .Y(n2063) );
  OAI21X1 U1732 ( .A(n1948), .B(n2018), .C(n2063), .Y(n2604) );
  NAND2X1 U1733 ( .A(\mem<23><12> ), .B(n5), .Y(n2064) );
  OAI21X1 U1734 ( .A(n1948), .B(n2020), .C(n2064), .Y(n2603) );
  NAND2X1 U1735 ( .A(\mem<23><13> ), .B(n5), .Y(n2065) );
  OAI21X1 U1736 ( .A(n1948), .B(n2022), .C(n2065), .Y(n2602) );
  NAND2X1 U1737 ( .A(\mem<23><14> ), .B(n5), .Y(n2066) );
  OAI21X1 U1738 ( .A(n1948), .B(n2024), .C(n2066), .Y(n2601) );
  NAND2X1 U1739 ( .A(\mem<23><15> ), .B(n5), .Y(n2067) );
  OAI21X1 U1740 ( .A(n1948), .B(n1376), .C(n2067), .Y(n2600) );
  NAND2X1 U1741 ( .A(\mem<22><0> ), .B(n7), .Y(n2068) );
  OAI21X1 U1742 ( .A(n1949), .B(n1996), .C(n2068), .Y(n2599) );
  NAND2X1 U1743 ( .A(\mem<22><1> ), .B(n7), .Y(n2069) );
  OAI21X1 U1744 ( .A(n1949), .B(n1997), .C(n2069), .Y(n2598) );
  NAND2X1 U1745 ( .A(\mem<22><2> ), .B(n7), .Y(n2070) );
  OAI21X1 U1746 ( .A(n1949), .B(n1999), .C(n2070), .Y(n2597) );
  NAND2X1 U1747 ( .A(\mem<22><3> ), .B(n7), .Y(n2071) );
  OAI21X1 U1748 ( .A(n1949), .B(n2001), .C(n2071), .Y(n2596) );
  NAND2X1 U1749 ( .A(\mem<22><4> ), .B(n7), .Y(n2072) );
  OAI21X1 U1750 ( .A(n1949), .B(n2003), .C(n2072), .Y(n2595) );
  NAND2X1 U1751 ( .A(\mem<22><5> ), .B(n7), .Y(n2073) );
  OAI21X1 U1752 ( .A(n1949), .B(n2005), .C(n2073), .Y(n2594) );
  NAND2X1 U1753 ( .A(\mem<22><6> ), .B(n7), .Y(n2074) );
  OAI21X1 U1754 ( .A(n1949), .B(n2007), .C(n2074), .Y(n2593) );
  NAND2X1 U1755 ( .A(\mem<22><7> ), .B(n7), .Y(n2075) );
  OAI21X1 U1756 ( .A(n1949), .B(n2009), .C(n2075), .Y(n2592) );
  NAND2X1 U1757 ( .A(\mem<22><8> ), .B(n7), .Y(n2076) );
  OAI21X1 U1758 ( .A(n1950), .B(n2011), .C(n2076), .Y(n2591) );
  NAND2X1 U1759 ( .A(\mem<22><9> ), .B(n7), .Y(n2077) );
  OAI21X1 U1760 ( .A(n1950), .B(n2013), .C(n2077), .Y(n2590) );
  NAND2X1 U1761 ( .A(\mem<22><10> ), .B(n7), .Y(n2078) );
  OAI21X1 U1762 ( .A(n1950), .B(n2015), .C(n2078), .Y(n2589) );
  NAND2X1 U1763 ( .A(\mem<22><11> ), .B(n7), .Y(n2079) );
  OAI21X1 U1764 ( .A(n1950), .B(n2018), .C(n2079), .Y(n2588) );
  NAND2X1 U1765 ( .A(\mem<22><12> ), .B(n7), .Y(n2080) );
  OAI21X1 U1766 ( .A(n1950), .B(n2020), .C(n2080), .Y(n2587) );
  NAND2X1 U1767 ( .A(\mem<22><13> ), .B(n7), .Y(n2081) );
  OAI21X1 U1768 ( .A(n1950), .B(n2022), .C(n2081), .Y(n2586) );
  NAND2X1 U1769 ( .A(\mem<22><14> ), .B(n7), .Y(n2082) );
  OAI21X1 U1770 ( .A(n1950), .B(n2024), .C(n2082), .Y(n2585) );
  NAND2X1 U1771 ( .A(\mem<22><15> ), .B(n7), .Y(n2083) );
  OAI21X1 U1772 ( .A(n1950), .B(n1377), .C(n2083), .Y(n2584) );
  NAND2X1 U1773 ( .A(\mem<21><0> ), .B(n9), .Y(n2084) );
  OAI21X1 U1774 ( .A(n1951), .B(n1996), .C(n2084), .Y(n2583) );
  NAND2X1 U1775 ( .A(\mem<21><1> ), .B(n9), .Y(n2085) );
  OAI21X1 U1776 ( .A(n1951), .B(n1997), .C(n2085), .Y(n2582) );
  NAND2X1 U1777 ( .A(\mem<21><2> ), .B(n9), .Y(n2086) );
  OAI21X1 U1778 ( .A(n1951), .B(n1999), .C(n2086), .Y(n2581) );
  NAND2X1 U1779 ( .A(\mem<21><3> ), .B(n9), .Y(n2087) );
  OAI21X1 U1780 ( .A(n1951), .B(n2001), .C(n2087), .Y(n2580) );
  NAND2X1 U1781 ( .A(\mem<21><4> ), .B(n9), .Y(n2088) );
  OAI21X1 U1782 ( .A(n1951), .B(n2003), .C(n2088), .Y(n2579) );
  NAND2X1 U1783 ( .A(\mem<21><5> ), .B(n9), .Y(n2089) );
  OAI21X1 U1784 ( .A(n1951), .B(n2005), .C(n2089), .Y(n2578) );
  NAND2X1 U1785 ( .A(\mem<21><6> ), .B(n9), .Y(n2090) );
  OAI21X1 U1786 ( .A(n1951), .B(n2007), .C(n2090), .Y(n2577) );
  NAND2X1 U1787 ( .A(\mem<21><7> ), .B(n9), .Y(n2091) );
  OAI21X1 U1788 ( .A(n1951), .B(n2009), .C(n2091), .Y(n2576) );
  NAND2X1 U1789 ( .A(\mem<21><8> ), .B(n9), .Y(n2092) );
  OAI21X1 U1790 ( .A(n1952), .B(n2011), .C(n2092), .Y(n2575) );
  NAND2X1 U1791 ( .A(\mem<21><9> ), .B(n9), .Y(n2093) );
  OAI21X1 U1792 ( .A(n1952), .B(n2013), .C(n2093), .Y(n2574) );
  NAND2X1 U1793 ( .A(\mem<21><10> ), .B(n9), .Y(n2094) );
  OAI21X1 U1794 ( .A(n1952), .B(n2015), .C(n2094), .Y(n2573) );
  NAND2X1 U1795 ( .A(\mem<21><11> ), .B(n9), .Y(n2095) );
  OAI21X1 U1796 ( .A(n1952), .B(n2018), .C(n2095), .Y(n2572) );
  NAND2X1 U1797 ( .A(\mem<21><12> ), .B(n9), .Y(n2096) );
  OAI21X1 U1798 ( .A(n1952), .B(n2020), .C(n2096), .Y(n2571) );
  NAND2X1 U1799 ( .A(\mem<21><13> ), .B(n9), .Y(n2097) );
  OAI21X1 U1800 ( .A(n1952), .B(n2022), .C(n2097), .Y(n2570) );
  NAND2X1 U1801 ( .A(\mem<21><14> ), .B(n9), .Y(n2098) );
  OAI21X1 U1802 ( .A(n1952), .B(n2024), .C(n2098), .Y(n2569) );
  NAND2X1 U1803 ( .A(\mem<21><15> ), .B(n9), .Y(n2099) );
  OAI21X1 U1804 ( .A(n1952), .B(n1378), .C(n2099), .Y(n2568) );
  NAND2X1 U1805 ( .A(\mem<20><0> ), .B(n11), .Y(n2100) );
  OAI21X1 U1806 ( .A(n1953), .B(n1996), .C(n2100), .Y(n2567) );
  NAND2X1 U1807 ( .A(\mem<20><1> ), .B(n11), .Y(n2101) );
  OAI21X1 U1808 ( .A(n1953), .B(n1997), .C(n2101), .Y(n2566) );
  NAND2X1 U1809 ( .A(\mem<20><2> ), .B(n11), .Y(n2102) );
  OAI21X1 U1810 ( .A(n1953), .B(n1999), .C(n2102), .Y(n2565) );
  NAND2X1 U1811 ( .A(\mem<20><3> ), .B(n11), .Y(n2103) );
  OAI21X1 U1812 ( .A(n1953), .B(n2001), .C(n2103), .Y(n2564) );
  NAND2X1 U1813 ( .A(\mem<20><4> ), .B(n11), .Y(n2104) );
  OAI21X1 U1814 ( .A(n1953), .B(n2003), .C(n2104), .Y(n2563) );
  NAND2X1 U1815 ( .A(\mem<20><5> ), .B(n11), .Y(n2105) );
  OAI21X1 U1816 ( .A(n1953), .B(n2005), .C(n2105), .Y(n2562) );
  NAND2X1 U1817 ( .A(\mem<20><6> ), .B(n11), .Y(n2106) );
  OAI21X1 U1818 ( .A(n1953), .B(n2007), .C(n2106), .Y(n2561) );
  NAND2X1 U1819 ( .A(\mem<20><7> ), .B(n11), .Y(n2107) );
  OAI21X1 U1820 ( .A(n1953), .B(n2009), .C(n2107), .Y(n2560) );
  NAND2X1 U1821 ( .A(\mem<20><8> ), .B(n11), .Y(n2108) );
  OAI21X1 U1822 ( .A(n1954), .B(n2011), .C(n2108), .Y(n2559) );
  NAND2X1 U1823 ( .A(\mem<20><9> ), .B(n11), .Y(n2109) );
  OAI21X1 U1824 ( .A(n1954), .B(n2013), .C(n2109), .Y(n2558) );
  NAND2X1 U1825 ( .A(\mem<20><10> ), .B(n11), .Y(n2110) );
  OAI21X1 U1826 ( .A(n1954), .B(n2015), .C(n2110), .Y(n2557) );
  NAND2X1 U1827 ( .A(\mem<20><11> ), .B(n11), .Y(n2111) );
  OAI21X1 U1828 ( .A(n1954), .B(n2018), .C(n2111), .Y(n2556) );
  NAND2X1 U1829 ( .A(\mem<20><12> ), .B(n11), .Y(n2112) );
  OAI21X1 U1830 ( .A(n1954), .B(n2020), .C(n2112), .Y(n2555) );
  NAND2X1 U1831 ( .A(\mem<20><13> ), .B(n11), .Y(n2113) );
  OAI21X1 U1832 ( .A(n1954), .B(n2022), .C(n2113), .Y(n2554) );
  NAND2X1 U1833 ( .A(\mem<20><14> ), .B(n11), .Y(n2114) );
  OAI21X1 U1834 ( .A(n1954), .B(n2024), .C(n2114), .Y(n2553) );
  NAND2X1 U1835 ( .A(\mem<20><15> ), .B(n11), .Y(n2115) );
  OAI21X1 U1836 ( .A(n1954), .B(n1379), .C(n2115), .Y(n2552) );
  NAND2X1 U1837 ( .A(\mem<19><0> ), .B(n13), .Y(n2116) );
  OAI21X1 U1838 ( .A(n1955), .B(n1996), .C(n2116), .Y(n2551) );
  NAND2X1 U1839 ( .A(\mem<19><1> ), .B(n13), .Y(n2117) );
  OAI21X1 U1840 ( .A(n1955), .B(n1997), .C(n2117), .Y(n2550) );
  NAND2X1 U1841 ( .A(\mem<19><2> ), .B(n13), .Y(n2118) );
  OAI21X1 U1842 ( .A(n1955), .B(n1999), .C(n2118), .Y(n2549) );
  NAND2X1 U1843 ( .A(\mem<19><3> ), .B(n13), .Y(n2119) );
  OAI21X1 U1844 ( .A(n1955), .B(n2001), .C(n2119), .Y(n2548) );
  NAND2X1 U1845 ( .A(\mem<19><4> ), .B(n13), .Y(n2120) );
  OAI21X1 U1846 ( .A(n1955), .B(n2003), .C(n2120), .Y(n2547) );
  NAND2X1 U1847 ( .A(\mem<19><5> ), .B(n13), .Y(n2121) );
  OAI21X1 U1848 ( .A(n1955), .B(n2005), .C(n2121), .Y(n2546) );
  NAND2X1 U1849 ( .A(\mem<19><6> ), .B(n13), .Y(n2122) );
  OAI21X1 U1850 ( .A(n1955), .B(n2007), .C(n2122), .Y(n2545) );
  NAND2X1 U1851 ( .A(\mem<19><7> ), .B(n13), .Y(n2123) );
  OAI21X1 U1852 ( .A(n1955), .B(n2009), .C(n2123), .Y(n2544) );
  OAI21X1 U1853 ( .A(n1956), .B(n2011), .C(n389), .Y(n2543) );
  OAI21X1 U1854 ( .A(n1956), .B(n2013), .C(n391), .Y(n2542) );
  OAI21X1 U1855 ( .A(n1956), .B(n2015), .C(n393), .Y(n2541) );
  OAI21X1 U1856 ( .A(n1956), .B(n2018), .C(n395), .Y(n2540) );
  OAI21X1 U1857 ( .A(n1956), .B(n2020), .C(n397), .Y(n2539) );
  OAI21X1 U1858 ( .A(n1956), .B(n2022), .C(n399), .Y(n2538) );
  OAI21X1 U1859 ( .A(n1956), .B(n2024), .C(n401), .Y(n2537) );
  OAI21X1 U1860 ( .A(n1956), .B(n1380), .C(n61), .Y(n2536) );
  NAND2X1 U1861 ( .A(\mem<18><0> ), .B(n15), .Y(n2124) );
  OAI21X1 U1862 ( .A(n1957), .B(n1996), .C(n2124), .Y(n2535) );
  NAND2X1 U1863 ( .A(\mem<18><1> ), .B(n15), .Y(n2125) );
  OAI21X1 U1864 ( .A(n1957), .B(n1997), .C(n2125), .Y(n2534) );
  NAND2X1 U1865 ( .A(\mem<18><2> ), .B(n15), .Y(n2126) );
  OAI21X1 U1866 ( .A(n1957), .B(n1999), .C(n2126), .Y(n2533) );
  NAND2X1 U1867 ( .A(\mem<18><3> ), .B(n15), .Y(n2127) );
  OAI21X1 U1868 ( .A(n1957), .B(n2001), .C(n2127), .Y(n2532) );
  NAND2X1 U1869 ( .A(\mem<18><4> ), .B(n15), .Y(n2128) );
  OAI21X1 U1870 ( .A(n1957), .B(n2003), .C(n2128), .Y(n2531) );
  NAND2X1 U1871 ( .A(\mem<18><5> ), .B(n15), .Y(n2129) );
  OAI21X1 U1872 ( .A(n1957), .B(n2005), .C(n2129), .Y(n2530) );
  NAND2X1 U1873 ( .A(\mem<18><6> ), .B(n15), .Y(n2130) );
  OAI21X1 U1874 ( .A(n1957), .B(n2007), .C(n2130), .Y(n2529) );
  NAND2X1 U1875 ( .A(\mem<18><7> ), .B(n15), .Y(n2131) );
  OAI21X1 U1876 ( .A(n1957), .B(n2009), .C(n2131), .Y(n2528) );
  OAI21X1 U1877 ( .A(n1958), .B(n2011), .C(n403), .Y(n2527) );
  OAI21X1 U1878 ( .A(n1958), .B(n2013), .C(n405), .Y(n2526) );
  OAI21X1 U1879 ( .A(n1958), .B(n2015), .C(n407), .Y(n2525) );
  OAI21X1 U1880 ( .A(n1958), .B(n2018), .C(n409), .Y(n2524) );
  OAI21X1 U1881 ( .A(n1958), .B(n2020), .C(n411), .Y(n2523) );
  OAI21X1 U1882 ( .A(n1958), .B(n2022), .C(n413), .Y(n2522) );
  OAI21X1 U1883 ( .A(n1958), .B(n2024), .C(n415), .Y(n2521) );
  OAI21X1 U1884 ( .A(n1958), .B(n1364), .C(n417), .Y(n2520) );
  NAND2X1 U1885 ( .A(\mem<17><0> ), .B(n17), .Y(n2132) );
  OAI21X1 U1886 ( .A(n1959), .B(n1996), .C(n2132), .Y(n2519) );
  NAND2X1 U1887 ( .A(\mem<17><1> ), .B(n17), .Y(n2133) );
  OAI21X1 U1888 ( .A(n1959), .B(n1997), .C(n2133), .Y(n2518) );
  NAND2X1 U1889 ( .A(\mem<17><2> ), .B(n17), .Y(n2134) );
  OAI21X1 U1890 ( .A(n1959), .B(n1999), .C(n2134), .Y(n2517) );
  NAND2X1 U1891 ( .A(\mem<17><3> ), .B(n17), .Y(n2135) );
  OAI21X1 U1892 ( .A(n1959), .B(n2001), .C(n2135), .Y(n2516) );
  NAND2X1 U1893 ( .A(\mem<17><4> ), .B(n17), .Y(n2136) );
  OAI21X1 U1894 ( .A(n1959), .B(n2003), .C(n2136), .Y(n2515) );
  NAND2X1 U1895 ( .A(\mem<17><5> ), .B(n17), .Y(n2137) );
  OAI21X1 U1896 ( .A(n1959), .B(n2005), .C(n2137), .Y(n2514) );
  NAND2X1 U1897 ( .A(\mem<17><6> ), .B(n17), .Y(n2138) );
  OAI21X1 U1898 ( .A(n1959), .B(n2007), .C(n2138), .Y(n2513) );
  NAND2X1 U1899 ( .A(\mem<17><7> ), .B(n17), .Y(n2139) );
  OAI21X1 U1900 ( .A(n1959), .B(n2009), .C(n2139), .Y(n2512) );
  OAI21X1 U1901 ( .A(n1960), .B(n2011), .C(n419), .Y(n2511) );
  OAI21X1 U1902 ( .A(n1960), .B(n2013), .C(n421), .Y(n2510) );
  OAI21X1 U1903 ( .A(n1960), .B(n2015), .C(n423), .Y(n2509) );
  OAI21X1 U1904 ( .A(n1960), .B(n2018), .C(n425), .Y(n2508) );
  OAI21X1 U1905 ( .A(n1960), .B(n2020), .C(n427), .Y(n2507) );
  OAI21X1 U1906 ( .A(n1960), .B(n2022), .C(n429), .Y(n2506) );
  OAI21X1 U1907 ( .A(n1960), .B(n2024), .C(n431), .Y(n2505) );
  OAI21X1 U1908 ( .A(n1960), .B(n1364), .C(n433), .Y(n2504) );
  NAND2X1 U1909 ( .A(\mem<16><0> ), .B(n19), .Y(n2140) );
  OAI21X1 U1910 ( .A(n1961), .B(n1996), .C(n2140), .Y(n2503) );
  NAND2X1 U1911 ( .A(\mem<16><1> ), .B(n19), .Y(n2141) );
  OAI21X1 U1912 ( .A(n1961), .B(n1997), .C(n2141), .Y(n2502) );
  NAND2X1 U1913 ( .A(\mem<16><2> ), .B(n19), .Y(n2142) );
  OAI21X1 U1914 ( .A(n1961), .B(n1999), .C(n2142), .Y(n2501) );
  NAND2X1 U1915 ( .A(\mem<16><3> ), .B(n19), .Y(n2143) );
  OAI21X1 U1916 ( .A(n1961), .B(n2001), .C(n2143), .Y(n2500) );
  NAND2X1 U1917 ( .A(\mem<16><4> ), .B(n19), .Y(n2144) );
  OAI21X1 U1918 ( .A(n1961), .B(n2003), .C(n2144), .Y(n2499) );
  NAND2X1 U1919 ( .A(\mem<16><5> ), .B(n19), .Y(n2145) );
  OAI21X1 U1920 ( .A(n1961), .B(n2005), .C(n2145), .Y(n2498) );
  NAND2X1 U1921 ( .A(\mem<16><6> ), .B(n19), .Y(n2146) );
  OAI21X1 U1922 ( .A(n1961), .B(n2007), .C(n2146), .Y(n2497) );
  NAND2X1 U1923 ( .A(\mem<16><7> ), .B(n19), .Y(n2147) );
  OAI21X1 U1924 ( .A(n1961), .B(n2009), .C(n2147), .Y(n2496) );
  OAI21X1 U1925 ( .A(n1961), .B(n2011), .C(n435), .Y(n2495) );
  OAI21X1 U1926 ( .A(n1961), .B(n2013), .C(n437), .Y(n2494) );
  OAI21X1 U1927 ( .A(n1961), .B(n2015), .C(n439), .Y(n2493) );
  OAI21X1 U1928 ( .A(n1961), .B(n2018), .C(n441), .Y(n2492) );
  OAI21X1 U1929 ( .A(n1961), .B(n2020), .C(n443), .Y(n2491) );
  OAI21X1 U1930 ( .A(n1961), .B(n2022), .C(n445), .Y(n2490) );
  OAI21X1 U1931 ( .A(n1961), .B(n2024), .C(n447), .Y(n2489) );
  NAND2X1 U1932 ( .A(\mem<16><15> ), .B(n19), .Y(n2148) );
  OAI21X1 U1933 ( .A(n1961), .B(n1368), .C(n2148), .Y(n2488) );
  NAND3X1 U1934 ( .A(n2033), .B(n2744), .C(n2036), .Y(n2149) );
  NAND2X1 U1935 ( .A(\mem<15><0> ), .B(n21), .Y(n2150) );
  OAI21X1 U1936 ( .A(n1962), .B(n1996), .C(n2150), .Y(n2487) );
  NAND2X1 U1937 ( .A(\mem<15><1> ), .B(n21), .Y(n2151) );
  OAI21X1 U1938 ( .A(n1962), .B(n1997), .C(n2151), .Y(n2486) );
  NAND2X1 U1939 ( .A(\mem<15><2> ), .B(n21), .Y(n2152) );
  OAI21X1 U1940 ( .A(n1962), .B(n1999), .C(n2152), .Y(n2485) );
  NAND2X1 U1941 ( .A(\mem<15><3> ), .B(n21), .Y(n2153) );
  OAI21X1 U1942 ( .A(n1962), .B(n2001), .C(n2153), .Y(n2484) );
  NAND2X1 U1943 ( .A(\mem<15><4> ), .B(n21), .Y(n2154) );
  OAI21X1 U1944 ( .A(n1962), .B(n2003), .C(n2154), .Y(n2483) );
  NAND2X1 U1945 ( .A(\mem<15><5> ), .B(n21), .Y(n2155) );
  OAI21X1 U1946 ( .A(n1962), .B(n2005), .C(n2155), .Y(n2482) );
  NAND2X1 U1947 ( .A(\mem<15><6> ), .B(n21), .Y(n2156) );
  OAI21X1 U1948 ( .A(n1962), .B(n2007), .C(n2156), .Y(n2481) );
  NAND2X1 U1949 ( .A(\mem<15><7> ), .B(n21), .Y(n2157) );
  OAI21X1 U1950 ( .A(n1962), .B(n2009), .C(n2157), .Y(n2480) );
  OAI21X1 U1951 ( .A(n1963), .B(n2011), .C(n449), .Y(n2479) );
  OAI21X1 U1952 ( .A(n1963), .B(n2013), .C(n451), .Y(n2478) );
  OAI21X1 U1953 ( .A(n1963), .B(n2015), .C(n453), .Y(n2477) );
  OAI21X1 U1954 ( .A(n1963), .B(n2018), .C(n455), .Y(n2476) );
  OAI21X1 U1955 ( .A(n1963), .B(n2020), .C(n457), .Y(n2475) );
  OAI21X1 U1956 ( .A(n1963), .B(n2022), .C(n459), .Y(n2474) );
  OAI21X1 U1957 ( .A(n1963), .B(n2024), .C(n461), .Y(n2473) );
  OAI21X1 U1958 ( .A(n1963), .B(n1367), .C(n63), .Y(n2472) );
  NAND2X1 U1959 ( .A(\mem<14><0> ), .B(n23), .Y(n2158) );
  OAI21X1 U1960 ( .A(n1964), .B(n1996), .C(n2158), .Y(n2471) );
  NAND2X1 U1961 ( .A(\mem<14><1> ), .B(n23), .Y(n2159) );
  OAI21X1 U1962 ( .A(n1964), .B(n1997), .C(n2159), .Y(n2470) );
  NAND2X1 U1963 ( .A(\mem<14><2> ), .B(n23), .Y(n2160) );
  OAI21X1 U1964 ( .A(n1964), .B(n1999), .C(n2160), .Y(n2469) );
  NAND2X1 U1965 ( .A(\mem<14><3> ), .B(n23), .Y(n2161) );
  OAI21X1 U1966 ( .A(n1964), .B(n2001), .C(n2161), .Y(n2468) );
  NAND2X1 U1967 ( .A(\mem<14><4> ), .B(n23), .Y(n2162) );
  OAI21X1 U1968 ( .A(n1964), .B(n2003), .C(n2162), .Y(n2467) );
  NAND2X1 U1969 ( .A(\mem<14><5> ), .B(n23), .Y(n2163) );
  OAI21X1 U1970 ( .A(n1964), .B(n2005), .C(n2163), .Y(n2466) );
  NAND2X1 U1971 ( .A(\mem<14><6> ), .B(n23), .Y(n2164) );
  OAI21X1 U1972 ( .A(n1964), .B(n2007), .C(n2164), .Y(n2465) );
  NAND2X1 U1973 ( .A(\mem<14><7> ), .B(n23), .Y(n2165) );
  OAI21X1 U1974 ( .A(n1964), .B(n2009), .C(n2165), .Y(n2464) );
  OAI21X1 U1975 ( .A(n1965), .B(n2011), .C(n463), .Y(n2463) );
  OAI21X1 U1976 ( .A(n1965), .B(n2013), .C(n465), .Y(n2462) );
  OAI21X1 U1977 ( .A(n1965), .B(n2015), .C(n467), .Y(n2461) );
  OAI21X1 U1978 ( .A(n1965), .B(n2018), .C(n469), .Y(n2460) );
  OAI21X1 U1979 ( .A(n1965), .B(n2020), .C(n471), .Y(n2459) );
  OAI21X1 U1980 ( .A(n1965), .B(n2022), .C(n473), .Y(n2458) );
  OAI21X1 U1981 ( .A(n1965), .B(n2024), .C(n475), .Y(n2457) );
  OAI21X1 U1982 ( .A(n1965), .B(n1368), .C(n65), .Y(n2456) );
  NAND2X1 U1983 ( .A(\mem<13><0> ), .B(n25), .Y(n2166) );
  OAI21X1 U1984 ( .A(n1966), .B(n1996), .C(n2166), .Y(n2455) );
  NAND2X1 U1985 ( .A(\mem<13><1> ), .B(n25), .Y(n2167) );
  OAI21X1 U1986 ( .A(n1966), .B(n1997), .C(n2167), .Y(n2454) );
  NAND2X1 U1987 ( .A(\mem<13><2> ), .B(n25), .Y(n2168) );
  OAI21X1 U1988 ( .A(n1966), .B(n1999), .C(n2168), .Y(n2453) );
  NAND2X1 U1989 ( .A(\mem<13><3> ), .B(n25), .Y(n2169) );
  OAI21X1 U1990 ( .A(n1966), .B(n2001), .C(n2169), .Y(n2452) );
  NAND2X1 U1991 ( .A(\mem<13><4> ), .B(n25), .Y(n2170) );
  OAI21X1 U1992 ( .A(n1966), .B(n2003), .C(n2170), .Y(n2451) );
  NAND2X1 U1993 ( .A(\mem<13><5> ), .B(n25), .Y(n2171) );
  OAI21X1 U1994 ( .A(n1966), .B(n2005), .C(n2171), .Y(n2450) );
  NAND2X1 U1995 ( .A(\mem<13><6> ), .B(n25), .Y(n2172) );
  OAI21X1 U1996 ( .A(n1966), .B(n2007), .C(n2172), .Y(n2449) );
  NAND2X1 U1997 ( .A(\mem<13><7> ), .B(n25), .Y(n2173) );
  OAI21X1 U1998 ( .A(n1966), .B(n2009), .C(n2173), .Y(n2448) );
  OAI21X1 U1999 ( .A(n1967), .B(n2011), .C(n477), .Y(n2447) );
  OAI21X1 U2000 ( .A(n1967), .B(n2013), .C(n479), .Y(n2446) );
  OAI21X1 U2001 ( .A(n1967), .B(n2015), .C(n481), .Y(n2445) );
  OAI21X1 U2002 ( .A(n1967), .B(n2018), .C(n483), .Y(n2444) );
  OAI21X1 U2003 ( .A(n1967), .B(n2020), .C(n485), .Y(n2443) );
  OAI21X1 U2004 ( .A(n1967), .B(n2022), .C(n487), .Y(n2442) );
  OAI21X1 U2005 ( .A(n1967), .B(n2024), .C(n489), .Y(n2441) );
  OAI21X1 U2006 ( .A(n1967), .B(n1369), .C(n67), .Y(n2440) );
  NAND2X1 U2007 ( .A(\mem<12><0> ), .B(n27), .Y(n2174) );
  OAI21X1 U2008 ( .A(n1968), .B(n1996), .C(n2174), .Y(n2439) );
  NAND2X1 U2009 ( .A(\mem<12><1> ), .B(n27), .Y(n2175) );
  OAI21X1 U2010 ( .A(n1968), .B(n1997), .C(n2175), .Y(n2438) );
  NAND2X1 U2011 ( .A(\mem<12><2> ), .B(n27), .Y(n2176) );
  OAI21X1 U2012 ( .A(n1968), .B(n1999), .C(n2176), .Y(n2437) );
  NAND2X1 U2013 ( .A(\mem<12><3> ), .B(n27), .Y(n2177) );
  OAI21X1 U2014 ( .A(n1968), .B(n2001), .C(n2177), .Y(n2436) );
  NAND2X1 U2015 ( .A(\mem<12><4> ), .B(n27), .Y(n2178) );
  OAI21X1 U2016 ( .A(n1968), .B(n2003), .C(n2178), .Y(n2435) );
  NAND2X1 U2017 ( .A(\mem<12><5> ), .B(n27), .Y(n2179) );
  OAI21X1 U2018 ( .A(n1968), .B(n2005), .C(n2179), .Y(n2434) );
  NAND2X1 U2019 ( .A(\mem<12><6> ), .B(n27), .Y(n2180) );
  OAI21X1 U2020 ( .A(n1968), .B(n2007), .C(n2180), .Y(n2433) );
  NAND2X1 U2021 ( .A(\mem<12><7> ), .B(n27), .Y(n2181) );
  OAI21X1 U2022 ( .A(n1968), .B(n2009), .C(n2181), .Y(n2432) );
  OAI21X1 U2023 ( .A(n1969), .B(n2011), .C(n491), .Y(n2431) );
  OAI21X1 U2024 ( .A(n1969), .B(n2013), .C(n493), .Y(n2430) );
  OAI21X1 U2025 ( .A(n1969), .B(n2015), .C(n495), .Y(n2429) );
  OAI21X1 U2026 ( .A(n1969), .B(n2018), .C(n497), .Y(n2428) );
  OAI21X1 U2027 ( .A(n1969), .B(n2020), .C(n499), .Y(n2427) );
  OAI21X1 U2028 ( .A(n1969), .B(n2022), .C(n501), .Y(n2426) );
  OAI21X1 U2029 ( .A(n1969), .B(n2024), .C(n503), .Y(n2425) );
  OAI21X1 U2030 ( .A(n1969), .B(n1370), .C(n69), .Y(n2424) );
  NAND2X1 U2031 ( .A(\mem<11><0> ), .B(n29), .Y(n2182) );
  OAI21X1 U2032 ( .A(n1970), .B(n1996), .C(n2182), .Y(n2423) );
  NAND2X1 U2033 ( .A(\mem<11><1> ), .B(n29), .Y(n2183) );
  OAI21X1 U2034 ( .A(n1970), .B(n1997), .C(n2183), .Y(n2422) );
  NAND2X1 U2035 ( .A(\mem<11><2> ), .B(n29), .Y(n2184) );
  OAI21X1 U2036 ( .A(n1970), .B(n1999), .C(n2184), .Y(n2421) );
  NAND2X1 U2037 ( .A(\mem<11><3> ), .B(n29), .Y(n2185) );
  OAI21X1 U2038 ( .A(n1970), .B(n2001), .C(n2185), .Y(n2420) );
  NAND2X1 U2039 ( .A(\mem<11><4> ), .B(n29), .Y(n2186) );
  OAI21X1 U2040 ( .A(n1970), .B(n2003), .C(n2186), .Y(n2419) );
  NAND2X1 U2041 ( .A(\mem<11><5> ), .B(n29), .Y(n2187) );
  OAI21X1 U2042 ( .A(n1970), .B(n2005), .C(n2187), .Y(n2418) );
  NAND2X1 U2043 ( .A(\mem<11><6> ), .B(n29), .Y(n2188) );
  OAI21X1 U2044 ( .A(n1970), .B(n2007), .C(n2188), .Y(n2417) );
  NAND2X1 U2045 ( .A(\mem<11><7> ), .B(n29), .Y(n2189) );
  OAI21X1 U2046 ( .A(n1970), .B(n2009), .C(n2189), .Y(n2416) );
  OAI21X1 U2047 ( .A(n1971), .B(n2011), .C(n505), .Y(n2415) );
  OAI21X1 U2048 ( .A(n1971), .B(n2013), .C(n507), .Y(n2414) );
  OAI21X1 U2049 ( .A(n1971), .B(n2015), .C(n509), .Y(n2413) );
  OAI21X1 U2050 ( .A(n1971), .B(n2017), .C(n511), .Y(n2412) );
  OAI21X1 U2051 ( .A(n1971), .B(n2019), .C(n513), .Y(n2411) );
  OAI21X1 U2052 ( .A(n1971), .B(n2021), .C(n515), .Y(n2410) );
  OAI21X1 U2053 ( .A(n1971), .B(n2023), .C(n517), .Y(n2409) );
  OAI21X1 U2054 ( .A(n1971), .B(n1372), .C(n71), .Y(n2408) );
  NAND2X1 U2055 ( .A(\mem<10><0> ), .B(n31), .Y(n2190) );
  OAI21X1 U2056 ( .A(n1972), .B(n1996), .C(n2190), .Y(n2407) );
  NAND2X1 U2057 ( .A(\mem<10><1> ), .B(n31), .Y(n2191) );
  OAI21X1 U2058 ( .A(n1972), .B(n1997), .C(n2191), .Y(n2406) );
  NAND2X1 U2059 ( .A(\mem<10><2> ), .B(n31), .Y(n2192) );
  OAI21X1 U2060 ( .A(n1972), .B(n1999), .C(n2192), .Y(n2405) );
  NAND2X1 U2061 ( .A(\mem<10><3> ), .B(n31), .Y(n2193) );
  OAI21X1 U2062 ( .A(n1972), .B(n2001), .C(n2193), .Y(n2404) );
  NAND2X1 U2063 ( .A(\mem<10><4> ), .B(n31), .Y(n2194) );
  OAI21X1 U2064 ( .A(n1972), .B(n2003), .C(n2194), .Y(n2403) );
  NAND2X1 U2065 ( .A(\mem<10><5> ), .B(n31), .Y(n2195) );
  OAI21X1 U2066 ( .A(n1972), .B(n2005), .C(n2195), .Y(n2402) );
  NAND2X1 U2067 ( .A(\mem<10><6> ), .B(n31), .Y(n2196) );
  OAI21X1 U2068 ( .A(n1972), .B(n2007), .C(n2196), .Y(n2401) );
  NAND2X1 U2069 ( .A(\mem<10><7> ), .B(n31), .Y(n2197) );
  OAI21X1 U2070 ( .A(n1972), .B(n2009), .C(n2197), .Y(n2400) );
  OAI21X1 U2071 ( .A(n1973), .B(n2011), .C(n519), .Y(n2399) );
  OAI21X1 U2072 ( .A(n1973), .B(n2013), .C(n521), .Y(n2398) );
  OAI21X1 U2073 ( .A(n1973), .B(n2015), .C(n523), .Y(n2397) );
  OAI21X1 U2074 ( .A(n1973), .B(n2017), .C(n525), .Y(n2396) );
  OAI21X1 U2075 ( .A(n1973), .B(n2019), .C(n527), .Y(n2395) );
  OAI21X1 U2076 ( .A(n1973), .B(n2021), .C(n529), .Y(n2394) );
  OAI21X1 U2077 ( .A(n1973), .B(n2023), .C(n531), .Y(n2393) );
  OAI21X1 U2078 ( .A(n1973), .B(n1373), .C(n73), .Y(n2392) );
  NAND2X1 U2079 ( .A(\mem<9><0> ), .B(n33), .Y(n2198) );
  OAI21X1 U2080 ( .A(n1974), .B(n1996), .C(n2198), .Y(n2391) );
  NAND2X1 U2081 ( .A(\mem<9><1> ), .B(n33), .Y(n2199) );
  OAI21X1 U2082 ( .A(n1974), .B(n1997), .C(n2199), .Y(n2390) );
  NAND2X1 U2083 ( .A(\mem<9><2> ), .B(n33), .Y(n2200) );
  OAI21X1 U2084 ( .A(n1974), .B(n1999), .C(n2200), .Y(n2389) );
  NAND2X1 U2085 ( .A(\mem<9><3> ), .B(n33), .Y(n2201) );
  OAI21X1 U2086 ( .A(n1974), .B(n2001), .C(n2201), .Y(n2388) );
  NAND2X1 U2087 ( .A(\mem<9><4> ), .B(n33), .Y(n2202) );
  OAI21X1 U2088 ( .A(n1974), .B(n2003), .C(n2202), .Y(n2387) );
  NAND2X1 U2089 ( .A(\mem<9><5> ), .B(n33), .Y(n2203) );
  OAI21X1 U2090 ( .A(n1974), .B(n2005), .C(n2203), .Y(n2386) );
  NAND2X1 U2091 ( .A(\mem<9><6> ), .B(n33), .Y(n2204) );
  OAI21X1 U2092 ( .A(n1974), .B(n2007), .C(n2204), .Y(n2385) );
  NAND2X1 U2093 ( .A(\mem<9><7> ), .B(n33), .Y(n2205) );
  OAI21X1 U2094 ( .A(n1974), .B(n2009), .C(n2205), .Y(n2384) );
  OAI21X1 U2095 ( .A(n1975), .B(n2011), .C(n383), .Y(n2383) );
  OAI21X1 U2096 ( .A(n1975), .B(n2013), .C(n385), .Y(n2382) );
  OAI21X1 U2097 ( .A(n1975), .B(n2015), .C(n533), .Y(n2381) );
  OAI21X1 U2098 ( .A(n1975), .B(n2017), .C(n535), .Y(n2380) );
  OAI21X1 U2099 ( .A(n1975), .B(n2019), .C(n537), .Y(n2379) );
  OAI21X1 U2100 ( .A(n1975), .B(n2021), .C(n539), .Y(n2378) );
  OAI21X1 U2101 ( .A(n1975), .B(n2023), .C(n541), .Y(n2377) );
  OAI21X1 U2102 ( .A(n1975), .B(n1374), .C(n75), .Y(n2376) );
  NAND2X1 U2103 ( .A(\mem<8><0> ), .B(n35), .Y(n2207) );
  OAI21X1 U2104 ( .A(n1976), .B(n1996), .C(n2207), .Y(n2375) );
  OAI21X1 U2105 ( .A(n1976), .B(n1997), .C(n543), .Y(n2374) );
  OAI21X1 U2106 ( .A(n1976), .B(n1999), .C(n545), .Y(n2373) );
  OAI21X1 U2107 ( .A(n1976), .B(n2001), .C(n547), .Y(n2372) );
  OAI21X1 U2108 ( .A(n1976), .B(n2003), .C(n549), .Y(n2371) );
  OAI21X1 U2109 ( .A(n1976), .B(n2005), .C(n551), .Y(n2370) );
  OAI21X1 U2110 ( .A(n1976), .B(n2007), .C(n553), .Y(n2369) );
  OAI21X1 U2111 ( .A(n1976), .B(n2009), .C(n555), .Y(n2368) );
  OAI21X1 U2112 ( .A(n1976), .B(n2012), .C(n557), .Y(n2367) );
  OAI21X1 U2113 ( .A(n1976), .B(n2014), .C(n559), .Y(n2366) );
  OAI21X1 U2114 ( .A(n1976), .B(n2016), .C(n561), .Y(n2365) );
  OAI21X1 U2115 ( .A(n1976), .B(n2017), .C(n563), .Y(n2364) );
  OAI21X1 U2116 ( .A(n1976), .B(n2019), .C(n565), .Y(n2363) );
  OAI21X1 U2117 ( .A(n1976), .B(n2021), .C(n567), .Y(n2362) );
  OAI21X1 U2118 ( .A(n1976), .B(n2023), .C(n569), .Y(n2361) );
  NAND2X1 U2119 ( .A(\mem<8><15> ), .B(n35), .Y(n2208) );
  OAI21X1 U2120 ( .A(n1976), .B(n1369), .C(n2208), .Y(n2360) );
  NAND3X1 U2121 ( .A(n2034), .B(n2744), .C(n2036), .Y(n2209) );
  OAI21X1 U2122 ( .A(n1977), .B(n1996), .C(n77), .Y(n2359) );
  OAI21X1 U2123 ( .A(n1977), .B(n1997), .C(n571), .Y(n2358) );
  OAI21X1 U2124 ( .A(n1977), .B(n1999), .C(n573), .Y(n2357) );
  OAI21X1 U2125 ( .A(n1977), .B(n2001), .C(n575), .Y(n2356) );
  OAI21X1 U2126 ( .A(n1977), .B(n2003), .C(n577), .Y(n2355) );
  OAI21X1 U2127 ( .A(n1977), .B(n2005), .C(n579), .Y(n2354) );
  OAI21X1 U2128 ( .A(n1977), .B(n2007), .C(n581), .Y(n2353) );
  OAI21X1 U2129 ( .A(n1977), .B(n2009), .C(n583), .Y(n2352) );
  OAI21X1 U2130 ( .A(n1978), .B(n2011), .C(n585), .Y(n2351) );
  OAI21X1 U2131 ( .A(n1978), .B(n2013), .C(n587), .Y(n2350) );
  OAI21X1 U2132 ( .A(n1978), .B(n2015), .C(n589), .Y(n2349) );
  OAI21X1 U2133 ( .A(n1978), .B(n2017), .C(n591), .Y(n2348) );
  OAI21X1 U2134 ( .A(n1978), .B(n2019), .C(n593), .Y(n2347) );
  OAI21X1 U2135 ( .A(n1978), .B(n2021), .C(n595), .Y(n2346) );
  OAI21X1 U2136 ( .A(n1978), .B(n2023), .C(n597), .Y(n2345) );
  OAI21X1 U2137 ( .A(n1978), .B(n1378), .C(n79), .Y(n2344) );
  NAND2X1 U2138 ( .A(\mem<6><0> ), .B(n39), .Y(n2210) );
  OAI21X1 U2139 ( .A(n1979), .B(n1996), .C(n2210), .Y(n2343) );
  OAI21X1 U2140 ( .A(n1979), .B(n1997), .C(n599), .Y(n2342) );
  OAI21X1 U2141 ( .A(n1979), .B(n1999), .C(n601), .Y(n2341) );
  OAI21X1 U2142 ( .A(n1979), .B(n2001), .C(n603), .Y(n2340) );
  OAI21X1 U2143 ( .A(n1979), .B(n2003), .C(n605), .Y(n2339) );
  OAI21X1 U2144 ( .A(n1979), .B(n2005), .C(n607), .Y(n2338) );
  OAI21X1 U2145 ( .A(n1979), .B(n2007), .C(n609), .Y(n2337) );
  OAI21X1 U2146 ( .A(n1979), .B(n2009), .C(n611), .Y(n2336) );
  OAI21X1 U2147 ( .A(n1980), .B(n2011), .C(n613), .Y(n2335) );
  OAI21X1 U2148 ( .A(n1980), .B(n2013), .C(n615), .Y(n2334) );
  OAI21X1 U2149 ( .A(n1980), .B(n2015), .C(n617), .Y(n2333) );
  OAI21X1 U2150 ( .A(n1980), .B(n2017), .C(n619), .Y(n2332) );
  OAI21X1 U2151 ( .A(n1980), .B(n2019), .C(n621), .Y(n2331) );
  OAI21X1 U2152 ( .A(n1980), .B(n2021), .C(n623), .Y(n2330) );
  OAI21X1 U2153 ( .A(n1980), .B(n2023), .C(n625), .Y(n2329) );
  OAI21X1 U2154 ( .A(n1980), .B(n1376), .C(n81), .Y(n2328) );
  NAND2X1 U2155 ( .A(\mem<5><0> ), .B(n41), .Y(n2212) );
  OAI21X1 U2156 ( .A(n1981), .B(n1996), .C(n2212), .Y(n2327) );
  OAI21X1 U2157 ( .A(n1981), .B(n1998), .C(n627), .Y(n2326) );
  OAI21X1 U2158 ( .A(n1981), .B(n2000), .C(n629), .Y(n2325) );
  OAI21X1 U2159 ( .A(n1981), .B(n2002), .C(n631), .Y(n2324) );
  OAI21X1 U2160 ( .A(n1981), .B(n2004), .C(n633), .Y(n2323) );
  OAI21X1 U2161 ( .A(n1981), .B(n2006), .C(n635), .Y(n2322) );
  OAI21X1 U2162 ( .A(n1981), .B(n2008), .C(n637), .Y(n2321) );
  OAI21X1 U2163 ( .A(n1981), .B(n2010), .C(n639), .Y(n2320) );
  OAI21X1 U2164 ( .A(n1982), .B(n2011), .C(n641), .Y(n2319) );
  OAI21X1 U2165 ( .A(n1982), .B(n2013), .C(n643), .Y(n2318) );
  OAI21X1 U2166 ( .A(n1982), .B(n2015), .C(n645), .Y(n2317) );
  OAI21X1 U2167 ( .A(n1982), .B(n2017), .C(n647), .Y(n2316) );
  OAI21X1 U2168 ( .A(n1982), .B(n2019), .C(n649), .Y(n2315) );
  OAI21X1 U2169 ( .A(n1982), .B(n2021), .C(n1163), .Y(n2314) );
  OAI21X1 U2170 ( .A(n1982), .B(n2023), .C(n1165), .Y(n2313) );
  OAI21X1 U2171 ( .A(n1982), .B(n1377), .C(n83), .Y(n2312) );
  NAND2X1 U2172 ( .A(\mem<4><0> ), .B(n43), .Y(n2214) );
  OAI21X1 U2173 ( .A(n1983), .B(n1996), .C(n2214), .Y(n2311) );
  OAI21X1 U2174 ( .A(n1983), .B(n1997), .C(n1167), .Y(n2310) );
  OAI21X1 U2175 ( .A(n1983), .B(n1999), .C(n1169), .Y(n2309) );
  OAI21X1 U2176 ( .A(n1983), .B(n2001), .C(n1171), .Y(n2308) );
  OAI21X1 U2177 ( .A(n1983), .B(n2003), .C(n1173), .Y(n2307) );
  OAI21X1 U2178 ( .A(n1983), .B(n2005), .C(n1175), .Y(n2306) );
  OAI21X1 U2179 ( .A(n1983), .B(n2007), .C(n1177), .Y(n2305) );
  OAI21X1 U2180 ( .A(n1983), .B(n2009), .C(n1179), .Y(n2304) );
  OAI21X1 U2181 ( .A(n1984), .B(n2011), .C(n1181), .Y(n2303) );
  OAI21X1 U2182 ( .A(n1984), .B(n2013), .C(n1183), .Y(n2302) );
  OAI21X1 U2183 ( .A(n1984), .B(n2015), .C(n1185), .Y(n2301) );
  OAI21X1 U2184 ( .A(n1984), .B(n2017), .C(n1187), .Y(n2300) );
  OAI21X1 U2185 ( .A(n1984), .B(n2019), .C(n1189), .Y(n2299) );
  OAI21X1 U2186 ( .A(n1984), .B(n2021), .C(n1191), .Y(n2298) );
  OAI21X1 U2187 ( .A(n1984), .B(n2023), .C(n1193), .Y(n2297) );
  OAI21X1 U2188 ( .A(n1984), .B(n1379), .C(n85), .Y(n2296) );
  NAND2X1 U2189 ( .A(\mem<3><0> ), .B(n45), .Y(n2216) );
  OAI21X1 U2190 ( .A(n1985), .B(n1996), .C(n2216), .Y(n2295) );
  OAI21X1 U2191 ( .A(n1985), .B(n1997), .C(n1195), .Y(n2294) );
  OAI21X1 U2192 ( .A(n1985), .B(n1999), .C(n1197), .Y(n2293) );
  OAI21X1 U2193 ( .A(n1985), .B(n2001), .C(n1199), .Y(n2292) );
  OAI21X1 U2194 ( .A(n1985), .B(n2003), .C(n1201), .Y(n2291) );
  OAI21X1 U2195 ( .A(n1985), .B(n2005), .C(n1203), .Y(n2290) );
  OAI21X1 U2196 ( .A(n1985), .B(n2007), .C(n1205), .Y(n2289) );
  OAI21X1 U2197 ( .A(n1985), .B(n2009), .C(n1207), .Y(n2288) );
  OAI21X1 U2198 ( .A(n1986), .B(n2012), .C(n1209), .Y(n2287) );
  OAI21X1 U2199 ( .A(n1986), .B(n2014), .C(n1211), .Y(n2286) );
  OAI21X1 U2200 ( .A(n1986), .B(n2016), .C(n1213), .Y(n2285) );
  OAI21X1 U2201 ( .A(n1986), .B(n2017), .C(n1215), .Y(n2284) );
  OAI21X1 U2202 ( .A(n1986), .B(n2019), .C(n1217), .Y(n2283) );
  OAI21X1 U2203 ( .A(n1986), .B(n2021), .C(n1219), .Y(n2282) );
  OAI21X1 U2204 ( .A(n1986), .B(n2023), .C(n1221), .Y(n2281) );
  OAI21X1 U2205 ( .A(n1986), .B(n1365), .C(n87), .Y(n2280) );
  NAND2X1 U2206 ( .A(\mem<2><0> ), .B(n47), .Y(n2218) );
  OAI21X1 U2207 ( .A(n1987), .B(n1996), .C(n2218), .Y(n2279) );
  OAI21X1 U2208 ( .A(n1987), .B(n1998), .C(n1223), .Y(n2278) );
  OAI21X1 U2209 ( .A(n1987), .B(n2000), .C(n1225), .Y(n2277) );
  OAI21X1 U2210 ( .A(n1987), .B(n2002), .C(n1227), .Y(n2276) );
  OAI21X1 U2211 ( .A(n1987), .B(n2004), .C(n1229), .Y(n2275) );
  OAI21X1 U2212 ( .A(n1987), .B(n2006), .C(n1231), .Y(n2274) );
  OAI21X1 U2213 ( .A(n1987), .B(n2008), .C(n1233), .Y(n2273) );
  OAI21X1 U2214 ( .A(n1987), .B(n2010), .C(n1235), .Y(n2272) );
  OAI21X1 U2215 ( .A(n1988), .B(n2011), .C(n1237), .Y(n2271) );
  OAI21X1 U2216 ( .A(n1988), .B(n2013), .C(n1239), .Y(n2270) );
  OAI21X1 U2217 ( .A(n1988), .B(n2015), .C(n1241), .Y(n2269) );
  OAI21X1 U2218 ( .A(n1988), .B(n2017), .C(n1243), .Y(n2268) );
  OAI21X1 U2219 ( .A(n1988), .B(n2019), .C(n1245), .Y(n2267) );
  OAI21X1 U2220 ( .A(n1988), .B(n2021), .C(n1247), .Y(n2266) );
  OAI21X1 U2221 ( .A(n1988), .B(n2023), .C(n1249), .Y(n2265) );
  OAI21X1 U2222 ( .A(n1988), .B(n1366), .C(n89), .Y(n2264) );
  NAND2X1 U2223 ( .A(\mem<1><0> ), .B(n49), .Y(n2220) );
  OAI21X1 U2224 ( .A(n1989), .B(n1996), .C(n2220), .Y(n2263) );
  OAI21X1 U2225 ( .A(n1989), .B(n1997), .C(n1251), .Y(n2262) );
  OAI21X1 U2226 ( .A(n1989), .B(n1999), .C(n1253), .Y(n2261) );
  OAI21X1 U2227 ( .A(n1989), .B(n2001), .C(n1255), .Y(n2260) );
  OAI21X1 U2228 ( .A(n1989), .B(n2003), .C(n1257), .Y(n2259) );
  OAI21X1 U2229 ( .A(n1989), .B(n2005), .C(n1259), .Y(n2258) );
  OAI21X1 U2230 ( .A(n1989), .B(n2007), .C(n1261), .Y(n2257) );
  OAI21X1 U2231 ( .A(n1989), .B(n2009), .C(n1263), .Y(n2256) );
  OAI21X1 U2232 ( .A(n1990), .B(n2011), .C(n1265), .Y(n2255) );
  OAI21X1 U2233 ( .A(n1990), .B(n2013), .C(n1267), .Y(n2254) );
  OAI21X1 U2234 ( .A(n1990), .B(n2015), .C(n1269), .Y(n2253) );
  OAI21X1 U2235 ( .A(n1990), .B(n2017), .C(n1271), .Y(n2252) );
  OAI21X1 U2236 ( .A(n1990), .B(n2019), .C(n1273), .Y(n2251) );
  OAI21X1 U2237 ( .A(n1990), .B(n2021), .C(n1275), .Y(n2250) );
  OAI21X1 U2238 ( .A(n1990), .B(n2023), .C(n1277), .Y(n2249) );
  OAI21X1 U2239 ( .A(n1990), .B(n1367), .C(n91), .Y(n2248) );
  NAND2X1 U2240 ( .A(\mem<0><0> ), .B(n51), .Y(n2223) );
  OAI21X1 U2241 ( .A(n1991), .B(n1996), .C(n2223), .Y(n2247) );
  NAND2X1 U2242 ( .A(\mem<0><1> ), .B(n51), .Y(n2224) );
  OAI21X1 U2243 ( .A(n1991), .B(n1997), .C(n2224), .Y(n2246) );
  NAND2X1 U2244 ( .A(\mem<0><2> ), .B(n51), .Y(n2225) );
  OAI21X1 U2245 ( .A(n1991), .B(n1999), .C(n2225), .Y(n2245) );
  NAND2X1 U2246 ( .A(\mem<0><3> ), .B(n51), .Y(n2226) );
  OAI21X1 U2247 ( .A(n1991), .B(n2001), .C(n2226), .Y(n2244) );
  NAND2X1 U2248 ( .A(\mem<0><4> ), .B(n51), .Y(n2227) );
  OAI21X1 U2249 ( .A(n1991), .B(n2003), .C(n2227), .Y(n2243) );
  NAND2X1 U2250 ( .A(\mem<0><5> ), .B(n51), .Y(n2228) );
  OAI21X1 U2251 ( .A(n1991), .B(n2005), .C(n2228), .Y(n2242) );
  NAND2X1 U2252 ( .A(\mem<0><6> ), .B(n51), .Y(n2229) );
  OAI21X1 U2253 ( .A(n1991), .B(n2007), .C(n2229), .Y(n2241) );
  NAND2X1 U2254 ( .A(\mem<0><7> ), .B(n51), .Y(n2230) );
  OAI21X1 U2255 ( .A(n1991), .B(n2009), .C(n2230), .Y(n2240) );
  OAI21X1 U2256 ( .A(n1991), .B(n2011), .C(n1279), .Y(n2239) );
  OAI21X1 U2257 ( .A(n1991), .B(n2013), .C(n1281), .Y(n2238) );
  OAI21X1 U2258 ( .A(n1991), .B(n2015), .C(n1283), .Y(n2237) );
  OAI21X1 U2259 ( .A(n1991), .B(n2017), .C(n1285), .Y(n2236) );
  OAI21X1 U2260 ( .A(n1991), .B(n2019), .C(n1287), .Y(n2235) );
  OAI21X1 U2261 ( .A(n1991), .B(n2021), .C(n1289), .Y(n2234) );
  OAI21X1 U2262 ( .A(n1991), .B(n2023), .C(n1291), .Y(n2233) );
  NAND2X1 U2263 ( .A(\mem<0><15> ), .B(n51), .Y(n2231) );
  OAI21X1 U2264 ( .A(n1991), .B(n1370), .C(n2231), .Y(n2232) );
endmodule


module memc_Size16_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2261), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2262), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2263), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2264), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2265), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2266), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2267), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2268), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2269), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2270), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2271), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2272), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2273), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2274), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2275), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2276), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2277), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2278), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2279), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2280), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2281), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2282), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2283), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2284), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2285), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2286), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2287), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2288), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2289), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2290), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2291), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2292), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2293), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2294), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2295), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2296), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2297), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2298), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2299), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2300), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2301), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2302), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2303), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2304), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2305), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2306), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2307), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2308), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2309), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2310), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2311), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2312), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2313), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2314), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2315), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2316), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2317), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2318), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2319), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2320), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2321), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2322), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2323), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2324), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2325), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2326), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2327), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2328), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2329), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2330), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2331), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2332), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2333), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2334), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2335), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2336), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2337), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2338), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2339), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2340), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2341), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2342), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2343), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2344), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2345), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2346), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2347), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2348), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2349), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2350), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2351), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2352), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2353), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2354), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2355), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2356), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2357), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2358), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2359), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2360), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2361), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2362), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2363), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2364), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2365), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2366), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2367), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2368), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2369), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2370), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2371), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2372), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2373), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2374), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2375), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2376), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2377), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2378), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2379), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2380), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2381), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2382), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2383), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2384), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2385), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2386), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2387), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2388), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2389), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2390), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2391), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2392), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2393), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2394), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2395), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2396), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2397), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2398), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2399), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2400), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2401), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2402), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2403), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2404), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2405), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2406), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2407), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2408), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2409), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2410), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2411), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2412), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2413), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2414), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2415), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2416), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2417), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2418), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2419), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2420), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2421), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2422), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2423), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2424), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2425), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2426), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2427), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2428), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2429), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2430), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2431), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2432), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2433), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2434), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2435), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2436), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2437), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2438), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2439), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2440), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2441), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2442), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2443), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2444), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2445), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2446), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2447), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2448), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2449), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2450), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2451), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2452), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2453), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2454), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2455), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2456), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2457), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2458), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2459), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2460), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2461), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2462), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2463), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2464), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2465), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2466), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2467), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2468), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2469), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2470), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2471), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2472), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2473), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2474), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2475), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2476), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2477), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2478), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2479), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2480), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2481), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2482), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2483), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2484), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2485), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2486), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2487), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2488), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2489), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2490), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2491), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2492), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2493), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2494), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2495), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2496), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2497), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2498), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2499), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2500), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2501), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2502), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2503), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2504), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2505), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2506), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2507), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2508), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2509), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2510), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2511), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2512), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2513), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2514), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2515), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2516), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2517), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2518), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2519), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2520), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2521), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2522), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2523), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2524), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2525), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2526), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2527), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2528), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2529), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2530), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2531), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2532), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2533), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2534), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2535), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2536), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2537), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2538), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2539), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2540), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2541), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2542), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2543), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2544), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2545), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2546), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2547), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2548), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2549), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2550), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2551), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2552), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2553), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2554), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2555), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2556), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2557), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2558), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2559), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2560), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2561), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2562), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2563), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2564), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2565), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2566), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2567), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2568), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2569), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2570), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2571), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2572), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2573), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2574), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2575), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2576), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2577), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2578), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2579), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2580), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2581), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2582), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2583), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2584), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2585), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2586), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2587), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2588), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2589), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2590), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2591), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2592), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2593), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2594), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2595), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2596), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2597), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2598), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2599), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2600), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2601), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2602), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2603), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2604), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2605), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2606), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2607), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2608), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2609), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2610), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2611), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2612), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2613), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2614), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2615), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2616), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2617), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2618), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2619), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2620), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2621), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2622), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2623), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2624), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2625), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2626), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2627), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2628), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2629), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2630), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2631), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2632), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2633), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2634), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2635), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2636), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2637), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2638), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2639), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2640), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2641), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2642), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2643), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2644), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2645), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2646), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2647), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2648), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2649), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2650), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2651), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2652), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2653), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2654), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2655), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2656), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2657), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2658), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2659), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2660), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2661), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2662), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2663), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2664), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2665), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2666), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2667), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2668), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2669), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2670), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2671), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2672), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2673), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2674), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2675), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2676), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2677), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2678), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2679), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2680), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2681), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2682), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2683), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2684), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2685), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2686), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2687), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2688), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2689), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2690), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2691), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2692), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2693), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2694), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2695), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2696), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2697), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2698), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2699), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2700), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2701), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2702), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2703), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2704), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2705), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2706), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2707), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2708), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2709), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2710), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2711), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2712), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2713), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2714), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2715), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2716), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2717), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2718), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2719), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2720), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2721), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2722), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2723), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2724), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2725), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2726), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2727), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2728), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2729), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2730), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2731), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2732), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2733), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2734), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2735), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2736), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2737), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2738), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2739), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2740), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2741), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2742), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2743), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2744), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2745), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2746), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2747), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2748), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2749), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2750), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2751), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2752), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2753), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2754), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2755), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2756), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2757), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2758), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2759), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2760), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2761), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2762), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2763), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2764), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2765), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2766), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2767), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2768), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2769), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2770), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2771), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2772), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2773) );
  INVX4 U2 ( .A(n270), .Y(n271) );
  INVX4 U3 ( .A(n268), .Y(n269) );
  INVX4 U4 ( .A(n266), .Y(n267) );
  INVX4 U5 ( .A(n264), .Y(n265) );
  INVX4 U6 ( .A(n262), .Y(n263) );
  INVX4 U7 ( .A(n260), .Y(n261) );
  INVX4 U8 ( .A(n258), .Y(n259) );
  INVX4 U9 ( .A(n256), .Y(n257) );
  INVX4 U10 ( .A(n205), .Y(n206) );
  INVX4 U11 ( .A(n203), .Y(n204) );
  INVX4 U12 ( .A(n201), .Y(n202) );
  INVX4 U13 ( .A(n199), .Y(n200) );
  INVX4 U14 ( .A(n197), .Y(n198) );
  INVX4 U15 ( .A(n195), .Y(n196) );
  INVX4 U16 ( .A(n193), .Y(n194) );
  INVX4 U17 ( .A(n191), .Y(n192) );
  INVX4 U18 ( .A(n189), .Y(n190) );
  INVX4 U19 ( .A(n187), .Y(n188) );
  INVX4 U20 ( .A(n185), .Y(n186) );
  INVX1 U21 ( .A(n2115), .Y(n1972) );
  INVX1 U22 ( .A(n2115), .Y(n1971) );
  INVX1 U23 ( .A(n2115), .Y(n1970) );
  INVX1 U24 ( .A(n1954), .Y(N31) );
  INVX1 U25 ( .A(n1955), .Y(N30) );
  INVX1 U26 ( .A(n1956), .Y(N29) );
  INVX1 U27 ( .A(n1958), .Y(N27) );
  INVX1 U28 ( .A(n1960), .Y(N25) );
  INVX1 U29 ( .A(n1966), .Y(N19) );
  INVX1 U30 ( .A(n1967), .Y(N18) );
  INVX1 U31 ( .A(n1968), .Y(N17) );
  INVX1 U32 ( .A(n1953), .Y(N32) );
  INVX1 U33 ( .A(n1957), .Y(N28) );
  INVX1 U34 ( .A(n1959), .Y(N26) );
  INVX1 U35 ( .A(n1961), .Y(N24) );
  INVX1 U36 ( .A(n1962), .Y(N23) );
  INVX1 U37 ( .A(n1963), .Y(N22) );
  INVX1 U38 ( .A(n1964), .Y(N21) );
  INVX1 U39 ( .A(n1965), .Y(N20) );
  BUFX2 U40 ( .A(n1389), .Y(n2013) );
  BUFX2 U41 ( .A(n1391), .Y(n2015) );
  BUFX2 U42 ( .A(n1393), .Y(n2017) );
  BUFX2 U43 ( .A(n1395), .Y(n2019) );
  BUFX2 U44 ( .A(n1397), .Y(n2021) );
  BUFX2 U45 ( .A(n1399), .Y(n2023) );
  BUFX2 U46 ( .A(n1401), .Y(n2025) );
  BUFX2 U47 ( .A(n1403), .Y(n2028) );
  BUFX2 U48 ( .A(n1405), .Y(n2030) );
  BUFX2 U49 ( .A(n1407), .Y(n2032) );
  BUFX2 U50 ( .A(n1409), .Y(n2034) );
  BUFX2 U51 ( .A(n1411), .Y(n2036) );
  BUFX2 U52 ( .A(n1413), .Y(n2039) );
  BUFX2 U53 ( .A(n1415), .Y(n2041) );
  BUFX2 U54 ( .A(n1417), .Y(n2044) );
  BUFX2 U55 ( .A(n1419), .Y(n2046) );
  BUFX2 U56 ( .A(n1421), .Y(n2048) );
  BUFX2 U57 ( .A(n1423), .Y(n2050) );
  BUFX2 U58 ( .A(n1425), .Y(n2052) );
  BUFX2 U59 ( .A(n1427), .Y(n2054) );
  BUFX2 U60 ( .A(n1429), .Y(n2056) );
  BUFX2 U61 ( .A(n1431), .Y(n2059) );
  BUFX2 U62 ( .A(n1433), .Y(n2061) );
  BUFX2 U63 ( .A(n1435), .Y(n2063) );
  BUFX2 U64 ( .A(n1437), .Y(n2065) );
  BUFX2 U65 ( .A(n1439), .Y(n2067) );
  BUFX2 U66 ( .A(n1441), .Y(n2069) );
  BUFX2 U67 ( .A(n1443), .Y(n2071) );
  INVX8 U68 ( .A(n2010), .Y(n2012) );
  INVX2 U69 ( .A(n2113), .Y(n1973) );
  INVX1 U70 ( .A(n2110), .Y(n1975) );
  INVX2 U71 ( .A(n1975), .Y(n1979) );
  INVX2 U72 ( .A(n1975), .Y(n1981) );
  INVX2 U73 ( .A(n1975), .Y(n1980) );
  INVX4 U74 ( .A(n2108), .Y(n2010) );
  INVX2 U75 ( .A(n2113), .Y(n1974) );
  INVX1 U76 ( .A(n2110), .Y(n1976) );
  INVX2 U77 ( .A(n1976), .Y(n1978) );
  INVX2 U78 ( .A(n1976), .Y(n1977) );
  INVX2 U79 ( .A(n1976), .Y(n1983) );
  BUFX2 U80 ( .A(n1389), .Y(n2014) );
  INVX1 U81 ( .A(n2110), .Y(n1984) );
  BUFX2 U82 ( .A(n1403), .Y(n2029) );
  BUFX2 U83 ( .A(n1417), .Y(n2045) );
  BUFX2 U84 ( .A(n1431), .Y(n2060) );
  BUFX2 U85 ( .A(n1437), .Y(n2066) );
  INVX1 U86 ( .A(n2010), .Y(n2011) );
  INVX1 U87 ( .A(n1387), .Y(n2073) );
  INVX1 U88 ( .A(n1386), .Y(n2058) );
  INVX1 U89 ( .A(write), .Y(n1469) );
  BUFX2 U90 ( .A(n1391), .Y(n2016) );
  BUFX2 U91 ( .A(n1411), .Y(n2037) );
  BUFX2 U92 ( .A(n1413), .Y(n2040) );
  BUFX2 U93 ( .A(n1415), .Y(n2042) );
  BUFX2 U94 ( .A(n1405), .Y(n2031) );
  BUFX2 U95 ( .A(n1407), .Y(n2033) );
  BUFX2 U96 ( .A(n1409), .Y(n2035) );
  BUFX2 U97 ( .A(n1393), .Y(n2018) );
  BUFX2 U98 ( .A(n1395), .Y(n2020) );
  BUFX2 U99 ( .A(n1397), .Y(n2022) );
  BUFX2 U100 ( .A(n1399), .Y(n2024) );
  BUFX2 U101 ( .A(n1401), .Y(n2026) );
  BUFX2 U102 ( .A(n1421), .Y(n2049) );
  BUFX2 U103 ( .A(n1423), .Y(n2051) );
  BUFX2 U104 ( .A(n1425), .Y(n2053) );
  BUFX2 U105 ( .A(n1427), .Y(n2055) );
  BUFX2 U106 ( .A(n1429), .Y(n2057) );
  BUFX2 U107 ( .A(n1433), .Y(n2062) );
  BUFX2 U108 ( .A(n1435), .Y(n2064) );
  BUFX2 U109 ( .A(n1439), .Y(n2068) );
  BUFX2 U110 ( .A(n1441), .Y(n2070) );
  BUFX2 U111 ( .A(n1443), .Y(n2072) );
  INVX1 U112 ( .A(n2115), .Y(n2114) );
  INVX1 U113 ( .A(N13), .Y(n2115) );
  INVX1 U114 ( .A(N14), .Y(n2116) );
  INVX1 U115 ( .A(n1384), .Y(n2027) );
  BUFX2 U116 ( .A(n1419), .Y(n2047) );
  INVX1 U117 ( .A(n1385), .Y(n2043) );
  INVX1 U118 ( .A(n2116), .Y(n1969) );
  AND2X2 U119 ( .A(\mem<31><0> ), .B(n209), .Y(n1) );
  INVX1 U120 ( .A(n1), .Y(n2) );
  AND2X2 U121 ( .A(\mem<31><1> ), .B(n209), .Y(n3) );
  INVX1 U122 ( .A(n3), .Y(n4) );
  AND2X2 U123 ( .A(\mem<31><2> ), .B(n209), .Y(n5) );
  INVX1 U124 ( .A(n5), .Y(n6) );
  AND2X2 U125 ( .A(\mem<31><3> ), .B(n209), .Y(n7) );
  INVX1 U126 ( .A(n7), .Y(n8) );
  AND2X2 U127 ( .A(\mem<31><4> ), .B(n209), .Y(n9) );
  INVX1 U128 ( .A(n9), .Y(n10) );
  AND2X2 U129 ( .A(\mem<31><5> ), .B(n209), .Y(n11) );
  INVX1 U130 ( .A(n11), .Y(n12) );
  AND2X2 U131 ( .A(\mem<31><6> ), .B(n209), .Y(n13) );
  INVX1 U132 ( .A(n13), .Y(n14) );
  AND2X2 U133 ( .A(\mem<30><8> ), .B(n211), .Y(n15) );
  INVX1 U134 ( .A(n15), .Y(n16) );
  AND2X2 U135 ( .A(\mem<30><9> ), .B(n211), .Y(n17) );
  INVX1 U136 ( .A(n17), .Y(n18) );
  AND2X2 U137 ( .A(\mem<30><10> ), .B(n211), .Y(n19) );
  INVX1 U138 ( .A(n19), .Y(n20) );
  AND2X2 U139 ( .A(\mem<30><11> ), .B(n211), .Y(n21) );
  INVX1 U140 ( .A(n21), .Y(n22) );
  AND2X2 U141 ( .A(\mem<30><12> ), .B(n211), .Y(n23) );
  INVX1 U142 ( .A(n23), .Y(n24) );
  AND2X2 U143 ( .A(\mem<30><13> ), .B(n211), .Y(n25) );
  INVX1 U144 ( .A(n25), .Y(n26) );
  AND2X2 U145 ( .A(\mem<30><14> ), .B(n211), .Y(n27) );
  INVX1 U146 ( .A(n27), .Y(n28) );
  AND2X2 U147 ( .A(\mem<29><8> ), .B(n213), .Y(n29) );
  INVX1 U148 ( .A(n29), .Y(n30) );
  AND2X2 U149 ( .A(\mem<29><9> ), .B(n213), .Y(n31) );
  INVX1 U150 ( .A(n31), .Y(n32) );
  AND2X2 U151 ( .A(\mem<29><10> ), .B(n213), .Y(n33) );
  INVX1 U152 ( .A(n33), .Y(n34) );
  AND2X2 U153 ( .A(\mem<29><11> ), .B(n213), .Y(n35) );
  INVX1 U154 ( .A(n35), .Y(n36) );
  AND2X2 U155 ( .A(\mem<29><12> ), .B(n213), .Y(n37) );
  INVX1 U156 ( .A(n37), .Y(n38) );
  AND2X2 U157 ( .A(\mem<29><13> ), .B(n213), .Y(n39) );
  INVX1 U158 ( .A(n39), .Y(n40) );
  AND2X2 U159 ( .A(\mem<29><14> ), .B(n213), .Y(n41) );
  INVX1 U160 ( .A(n41), .Y(n42) );
  AND2X2 U161 ( .A(\mem<28><8> ), .B(n216), .Y(n43) );
  INVX1 U162 ( .A(n43), .Y(n44) );
  AND2X2 U163 ( .A(\mem<28><9> ), .B(n216), .Y(n45) );
  INVX1 U164 ( .A(n45), .Y(n46) );
  AND2X2 U165 ( .A(\mem<28><10> ), .B(n216), .Y(n47) );
  INVX1 U166 ( .A(n47), .Y(n48) );
  AND2X2 U167 ( .A(\mem<28><11> ), .B(n216), .Y(n49) );
  INVX1 U168 ( .A(n49), .Y(n50) );
  AND2X2 U169 ( .A(\mem<28><12> ), .B(n216), .Y(n51) );
  INVX1 U170 ( .A(n51), .Y(n52) );
  AND2X2 U171 ( .A(\mem<28><13> ), .B(n216), .Y(n53) );
  INVX1 U172 ( .A(n53), .Y(n54) );
  AND2X2 U173 ( .A(\mem<28><14> ), .B(n216), .Y(n55) );
  INVX1 U174 ( .A(n55), .Y(n56) );
  AND2X2 U175 ( .A(\mem<27><8> ), .B(n218), .Y(n57) );
  INVX1 U176 ( .A(n57), .Y(n58) );
  AND2X2 U177 ( .A(\mem<27><9> ), .B(n218), .Y(n59) );
  INVX1 U178 ( .A(n59), .Y(n60) );
  AND2X2 U179 ( .A(\mem<27><10> ), .B(n218), .Y(n61) );
  INVX1 U180 ( .A(n61), .Y(n62) );
  AND2X2 U181 ( .A(\mem<27><11> ), .B(n218), .Y(n63) );
  INVX1 U182 ( .A(n63), .Y(n64) );
  AND2X2 U183 ( .A(\mem<27><12> ), .B(n218), .Y(n65) );
  INVX1 U184 ( .A(n65), .Y(n66) );
  AND2X2 U185 ( .A(\mem<27><13> ), .B(n218), .Y(n67) );
  INVX1 U186 ( .A(n67), .Y(n68) );
  AND2X2 U187 ( .A(\mem<27><14> ), .B(n218), .Y(n69) );
  INVX1 U188 ( .A(n69), .Y(n70) );
  AND2X2 U189 ( .A(\mem<26><8> ), .B(n220), .Y(n71) );
  INVX1 U190 ( .A(n71), .Y(n72) );
  AND2X2 U191 ( .A(\mem<26><9> ), .B(n220), .Y(n73) );
  INVX1 U192 ( .A(n73), .Y(n74) );
  AND2X2 U193 ( .A(\mem<26><10> ), .B(n220), .Y(n75) );
  INVX1 U194 ( .A(n75), .Y(n76) );
  AND2X2 U195 ( .A(\mem<26><11> ), .B(n220), .Y(n77) );
  INVX1 U196 ( .A(n77), .Y(n78) );
  AND2X2 U197 ( .A(\mem<26><12> ), .B(n220), .Y(n79) );
  INVX1 U198 ( .A(n79), .Y(n80) );
  AND2X2 U199 ( .A(\mem<26><13> ), .B(n220), .Y(n81) );
  INVX1 U200 ( .A(n81), .Y(n82) );
  AND2X2 U201 ( .A(\mem<26><14> ), .B(n220), .Y(n83) );
  INVX1 U202 ( .A(n83), .Y(n84) );
  AND2X2 U203 ( .A(\mem<25><8> ), .B(n222), .Y(n85) );
  INVX1 U204 ( .A(n85), .Y(n86) );
  AND2X2 U205 ( .A(\mem<25><9> ), .B(n222), .Y(n87) );
  INVX1 U206 ( .A(n87), .Y(n88) );
  AND2X2 U207 ( .A(\mem<25><10> ), .B(n222), .Y(n89) );
  INVX1 U208 ( .A(n89), .Y(n90) );
  AND2X2 U209 ( .A(\mem<25><11> ), .B(n222), .Y(n91) );
  INVX1 U210 ( .A(n91), .Y(n92) );
  AND2X2 U211 ( .A(\mem<25><12> ), .B(n222), .Y(n93) );
  INVX1 U212 ( .A(n93), .Y(n94) );
  AND2X2 U213 ( .A(\mem<25><13> ), .B(n222), .Y(n95) );
  INVX1 U214 ( .A(n95), .Y(n96) );
  AND2X2 U215 ( .A(\mem<25><14> ), .B(n222), .Y(n97) );
  INVX1 U216 ( .A(n97), .Y(n98) );
  AND2X2 U217 ( .A(\mem<24><8> ), .B(n224), .Y(n99) );
  INVX1 U218 ( .A(n99), .Y(n100) );
  AND2X2 U219 ( .A(\mem<24><9> ), .B(n224), .Y(n101) );
  INVX1 U220 ( .A(n101), .Y(n102) );
  AND2X2 U221 ( .A(\mem<24><10> ), .B(n224), .Y(n103) );
  INVX1 U222 ( .A(n103), .Y(n104) );
  AND2X2 U223 ( .A(\mem<24><11> ), .B(n224), .Y(n105) );
  INVX1 U224 ( .A(n105), .Y(n106) );
  AND2X2 U225 ( .A(\mem<24><12> ), .B(n224), .Y(n107) );
  INVX1 U226 ( .A(n107), .Y(n108) );
  AND2X2 U227 ( .A(\mem<24><13> ), .B(n224), .Y(n109) );
  INVX1 U228 ( .A(n109), .Y(n110) );
  AND2X2 U229 ( .A(\mem<24><15> ), .B(n224), .Y(n111) );
  INVX1 U230 ( .A(n111), .Y(n112) );
  AND2X2 U231 ( .A(\mem<23><8> ), .B(n226), .Y(n113) );
  INVX1 U232 ( .A(n113), .Y(n114) );
  AND2X2 U233 ( .A(\mem<23><9> ), .B(n226), .Y(n115) );
  INVX1 U234 ( .A(n115), .Y(n116) );
  AND2X2 U235 ( .A(\mem<23><10> ), .B(n226), .Y(n117) );
  INVX1 U236 ( .A(n117), .Y(n118) );
  AND2X2 U237 ( .A(\mem<23><11> ), .B(n226), .Y(n119) );
  INVX1 U238 ( .A(n119), .Y(n120) );
  AND2X2 U239 ( .A(\mem<23><12> ), .B(n226), .Y(n121) );
  INVX1 U240 ( .A(n121), .Y(n122) );
  AND2X2 U241 ( .A(\mem<23><13> ), .B(n226), .Y(n123) );
  INVX1 U242 ( .A(n123), .Y(n124) );
  AND2X2 U243 ( .A(\mem<23><14> ), .B(n226), .Y(n125) );
  INVX1 U244 ( .A(n125), .Y(n126) );
  AND2X2 U245 ( .A(\mem<22><8> ), .B(n228), .Y(n127) );
  INVX1 U246 ( .A(n127), .Y(n128) );
  AND2X2 U247 ( .A(\mem<22><9> ), .B(n228), .Y(n129) );
  INVX1 U248 ( .A(n129), .Y(n130) );
  AND2X2 U249 ( .A(\mem<22><10> ), .B(n228), .Y(n131) );
  INVX1 U250 ( .A(n131), .Y(n132) );
  AND2X2 U251 ( .A(\mem<22><11> ), .B(n228), .Y(n133) );
  INVX1 U252 ( .A(n133), .Y(n134) );
  AND2X2 U253 ( .A(\mem<22><12> ), .B(n228), .Y(n135) );
  INVX1 U254 ( .A(n135), .Y(n136) );
  AND2X2 U255 ( .A(\mem<22><13> ), .B(n228), .Y(n137) );
  INVX1 U256 ( .A(n137), .Y(n138) );
  AND2X2 U257 ( .A(\mem<22><14> ), .B(n228), .Y(n139) );
  INVX1 U258 ( .A(n139), .Y(n140) );
  AND2X2 U259 ( .A(\mem<21><8> ), .B(n230), .Y(n141) );
  INVX1 U260 ( .A(n141), .Y(n142) );
  AND2X2 U261 ( .A(\mem<21><9> ), .B(n230), .Y(n143) );
  INVX1 U262 ( .A(n143), .Y(n144) );
  AND2X2 U263 ( .A(\mem<21><10> ), .B(n230), .Y(n145) );
  INVX1 U264 ( .A(n145), .Y(n146) );
  AND2X2 U265 ( .A(\mem<21><11> ), .B(n230), .Y(n147) );
  INVX1 U266 ( .A(n147), .Y(n148) );
  AND2X2 U267 ( .A(\mem<21><12> ), .B(n230), .Y(n149) );
  INVX1 U268 ( .A(n149), .Y(n150) );
  AND2X2 U269 ( .A(\mem<21><13> ), .B(n230), .Y(n151) );
  INVX1 U270 ( .A(n151), .Y(n152) );
  AND2X2 U271 ( .A(\mem<21><14> ), .B(n230), .Y(n153) );
  INVX1 U272 ( .A(n153), .Y(n154) );
  AND2X2 U273 ( .A(\mem<20><8> ), .B(n232), .Y(n155) );
  INVX1 U274 ( .A(n155), .Y(n156) );
  AND2X2 U275 ( .A(\mem<20><9> ), .B(n232), .Y(n157) );
  INVX1 U276 ( .A(n157), .Y(n158) );
  AND2X2 U277 ( .A(\mem<20><10> ), .B(n232), .Y(n159) );
  INVX1 U278 ( .A(n159), .Y(n160) );
  AND2X2 U279 ( .A(\mem<20><11> ), .B(n232), .Y(n161) );
  INVX1 U280 ( .A(n161), .Y(n162) );
  AND2X2 U281 ( .A(\mem<20><12> ), .B(n232), .Y(n163) );
  INVX1 U282 ( .A(n163), .Y(n164) );
  AND2X2 U283 ( .A(\mem<20><13> ), .B(n232), .Y(n165) );
  INVX1 U284 ( .A(n165), .Y(n166) );
  AND2X2 U285 ( .A(\mem<20><14> ), .B(n232), .Y(n167) );
  INVX1 U286 ( .A(n167), .Y(n168) );
  AND2X2 U287 ( .A(\mem<7><7> ), .B(n259), .Y(n169) );
  INVX1 U288 ( .A(n169), .Y(n170) );
  AND2X2 U289 ( .A(\mem<6><7> ), .B(n261), .Y(n171) );
  INVX1 U290 ( .A(n171), .Y(n172) );
  AND2X2 U291 ( .A(\mem<5><7> ), .B(n263), .Y(n173) );
  INVX1 U292 ( .A(n173), .Y(n174) );
  AND2X2 U293 ( .A(\mem<4><7> ), .B(n265), .Y(n175) );
  INVX1 U294 ( .A(n175), .Y(n176) );
  AND2X2 U295 ( .A(\mem<3><7> ), .B(n267), .Y(n177) );
  INVX1 U296 ( .A(n177), .Y(n178) );
  AND2X2 U297 ( .A(\mem<2><7> ), .B(n269), .Y(n179) );
  INVX1 U298 ( .A(n179), .Y(n180) );
  AND2X2 U299 ( .A(\mem<1><7> ), .B(n271), .Y(n181) );
  INVX1 U300 ( .A(n181), .Y(n182) );
  INVX4 U301 ( .A(n208), .Y(n209) );
  INVX4 U302 ( .A(n210), .Y(n211) );
  INVX4 U303 ( .A(n212), .Y(n213) );
  INVX4 U304 ( .A(n215), .Y(n216) );
  INVX4 U305 ( .A(n217), .Y(n218) );
  INVX4 U306 ( .A(n219), .Y(n220) );
  INVX4 U307 ( .A(n221), .Y(n222) );
  INVX4 U308 ( .A(n223), .Y(n224) );
  INVX4 U309 ( .A(n225), .Y(n226) );
  INVX4 U310 ( .A(n227), .Y(n228) );
  INVX4 U311 ( .A(n229), .Y(n230) );
  INVX4 U312 ( .A(n231), .Y(n232) );
  AND2X2 U313 ( .A(n2074), .B(n1410), .Y(n183) );
  INVX1 U314 ( .A(n183), .Y(n184) );
  AND2X2 U315 ( .A(n2074), .B(n1412), .Y(n185) );
  AND2X2 U316 ( .A(n2074), .B(n1414), .Y(n187) );
  AND2X2 U317 ( .A(n2074), .B(n1385), .Y(n189) );
  AND2X2 U318 ( .A(n2074), .B(n1416), .Y(n191) );
  AND2X2 U319 ( .A(n2074), .B(n1418), .Y(n193) );
  AND2X2 U320 ( .A(n2074), .B(n1420), .Y(n195) );
  AND2X2 U321 ( .A(n2074), .B(n1422), .Y(n197) );
  AND2X2 U322 ( .A(n2074), .B(n1424), .Y(n199) );
  AND2X2 U323 ( .A(n2074), .B(n1426), .Y(n201) );
  AND2X2 U324 ( .A(n2074), .B(n1428), .Y(n203) );
  AND2X2 U325 ( .A(n2074), .B(n1387), .Y(n205) );
  INVX1 U326 ( .A(n233), .Y(n207) );
  AND2X2 U327 ( .A(n2075), .B(n1388), .Y(n208) );
  AND2X2 U328 ( .A(n2075), .B(n1390), .Y(n210) );
  AND2X2 U329 ( .A(n2075), .B(n1392), .Y(n212) );
  AND2X2 U330 ( .A(n2075), .B(n1394), .Y(n215) );
  AND2X2 U331 ( .A(n2075), .B(n1396), .Y(n217) );
  AND2X2 U332 ( .A(n2075), .B(n1398), .Y(n219) );
  AND2X2 U333 ( .A(n2075), .B(n1400), .Y(n221) );
  AND2X2 U334 ( .A(n2075), .B(n1384), .Y(n223) );
  AND2X2 U335 ( .A(n2075), .B(n1402), .Y(n225) );
  AND2X2 U336 ( .A(n2075), .B(n1404), .Y(n227) );
  AND2X2 U337 ( .A(n2075), .B(n1406), .Y(n229) );
  AND2X2 U338 ( .A(n2075), .B(n1408), .Y(n231) );
  AND2X2 U339 ( .A(\data_in<7> ), .B(n2076), .Y(n233) );
  AND2X2 U340 ( .A(\mem<19><7> ), .B(n2038), .Y(n234) );
  INVX1 U341 ( .A(n234), .Y(n235) );
  AND2X2 U342 ( .A(\mem<19><15> ), .B(n2038), .Y(n236) );
  INVX1 U343 ( .A(n236), .Y(n237) );
  AND2X2 U344 ( .A(\mem<15><15> ), .B(n192), .Y(n238) );
  INVX1 U345 ( .A(n238), .Y(n239) );
  AND2X2 U346 ( .A(\mem<14><15> ), .B(n194), .Y(n240) );
  INVX1 U347 ( .A(n240), .Y(n241) );
  AND2X2 U348 ( .A(\mem<13><15> ), .B(n196), .Y(n242) );
  INVX1 U349 ( .A(n242), .Y(n243) );
  AND2X2 U350 ( .A(\mem<12><15> ), .B(n198), .Y(n244) );
  INVX1 U351 ( .A(n244), .Y(n245) );
  AND2X2 U352 ( .A(\mem<11><15> ), .B(n200), .Y(n246) );
  INVX1 U353 ( .A(n246), .Y(n247) );
  AND2X2 U354 ( .A(\mem<10><15> ), .B(n202), .Y(n248) );
  INVX1 U355 ( .A(n248), .Y(n249) );
  AND2X2 U356 ( .A(\mem<9><15> ), .B(n204), .Y(n250) );
  INVX1 U357 ( .A(n250), .Y(n251) );
  AND2X2 U358 ( .A(\mem<8><7> ), .B(n257), .Y(n252) );
  INVX1 U359 ( .A(n252), .Y(n253) );
  AND2X2 U360 ( .A(\mem<8><15> ), .B(n257), .Y(n254) );
  INVX1 U361 ( .A(n254), .Y(n255) );
  AND2X2 U362 ( .A(n2075), .B(n1386), .Y(n256) );
  AND2X2 U363 ( .A(n2075), .B(n1430), .Y(n258) );
  AND2X2 U364 ( .A(n2075), .B(n1432), .Y(n260) );
  AND2X2 U365 ( .A(n2075), .B(n1434), .Y(n262) );
  AND2X2 U366 ( .A(n2075), .B(n1436), .Y(n264) );
  AND2X2 U367 ( .A(n2075), .B(n1438), .Y(n266) );
  AND2X2 U368 ( .A(n2075), .B(n1440), .Y(n268) );
  AND2X2 U369 ( .A(n2075), .B(n1442), .Y(n270) );
  INVX1 U370 ( .A(n274), .Y(n272) );
  INVX1 U371 ( .A(n274), .Y(n273) );
  AND2X2 U372 ( .A(\data_in<15> ), .B(n2075), .Y(n274) );
  INVX1 U373 ( .A(n233), .Y(n275) );
  INVX1 U374 ( .A(n274), .Y(n276) );
  AND2X2 U375 ( .A(\data_in<0> ), .B(n2076), .Y(n277) );
  AND2X2 U376 ( .A(\data_in<1> ), .B(n2076), .Y(n278) );
  AND2X2 U377 ( .A(\data_in<2> ), .B(n2076), .Y(n279) );
  AND2X2 U378 ( .A(\data_in<3> ), .B(n2076), .Y(n280) );
  AND2X2 U379 ( .A(\data_in<4> ), .B(n2076), .Y(n281) );
  AND2X2 U380 ( .A(\data_in<5> ), .B(n2076), .Y(n282) );
  AND2X2 U381 ( .A(\data_in<6> ), .B(n2076), .Y(n283) );
  AND2X2 U382 ( .A(\data_in<8> ), .B(n2076), .Y(n284) );
  AND2X2 U383 ( .A(\data_in<9> ), .B(n2076), .Y(n285) );
  AND2X2 U384 ( .A(\data_in<10> ), .B(n2076), .Y(n286) );
  AND2X2 U385 ( .A(\data_in<11> ), .B(n2075), .Y(n287) );
  AND2X2 U386 ( .A(\data_in<12> ), .B(n2075), .Y(n288) );
  AND2X2 U387 ( .A(\data_in<13> ), .B(n2075), .Y(n289) );
  AND2X2 U388 ( .A(\data_in<14> ), .B(n2075), .Y(n290) );
  AND2X2 U389 ( .A(write), .B(n2107), .Y(n291) );
  AND2X2 U390 ( .A(n1469), .B(n2107), .Y(n292) );
  AND2X2 U391 ( .A(\mem<4><15> ), .B(n265), .Y(n293) );
  INVX1 U392 ( .A(n293), .Y(n294) );
  INVX1 U393 ( .A(n2109), .Y(n2108) );
  AND2X1 U394 ( .A(n2112), .B(n2110), .Y(n295) );
  INVX1 U395 ( .A(n2111), .Y(n2110) );
  INVX1 U396 ( .A(n2113), .Y(n2112) );
  AND2X1 U397 ( .A(n2773), .B(N14), .Y(n296) );
  AND2X2 U398 ( .A(\mem<19><0> ), .B(n2038), .Y(n297) );
  INVX1 U399 ( .A(n297), .Y(n298) );
  AND2X2 U400 ( .A(\mem<19><1> ), .B(n2038), .Y(n299) );
  INVX1 U401 ( .A(n299), .Y(n300) );
  AND2X2 U402 ( .A(\mem<19><2> ), .B(n2038), .Y(n301) );
  INVX1 U403 ( .A(n301), .Y(n302) );
  AND2X2 U404 ( .A(\mem<19><3> ), .B(n2038), .Y(n303) );
  INVX1 U405 ( .A(n303), .Y(n304) );
  AND2X2 U406 ( .A(\mem<19><4> ), .B(n2038), .Y(n305) );
  INVX1 U407 ( .A(n305), .Y(n306) );
  AND2X2 U408 ( .A(\mem<19><5> ), .B(n2038), .Y(n307) );
  INVX1 U409 ( .A(n307), .Y(n308) );
  AND2X2 U410 ( .A(\mem<19><6> ), .B(n2038), .Y(n309) );
  INVX1 U411 ( .A(n309), .Y(n310) );
  AND2X2 U412 ( .A(\mem<19><8> ), .B(n2038), .Y(n311) );
  INVX1 U413 ( .A(n311), .Y(n312) );
  AND2X2 U414 ( .A(\mem<19><9> ), .B(n2038), .Y(n313) );
  INVX1 U415 ( .A(n313), .Y(n314) );
  AND2X2 U416 ( .A(\mem<19><10> ), .B(n2038), .Y(n315) );
  INVX1 U417 ( .A(n315), .Y(n316) );
  AND2X2 U418 ( .A(\mem<19><11> ), .B(n2038), .Y(n317) );
  INVX1 U419 ( .A(n317), .Y(n318) );
  AND2X2 U420 ( .A(\mem<19><12> ), .B(n2038), .Y(n319) );
  INVX1 U421 ( .A(n319), .Y(n320) );
  AND2X2 U422 ( .A(\mem<19><13> ), .B(n2038), .Y(n321) );
  INVX1 U423 ( .A(n321), .Y(n322) );
  AND2X2 U424 ( .A(\mem<19><14> ), .B(n2038), .Y(n323) );
  INVX1 U425 ( .A(n323), .Y(n324) );
  AND2X2 U426 ( .A(\mem<18><0> ), .B(n186), .Y(n325) );
  INVX1 U427 ( .A(n325), .Y(n326) );
  AND2X2 U428 ( .A(\mem<18><1> ), .B(n186), .Y(n327) );
  INVX1 U429 ( .A(n327), .Y(n328) );
  AND2X2 U430 ( .A(\mem<18><2> ), .B(n186), .Y(n329) );
  INVX1 U431 ( .A(n329), .Y(n330) );
  AND2X2 U432 ( .A(\mem<18><3> ), .B(n186), .Y(n331) );
  INVX1 U433 ( .A(n331), .Y(n332) );
  AND2X2 U434 ( .A(\mem<18><4> ), .B(n186), .Y(n333) );
  INVX1 U435 ( .A(n333), .Y(n334) );
  AND2X2 U436 ( .A(\mem<18><5> ), .B(n186), .Y(n335) );
  INVX1 U437 ( .A(n335), .Y(n336) );
  AND2X2 U438 ( .A(\mem<18><6> ), .B(n186), .Y(n337) );
  INVX1 U439 ( .A(n337), .Y(n338) );
  AND2X2 U440 ( .A(\mem<18><8> ), .B(n186), .Y(n339) );
  INVX1 U441 ( .A(n339), .Y(n340) );
  AND2X2 U442 ( .A(\mem<18><9> ), .B(n186), .Y(n341) );
  INVX1 U443 ( .A(n341), .Y(n342) );
  AND2X2 U444 ( .A(\mem<18><10> ), .B(n186), .Y(n343) );
  INVX1 U445 ( .A(n343), .Y(n344) );
  AND2X2 U446 ( .A(\mem<18><11> ), .B(n186), .Y(n345) );
  INVX1 U447 ( .A(n345), .Y(n346) );
  AND2X2 U448 ( .A(\mem<18><12> ), .B(n186), .Y(n347) );
  INVX1 U449 ( .A(n347), .Y(n348) );
  AND2X2 U450 ( .A(\mem<18><13> ), .B(n186), .Y(n349) );
  INVX1 U451 ( .A(n349), .Y(n350) );
  AND2X2 U452 ( .A(\mem<18><14> ), .B(n186), .Y(n351) );
  INVX1 U453 ( .A(n351), .Y(n352) );
  AND2X2 U454 ( .A(\mem<18><15> ), .B(n186), .Y(n353) );
  INVX1 U455 ( .A(n353), .Y(n354) );
  AND2X2 U456 ( .A(\mem<17><0> ), .B(n188), .Y(n355) );
  INVX1 U457 ( .A(n355), .Y(n356) );
  AND2X2 U458 ( .A(\mem<17><1> ), .B(n188), .Y(n357) );
  INVX1 U459 ( .A(n357), .Y(n358) );
  AND2X2 U460 ( .A(\mem<17><2> ), .B(n188), .Y(n359) );
  INVX1 U461 ( .A(n359), .Y(n360) );
  AND2X2 U462 ( .A(\mem<17><3> ), .B(n188), .Y(n361) );
  INVX1 U463 ( .A(n361), .Y(n362) );
  AND2X2 U464 ( .A(\mem<17><4> ), .B(n188), .Y(n363) );
  INVX1 U465 ( .A(n363), .Y(n364) );
  AND2X2 U466 ( .A(\mem<17><5> ), .B(n188), .Y(n365) );
  INVX1 U467 ( .A(n365), .Y(n366) );
  AND2X2 U468 ( .A(\mem<17><6> ), .B(n188), .Y(n367) );
  INVX1 U469 ( .A(n367), .Y(n368) );
  AND2X2 U470 ( .A(\mem<17><8> ), .B(n188), .Y(n369) );
  INVX1 U471 ( .A(n369), .Y(n370) );
  AND2X2 U472 ( .A(\mem<17><9> ), .B(n188), .Y(n371) );
  INVX1 U473 ( .A(n371), .Y(n372) );
  AND2X2 U474 ( .A(\mem<17><10> ), .B(n188), .Y(n373) );
  INVX1 U475 ( .A(n373), .Y(n374) );
  AND2X2 U476 ( .A(\mem<17><11> ), .B(n188), .Y(n375) );
  INVX1 U477 ( .A(n375), .Y(n376) );
  AND2X2 U478 ( .A(\mem<17><12> ), .B(n188), .Y(n377) );
  INVX1 U479 ( .A(n377), .Y(n378) );
  AND2X2 U480 ( .A(\mem<17><13> ), .B(n188), .Y(n379) );
  INVX1 U481 ( .A(n379), .Y(n380) );
  AND2X2 U482 ( .A(\mem<17><14> ), .B(n188), .Y(n381) );
  INVX1 U483 ( .A(n381), .Y(n382) );
  AND2X2 U484 ( .A(\mem<17><15> ), .B(n188), .Y(n383) );
  INVX1 U485 ( .A(n383), .Y(n384) );
  AND2X2 U486 ( .A(\mem<16><0> ), .B(n190), .Y(n385) );
  INVX1 U487 ( .A(n385), .Y(n386) );
  AND2X2 U488 ( .A(\mem<16><1> ), .B(n190), .Y(n387) );
  INVX1 U489 ( .A(n387), .Y(n388) );
  AND2X2 U490 ( .A(\mem<16><2> ), .B(n190), .Y(n389) );
  INVX1 U491 ( .A(n389), .Y(n390) );
  AND2X2 U492 ( .A(\mem<16><3> ), .B(n190), .Y(n391) );
  INVX1 U493 ( .A(n391), .Y(n392) );
  AND2X2 U494 ( .A(\mem<16><4> ), .B(n190), .Y(n393) );
  INVX1 U495 ( .A(n393), .Y(n394) );
  AND2X2 U496 ( .A(\mem<16><5> ), .B(n190), .Y(n395) );
  INVX1 U497 ( .A(n395), .Y(n396) );
  AND2X2 U498 ( .A(\mem<16><6> ), .B(n190), .Y(n397) );
  INVX1 U499 ( .A(n397), .Y(n398) );
  AND2X2 U500 ( .A(\mem<16><8> ), .B(n190), .Y(n399) );
  INVX1 U501 ( .A(n399), .Y(n400) );
  AND2X2 U502 ( .A(\mem<16><9> ), .B(n190), .Y(n401) );
  INVX1 U503 ( .A(n401), .Y(n402) );
  AND2X2 U504 ( .A(\mem<16><10> ), .B(n190), .Y(n403) );
  INVX1 U505 ( .A(n403), .Y(n404) );
  AND2X2 U506 ( .A(\mem<16><11> ), .B(n190), .Y(n405) );
  INVX1 U507 ( .A(n405), .Y(n406) );
  AND2X2 U508 ( .A(\mem<16><12> ), .B(n190), .Y(n407) );
  INVX1 U509 ( .A(n407), .Y(n408) );
  AND2X2 U510 ( .A(\mem<16><13> ), .B(n190), .Y(n409) );
  INVX1 U511 ( .A(n409), .Y(n410) );
  AND2X2 U512 ( .A(\mem<16><14> ), .B(n190), .Y(n411) );
  INVX1 U513 ( .A(n411), .Y(n412) );
  AND2X2 U514 ( .A(\mem<15><0> ), .B(n192), .Y(n413) );
  INVX1 U515 ( .A(n413), .Y(n414) );
  AND2X2 U516 ( .A(\mem<15><1> ), .B(n192), .Y(n415) );
  INVX1 U517 ( .A(n415), .Y(n416) );
  AND2X2 U518 ( .A(\mem<15><2> ), .B(n192), .Y(n417) );
  INVX1 U519 ( .A(n417), .Y(n418) );
  AND2X2 U520 ( .A(\mem<15><3> ), .B(n192), .Y(n419) );
  INVX1 U521 ( .A(n419), .Y(n420) );
  AND2X2 U522 ( .A(\mem<15><4> ), .B(n192), .Y(n421) );
  INVX1 U523 ( .A(n421), .Y(n422) );
  AND2X2 U524 ( .A(\mem<15><5> ), .B(n192), .Y(n423) );
  INVX1 U525 ( .A(n423), .Y(n424) );
  AND2X2 U526 ( .A(\mem<15><6> ), .B(n192), .Y(n425) );
  INVX1 U527 ( .A(n425), .Y(n426) );
  AND2X2 U528 ( .A(\mem<15><8> ), .B(n192), .Y(n427) );
  INVX1 U529 ( .A(n427), .Y(n428) );
  AND2X2 U530 ( .A(\mem<15><9> ), .B(n192), .Y(n429) );
  INVX1 U531 ( .A(n429), .Y(n430) );
  AND2X2 U532 ( .A(\mem<15><10> ), .B(n192), .Y(n431) );
  INVX1 U533 ( .A(n431), .Y(n432) );
  AND2X2 U534 ( .A(\mem<15><11> ), .B(n192), .Y(n433) );
  INVX1 U535 ( .A(n433), .Y(n434) );
  AND2X2 U536 ( .A(\mem<15><12> ), .B(n192), .Y(n435) );
  INVX1 U537 ( .A(n435), .Y(n436) );
  AND2X2 U538 ( .A(\mem<15><13> ), .B(n192), .Y(n437) );
  INVX1 U539 ( .A(n437), .Y(n438) );
  AND2X2 U540 ( .A(\mem<15><14> ), .B(n192), .Y(n439) );
  INVX1 U541 ( .A(n439), .Y(n440) );
  AND2X2 U542 ( .A(\mem<14><0> ), .B(n194), .Y(n441) );
  INVX1 U543 ( .A(n441), .Y(n442) );
  AND2X2 U544 ( .A(\mem<14><1> ), .B(n194), .Y(n443) );
  INVX1 U545 ( .A(n443), .Y(n444) );
  AND2X2 U546 ( .A(\mem<14><2> ), .B(n194), .Y(n445) );
  INVX1 U547 ( .A(n445), .Y(n446) );
  AND2X2 U548 ( .A(\mem<14><3> ), .B(n194), .Y(n447) );
  INVX1 U549 ( .A(n447), .Y(n448) );
  AND2X2 U550 ( .A(\mem<14><4> ), .B(n194), .Y(n449) );
  INVX1 U551 ( .A(n449), .Y(n450) );
  AND2X2 U552 ( .A(\mem<14><5> ), .B(n194), .Y(n451) );
  INVX1 U553 ( .A(n451), .Y(n452) );
  AND2X2 U554 ( .A(\mem<14><6> ), .B(n194), .Y(n453) );
  INVX1 U555 ( .A(n453), .Y(n454) );
  AND2X2 U556 ( .A(\mem<14><8> ), .B(n194), .Y(n455) );
  INVX1 U557 ( .A(n455), .Y(n456) );
  AND2X2 U558 ( .A(\mem<14><9> ), .B(n194), .Y(n457) );
  INVX1 U559 ( .A(n457), .Y(n458) );
  AND2X2 U560 ( .A(\mem<14><10> ), .B(n194), .Y(n459) );
  INVX1 U561 ( .A(n459), .Y(n460) );
  AND2X2 U562 ( .A(\mem<14><11> ), .B(n194), .Y(n461) );
  INVX1 U563 ( .A(n461), .Y(n462) );
  AND2X2 U564 ( .A(\mem<14><12> ), .B(n194), .Y(n463) );
  INVX1 U565 ( .A(n463), .Y(n464) );
  AND2X2 U566 ( .A(\mem<14><13> ), .B(n194), .Y(n465) );
  INVX1 U567 ( .A(n465), .Y(n466) );
  AND2X2 U568 ( .A(\mem<14><14> ), .B(n194), .Y(n467) );
  INVX1 U569 ( .A(n467), .Y(n468) );
  AND2X2 U570 ( .A(\mem<13><0> ), .B(n196), .Y(n469) );
  INVX1 U571 ( .A(n469), .Y(n470) );
  AND2X2 U572 ( .A(\mem<13><1> ), .B(n196), .Y(n471) );
  INVX1 U573 ( .A(n471), .Y(n472) );
  AND2X2 U574 ( .A(\mem<13><2> ), .B(n196), .Y(n473) );
  INVX1 U575 ( .A(n473), .Y(n474) );
  AND2X2 U576 ( .A(\mem<13><3> ), .B(n196), .Y(n475) );
  INVX1 U577 ( .A(n475), .Y(n476) );
  AND2X2 U578 ( .A(\mem<13><4> ), .B(n196), .Y(n477) );
  INVX1 U579 ( .A(n477), .Y(n478) );
  AND2X2 U580 ( .A(\mem<13><5> ), .B(n196), .Y(n479) );
  INVX1 U581 ( .A(n479), .Y(n480) );
  AND2X2 U582 ( .A(\mem<13><6> ), .B(n196), .Y(n481) );
  INVX1 U583 ( .A(n481), .Y(n482) );
  AND2X2 U584 ( .A(\mem<13><8> ), .B(n196), .Y(n483) );
  INVX1 U585 ( .A(n483), .Y(n484) );
  AND2X2 U586 ( .A(\mem<13><9> ), .B(n196), .Y(n485) );
  INVX1 U587 ( .A(n485), .Y(n486) );
  AND2X2 U588 ( .A(\mem<13><10> ), .B(n196), .Y(n487) );
  INVX1 U589 ( .A(n487), .Y(n488) );
  AND2X2 U590 ( .A(\mem<13><11> ), .B(n196), .Y(n489) );
  INVX1 U591 ( .A(n489), .Y(n490) );
  AND2X2 U592 ( .A(\mem<13><12> ), .B(n196), .Y(n491) );
  INVX1 U593 ( .A(n491), .Y(n492) );
  AND2X2 U594 ( .A(\mem<13><13> ), .B(n196), .Y(n493) );
  INVX1 U595 ( .A(n493), .Y(n494) );
  AND2X2 U596 ( .A(\mem<13><14> ), .B(n196), .Y(n495) );
  INVX1 U597 ( .A(n495), .Y(n496) );
  AND2X2 U598 ( .A(\mem<12><0> ), .B(n198), .Y(n497) );
  INVX1 U599 ( .A(n497), .Y(n498) );
  AND2X2 U600 ( .A(\mem<12><1> ), .B(n198), .Y(n499) );
  INVX1 U601 ( .A(n499), .Y(n500) );
  AND2X2 U602 ( .A(\mem<12><2> ), .B(n198), .Y(n501) );
  INVX1 U603 ( .A(n501), .Y(n502) );
  AND2X2 U604 ( .A(\mem<12><3> ), .B(n198), .Y(n503) );
  INVX1 U605 ( .A(n503), .Y(n504) );
  AND2X2 U606 ( .A(\mem<12><4> ), .B(n198), .Y(n505) );
  INVX1 U607 ( .A(n505), .Y(n506) );
  AND2X2 U608 ( .A(\mem<12><5> ), .B(n198), .Y(n507) );
  INVX1 U609 ( .A(n507), .Y(n508) );
  AND2X2 U610 ( .A(\mem<12><6> ), .B(n198), .Y(n509) );
  INVX1 U611 ( .A(n509), .Y(n510) );
  AND2X2 U612 ( .A(\mem<12><8> ), .B(n198), .Y(n511) );
  INVX1 U613 ( .A(n511), .Y(n512) );
  AND2X2 U614 ( .A(\mem<12><9> ), .B(n198), .Y(n513) );
  INVX1 U615 ( .A(n513), .Y(n514) );
  AND2X2 U616 ( .A(\mem<12><10> ), .B(n198), .Y(n515) );
  INVX1 U617 ( .A(n515), .Y(n516) );
  AND2X2 U618 ( .A(\mem<12><11> ), .B(n198), .Y(n517) );
  INVX1 U619 ( .A(n517), .Y(n518) );
  AND2X2 U620 ( .A(\mem<12><12> ), .B(n198), .Y(n519) );
  INVX1 U621 ( .A(n519), .Y(n520) );
  AND2X2 U622 ( .A(\mem<12><13> ), .B(n198), .Y(n521) );
  INVX1 U623 ( .A(n521), .Y(n522) );
  AND2X2 U624 ( .A(\mem<12><14> ), .B(n198), .Y(n523) );
  INVX1 U625 ( .A(n523), .Y(n524) );
  AND2X2 U626 ( .A(\mem<11><0> ), .B(n200), .Y(n525) );
  INVX1 U627 ( .A(n525), .Y(n526) );
  AND2X2 U628 ( .A(\mem<11><1> ), .B(n200), .Y(n527) );
  INVX1 U629 ( .A(n527), .Y(n528) );
  AND2X2 U630 ( .A(\mem<11><2> ), .B(n200), .Y(n529) );
  INVX1 U631 ( .A(n529), .Y(n530) );
  AND2X2 U632 ( .A(\mem<11><3> ), .B(n200), .Y(n531) );
  INVX1 U633 ( .A(n531), .Y(n532) );
  AND2X2 U634 ( .A(\mem<11><4> ), .B(n200), .Y(n533) );
  INVX1 U635 ( .A(n533), .Y(n534) );
  AND2X2 U636 ( .A(\mem<11><5> ), .B(n200), .Y(n535) );
  INVX1 U637 ( .A(n535), .Y(n536) );
  AND2X2 U638 ( .A(\mem<11><6> ), .B(n200), .Y(n537) );
  INVX1 U639 ( .A(n537), .Y(n538) );
  AND2X2 U640 ( .A(\mem<11><8> ), .B(n200), .Y(n539) );
  INVX1 U641 ( .A(n539), .Y(n540) );
  AND2X2 U642 ( .A(\mem<11><9> ), .B(n200), .Y(n541) );
  INVX1 U643 ( .A(n541), .Y(n542) );
  AND2X2 U644 ( .A(\mem<11><10> ), .B(n200), .Y(n543) );
  INVX1 U645 ( .A(n543), .Y(n544) );
  AND2X2 U646 ( .A(\mem<11><11> ), .B(n200), .Y(n545) );
  INVX1 U647 ( .A(n545), .Y(n546) );
  AND2X2 U648 ( .A(\mem<11><12> ), .B(n200), .Y(n547) );
  INVX1 U649 ( .A(n547), .Y(n548) );
  AND2X2 U650 ( .A(\mem<11><13> ), .B(n200), .Y(n549) );
  INVX1 U651 ( .A(n549), .Y(n550) );
  AND2X2 U652 ( .A(\mem<11><14> ), .B(n200), .Y(n551) );
  INVX1 U653 ( .A(n551), .Y(n552) );
  AND2X2 U654 ( .A(\mem<10><0> ), .B(n202), .Y(n553) );
  INVX1 U655 ( .A(n553), .Y(n554) );
  AND2X2 U656 ( .A(\mem<10><1> ), .B(n202), .Y(n555) );
  INVX1 U657 ( .A(n555), .Y(n556) );
  AND2X2 U658 ( .A(\mem<10><2> ), .B(n202), .Y(n557) );
  INVX1 U659 ( .A(n557), .Y(n558) );
  AND2X2 U660 ( .A(\mem<10><3> ), .B(n202), .Y(n559) );
  INVX1 U661 ( .A(n559), .Y(n560) );
  AND2X2 U662 ( .A(\mem<10><4> ), .B(n202), .Y(n561) );
  INVX1 U663 ( .A(n561), .Y(n562) );
  AND2X2 U664 ( .A(\mem<10><5> ), .B(n202), .Y(n563) );
  INVX1 U665 ( .A(n563), .Y(n564) );
  AND2X2 U666 ( .A(\mem<10><6> ), .B(n202), .Y(n565) );
  INVX1 U667 ( .A(n565), .Y(n566) );
  AND2X2 U668 ( .A(\mem<10><8> ), .B(n202), .Y(n567) );
  INVX1 U669 ( .A(n567), .Y(n568) );
  AND2X2 U670 ( .A(\mem<10><9> ), .B(n202), .Y(n569) );
  INVX1 U671 ( .A(n569), .Y(n570) );
  AND2X2 U672 ( .A(\mem<10><10> ), .B(n202), .Y(n571) );
  INVX1 U673 ( .A(n571), .Y(n572) );
  AND2X2 U674 ( .A(\mem<10><11> ), .B(n202), .Y(n573) );
  INVX1 U675 ( .A(n573), .Y(n574) );
  AND2X2 U676 ( .A(\mem<10><12> ), .B(n202), .Y(n575) );
  INVX1 U677 ( .A(n575), .Y(n576) );
  AND2X2 U678 ( .A(\mem<10><13> ), .B(n202), .Y(n577) );
  INVX1 U679 ( .A(n577), .Y(n578) );
  AND2X2 U680 ( .A(\mem<10><14> ), .B(n202), .Y(n579) );
  INVX1 U681 ( .A(n579), .Y(n580) );
  AND2X2 U682 ( .A(\mem<9><0> ), .B(n204), .Y(n581) );
  INVX1 U683 ( .A(n581), .Y(n582) );
  AND2X2 U684 ( .A(\mem<9><1> ), .B(n204), .Y(n583) );
  INVX1 U685 ( .A(n583), .Y(n584) );
  AND2X2 U686 ( .A(\mem<9><2> ), .B(n204), .Y(n585) );
  INVX1 U687 ( .A(n585), .Y(n586) );
  AND2X2 U688 ( .A(\mem<9><3> ), .B(n204), .Y(n587) );
  INVX1 U689 ( .A(n587), .Y(n588) );
  AND2X2 U690 ( .A(\mem<9><4> ), .B(n204), .Y(n589) );
  INVX1 U691 ( .A(n589), .Y(n590) );
  AND2X2 U692 ( .A(\mem<9><5> ), .B(n204), .Y(n591) );
  INVX1 U693 ( .A(n591), .Y(n592) );
  AND2X2 U694 ( .A(\mem<9><6> ), .B(n204), .Y(n593) );
  INVX1 U695 ( .A(n593), .Y(n594) );
  AND2X2 U696 ( .A(\mem<9><8> ), .B(n204), .Y(n595) );
  INVX1 U697 ( .A(n595), .Y(n596) );
  AND2X2 U698 ( .A(\mem<9><9> ), .B(n204), .Y(n597) );
  INVX1 U699 ( .A(n597), .Y(n598) );
  AND2X2 U700 ( .A(\mem<9><10> ), .B(n204), .Y(n599) );
  INVX1 U701 ( .A(n599), .Y(n600) );
  AND2X2 U702 ( .A(\mem<9><11> ), .B(n204), .Y(n601) );
  INVX1 U703 ( .A(n601), .Y(n602) );
  AND2X2 U704 ( .A(\mem<9><12> ), .B(n204), .Y(n603) );
  INVX1 U705 ( .A(n603), .Y(n604) );
  AND2X2 U706 ( .A(\mem<9><13> ), .B(n204), .Y(n605) );
  INVX1 U707 ( .A(n605), .Y(n606) );
  AND2X2 U708 ( .A(\mem<9><14> ), .B(n204), .Y(n607) );
  INVX1 U709 ( .A(n607), .Y(n608) );
  AND2X2 U710 ( .A(\mem<8><0> ), .B(n257), .Y(n609) );
  INVX1 U711 ( .A(n609), .Y(n610) );
  AND2X2 U712 ( .A(\mem<8><1> ), .B(n257), .Y(n611) );
  INVX1 U713 ( .A(n611), .Y(n612) );
  AND2X2 U714 ( .A(\mem<8><2> ), .B(n257), .Y(n613) );
  INVX1 U715 ( .A(n613), .Y(n614) );
  AND2X2 U716 ( .A(\mem<8><3> ), .B(n257), .Y(n615) );
  INVX1 U717 ( .A(n615), .Y(n616) );
  AND2X2 U718 ( .A(\mem<8><4> ), .B(n257), .Y(n617) );
  INVX1 U719 ( .A(n617), .Y(n618) );
  AND2X2 U720 ( .A(\mem<8><5> ), .B(n257), .Y(n619) );
  INVX1 U721 ( .A(n619), .Y(n620) );
  AND2X2 U722 ( .A(\mem<8><6> ), .B(n257), .Y(n621) );
  INVX1 U723 ( .A(n621), .Y(n622) );
  AND2X2 U724 ( .A(\mem<8><8> ), .B(n257), .Y(n623) );
  INVX1 U725 ( .A(n623), .Y(n624) );
  AND2X2 U726 ( .A(\mem<8><9> ), .B(n257), .Y(n625) );
  INVX1 U727 ( .A(n625), .Y(n626) );
  AND2X2 U728 ( .A(\mem<8><10> ), .B(n257), .Y(n627) );
  INVX1 U729 ( .A(n627), .Y(n628) );
  AND2X2 U730 ( .A(\mem<8><11> ), .B(n257), .Y(n629) );
  INVX1 U731 ( .A(n629), .Y(n630) );
  AND2X2 U732 ( .A(\mem<8><12> ), .B(n257), .Y(n631) );
  INVX1 U733 ( .A(n631), .Y(n632) );
  AND2X2 U734 ( .A(\mem<8><13> ), .B(n257), .Y(n633) );
  INVX1 U735 ( .A(n633), .Y(n634) );
  AND2X2 U736 ( .A(\mem<8><14> ), .B(n257), .Y(n635) );
  INVX1 U737 ( .A(n635), .Y(n636) );
  AND2X2 U738 ( .A(\mem<7><0> ), .B(n259), .Y(n637) );
  INVX1 U739 ( .A(n637), .Y(n638) );
  AND2X2 U740 ( .A(\mem<7><1> ), .B(n259), .Y(n639) );
  INVX1 U741 ( .A(n639), .Y(n640) );
  AND2X2 U742 ( .A(\mem<7><2> ), .B(n259), .Y(n641) );
  INVX1 U743 ( .A(n641), .Y(n642) );
  AND2X2 U744 ( .A(\mem<7><3> ), .B(n259), .Y(n643) );
  INVX1 U745 ( .A(n643), .Y(n644) );
  AND2X2 U746 ( .A(\mem<7><4> ), .B(n259), .Y(n645) );
  INVX1 U747 ( .A(n645), .Y(n646) );
  AND2X2 U748 ( .A(\mem<7><5> ), .B(n259), .Y(n647) );
  INVX1 U749 ( .A(n647), .Y(n648) );
  AND2X2 U750 ( .A(\mem<7><6> ), .B(n259), .Y(n649) );
  INVX1 U751 ( .A(n649), .Y(n650) );
  AND2X2 U752 ( .A(\mem<7><8> ), .B(n259), .Y(n1163) );
  INVX1 U753 ( .A(n1163), .Y(n1164) );
  AND2X2 U754 ( .A(\mem<7><9> ), .B(n259), .Y(n1165) );
  INVX1 U755 ( .A(n1165), .Y(n1166) );
  AND2X2 U756 ( .A(\mem<7><10> ), .B(n259), .Y(n1167) );
  INVX1 U757 ( .A(n1167), .Y(n1168) );
  AND2X2 U758 ( .A(\mem<7><11> ), .B(n259), .Y(n1169) );
  INVX1 U759 ( .A(n1169), .Y(n1170) );
  AND2X2 U760 ( .A(\mem<7><12> ), .B(n259), .Y(n1171) );
  INVX1 U761 ( .A(n1171), .Y(n1172) );
  AND2X2 U762 ( .A(\mem<7><13> ), .B(n259), .Y(n1173) );
  INVX1 U763 ( .A(n1173), .Y(n1174) );
  AND2X2 U764 ( .A(\mem<7><14> ), .B(n259), .Y(n1175) );
  INVX1 U765 ( .A(n1175), .Y(n1176) );
  AND2X2 U766 ( .A(\mem<6><0> ), .B(n261), .Y(n1177) );
  INVX1 U767 ( .A(n1177), .Y(n1178) );
  AND2X2 U768 ( .A(\mem<6><1> ), .B(n261), .Y(n1179) );
  INVX1 U769 ( .A(n1179), .Y(n1180) );
  AND2X2 U770 ( .A(\mem<6><2> ), .B(n261), .Y(n1181) );
  INVX1 U771 ( .A(n1181), .Y(n1182) );
  AND2X2 U772 ( .A(\mem<6><3> ), .B(n261), .Y(n1183) );
  INVX1 U773 ( .A(n1183), .Y(n1184) );
  AND2X2 U774 ( .A(\mem<6><4> ), .B(n261), .Y(n1185) );
  INVX1 U775 ( .A(n1185), .Y(n1186) );
  AND2X2 U776 ( .A(\mem<6><5> ), .B(n261), .Y(n1187) );
  INVX1 U777 ( .A(n1187), .Y(n1188) );
  AND2X2 U778 ( .A(\mem<6><6> ), .B(n261), .Y(n1189) );
  INVX1 U779 ( .A(n1189), .Y(n1190) );
  AND2X2 U780 ( .A(\mem<6><8> ), .B(n261), .Y(n1191) );
  INVX1 U781 ( .A(n1191), .Y(n1192) );
  AND2X2 U782 ( .A(\mem<6><9> ), .B(n261), .Y(n1193) );
  INVX1 U783 ( .A(n1193), .Y(n1194) );
  AND2X2 U784 ( .A(\mem<6><10> ), .B(n261), .Y(n1195) );
  INVX1 U785 ( .A(n1195), .Y(n1196) );
  AND2X2 U786 ( .A(\mem<6><11> ), .B(n261), .Y(n1197) );
  INVX1 U787 ( .A(n1197), .Y(n1198) );
  AND2X2 U788 ( .A(\mem<6><12> ), .B(n261), .Y(n1199) );
  INVX1 U789 ( .A(n1199), .Y(n1200) );
  AND2X2 U790 ( .A(\mem<6><13> ), .B(n261), .Y(n1201) );
  INVX1 U791 ( .A(n1201), .Y(n1202) );
  AND2X2 U792 ( .A(\mem<6><14> ), .B(n261), .Y(n1203) );
  INVX1 U793 ( .A(n1203), .Y(n1204) );
  AND2X2 U794 ( .A(\mem<5><0> ), .B(n263), .Y(n1205) );
  INVX1 U795 ( .A(n1205), .Y(n1206) );
  AND2X2 U796 ( .A(\mem<5><1> ), .B(n263), .Y(n1207) );
  INVX1 U797 ( .A(n1207), .Y(n1208) );
  AND2X2 U798 ( .A(\mem<5><2> ), .B(n263), .Y(n1209) );
  INVX1 U799 ( .A(n1209), .Y(n1210) );
  AND2X2 U800 ( .A(\mem<5><3> ), .B(n263), .Y(n1211) );
  INVX1 U801 ( .A(n1211), .Y(n1212) );
  AND2X2 U802 ( .A(\mem<5><4> ), .B(n263), .Y(n1213) );
  INVX1 U803 ( .A(n1213), .Y(n1214) );
  AND2X2 U804 ( .A(\mem<5><5> ), .B(n263), .Y(n1215) );
  INVX1 U805 ( .A(n1215), .Y(n1216) );
  AND2X2 U806 ( .A(\mem<5><6> ), .B(n263), .Y(n1217) );
  INVX1 U807 ( .A(n1217), .Y(n1218) );
  AND2X2 U808 ( .A(\mem<5><8> ), .B(n263), .Y(n1219) );
  INVX1 U809 ( .A(n1219), .Y(n1220) );
  AND2X2 U810 ( .A(\mem<5><9> ), .B(n263), .Y(n1221) );
  INVX1 U811 ( .A(n1221), .Y(n1222) );
  AND2X2 U812 ( .A(\mem<5><10> ), .B(n263), .Y(n1223) );
  INVX1 U813 ( .A(n1223), .Y(n1224) );
  AND2X2 U814 ( .A(\mem<5><11> ), .B(n263), .Y(n1225) );
  INVX1 U815 ( .A(n1225), .Y(n1226) );
  AND2X2 U816 ( .A(\mem<5><12> ), .B(n263), .Y(n1227) );
  INVX1 U817 ( .A(n1227), .Y(n1228) );
  AND2X2 U818 ( .A(\mem<5><13> ), .B(n263), .Y(n1229) );
  INVX1 U819 ( .A(n1229), .Y(n1230) );
  AND2X2 U820 ( .A(\mem<5><14> ), .B(n263), .Y(n1231) );
  INVX1 U821 ( .A(n1231), .Y(n1232) );
  AND2X2 U822 ( .A(\mem<4><0> ), .B(n265), .Y(n1233) );
  INVX1 U823 ( .A(n1233), .Y(n1234) );
  AND2X2 U824 ( .A(\mem<4><1> ), .B(n265), .Y(n1235) );
  INVX1 U825 ( .A(n1235), .Y(n1236) );
  AND2X2 U826 ( .A(\mem<4><2> ), .B(n265), .Y(n1237) );
  INVX1 U827 ( .A(n1237), .Y(n1238) );
  AND2X2 U828 ( .A(\mem<4><3> ), .B(n265), .Y(n1239) );
  INVX1 U829 ( .A(n1239), .Y(n1240) );
  AND2X2 U830 ( .A(\mem<4><4> ), .B(n265), .Y(n1241) );
  INVX1 U831 ( .A(n1241), .Y(n1242) );
  AND2X2 U832 ( .A(\mem<4><5> ), .B(n265), .Y(n1243) );
  INVX1 U833 ( .A(n1243), .Y(n1244) );
  AND2X2 U834 ( .A(\mem<4><6> ), .B(n265), .Y(n1245) );
  INVX1 U835 ( .A(n1245), .Y(n1246) );
  AND2X2 U836 ( .A(\mem<4><8> ), .B(n265), .Y(n1247) );
  INVX1 U837 ( .A(n1247), .Y(n1248) );
  AND2X2 U838 ( .A(\mem<4><9> ), .B(n265), .Y(n1249) );
  INVX1 U839 ( .A(n1249), .Y(n1250) );
  AND2X2 U840 ( .A(\mem<4><10> ), .B(n265), .Y(n1251) );
  INVX1 U841 ( .A(n1251), .Y(n1252) );
  AND2X2 U842 ( .A(\mem<4><11> ), .B(n265), .Y(n1253) );
  INVX1 U843 ( .A(n1253), .Y(n1254) );
  AND2X2 U844 ( .A(\mem<4><12> ), .B(n265), .Y(n1255) );
  INVX1 U845 ( .A(n1255), .Y(n1256) );
  AND2X2 U846 ( .A(\mem<4><13> ), .B(n265), .Y(n1257) );
  INVX1 U847 ( .A(n1257), .Y(n1258) );
  AND2X2 U848 ( .A(\mem<4><14> ), .B(n265), .Y(n1259) );
  INVX1 U849 ( .A(n1259), .Y(n1260) );
  AND2X2 U850 ( .A(\mem<3><0> ), .B(n267), .Y(n1261) );
  INVX1 U851 ( .A(n1261), .Y(n1262) );
  AND2X2 U852 ( .A(\mem<3><1> ), .B(n267), .Y(n1263) );
  INVX1 U853 ( .A(n1263), .Y(n1264) );
  AND2X2 U854 ( .A(\mem<3><2> ), .B(n267), .Y(n1265) );
  INVX1 U855 ( .A(n1265), .Y(n1266) );
  AND2X2 U856 ( .A(\mem<3><3> ), .B(n267), .Y(n1267) );
  INVX1 U857 ( .A(n1267), .Y(n1268) );
  AND2X2 U858 ( .A(\mem<3><4> ), .B(n267), .Y(n1269) );
  INVX1 U859 ( .A(n1269), .Y(n1270) );
  AND2X2 U860 ( .A(\mem<3><5> ), .B(n267), .Y(n1271) );
  INVX1 U861 ( .A(n1271), .Y(n1272) );
  AND2X2 U862 ( .A(\mem<3><6> ), .B(n267), .Y(n1273) );
  INVX1 U863 ( .A(n1273), .Y(n1274) );
  AND2X2 U864 ( .A(\mem<3><8> ), .B(n267), .Y(n1275) );
  INVX1 U865 ( .A(n1275), .Y(n1276) );
  AND2X2 U866 ( .A(\mem<3><9> ), .B(n267), .Y(n1277) );
  INVX1 U867 ( .A(n1277), .Y(n1278) );
  AND2X2 U868 ( .A(\mem<3><10> ), .B(n267), .Y(n1279) );
  INVX1 U869 ( .A(n1279), .Y(n1280) );
  AND2X2 U870 ( .A(\mem<3><11> ), .B(n267), .Y(n1281) );
  INVX1 U871 ( .A(n1281), .Y(n1282) );
  AND2X2 U872 ( .A(\mem<3><12> ), .B(n267), .Y(n1283) );
  INVX1 U873 ( .A(n1283), .Y(n1284) );
  AND2X2 U874 ( .A(\mem<3><13> ), .B(n267), .Y(n1285) );
  INVX1 U875 ( .A(n1285), .Y(n1286) );
  AND2X2 U876 ( .A(\mem<3><14> ), .B(n267), .Y(n1287) );
  INVX1 U877 ( .A(n1287), .Y(n1288) );
  AND2X2 U878 ( .A(\mem<2><0> ), .B(n269), .Y(n1289) );
  INVX1 U879 ( .A(n1289), .Y(n1290) );
  AND2X2 U880 ( .A(\mem<2><1> ), .B(n269), .Y(n1291) );
  INVX1 U881 ( .A(n1291), .Y(n1292) );
  AND2X2 U882 ( .A(\mem<2><2> ), .B(n269), .Y(n1293) );
  INVX1 U883 ( .A(n1293), .Y(n1294) );
  AND2X2 U884 ( .A(\mem<2><3> ), .B(n269), .Y(n1295) );
  INVX1 U885 ( .A(n1295), .Y(n1296) );
  AND2X2 U886 ( .A(\mem<2><4> ), .B(n269), .Y(n1297) );
  INVX1 U887 ( .A(n1297), .Y(n1298) );
  AND2X2 U888 ( .A(\mem<2><5> ), .B(n269), .Y(n1299) );
  INVX1 U889 ( .A(n1299), .Y(n1300) );
  AND2X2 U890 ( .A(\mem<2><6> ), .B(n269), .Y(n1301) );
  INVX1 U891 ( .A(n1301), .Y(n1302) );
  AND2X2 U892 ( .A(\mem<2><8> ), .B(n269), .Y(n1303) );
  INVX1 U893 ( .A(n1303), .Y(n1304) );
  AND2X2 U894 ( .A(\mem<2><9> ), .B(n269), .Y(n1305) );
  INVX1 U895 ( .A(n1305), .Y(n1306) );
  AND2X2 U896 ( .A(\mem<2><10> ), .B(n269), .Y(n1307) );
  INVX1 U897 ( .A(n1307), .Y(n1308) );
  AND2X2 U898 ( .A(\mem<2><11> ), .B(n269), .Y(n1309) );
  INVX1 U899 ( .A(n1309), .Y(n1310) );
  AND2X2 U900 ( .A(\mem<2><12> ), .B(n269), .Y(n1311) );
  INVX1 U901 ( .A(n1311), .Y(n1312) );
  AND2X2 U902 ( .A(\mem<2><13> ), .B(n269), .Y(n1313) );
  INVX1 U903 ( .A(n1313), .Y(n1314) );
  AND2X2 U904 ( .A(\mem<2><14> ), .B(n269), .Y(n1315) );
  INVX1 U905 ( .A(n1315), .Y(n1316) );
  AND2X2 U906 ( .A(\mem<1><0> ), .B(n271), .Y(n1317) );
  INVX1 U907 ( .A(n1317), .Y(n1318) );
  AND2X2 U908 ( .A(\mem<1><1> ), .B(n271), .Y(n1319) );
  INVX1 U909 ( .A(n1319), .Y(n1320) );
  AND2X2 U910 ( .A(\mem<1><2> ), .B(n271), .Y(n1321) );
  INVX1 U911 ( .A(n1321), .Y(n1322) );
  AND2X2 U912 ( .A(\mem<1><3> ), .B(n271), .Y(n1323) );
  INVX1 U913 ( .A(n1323), .Y(n1324) );
  AND2X2 U914 ( .A(\mem<1><4> ), .B(n271), .Y(n1325) );
  INVX1 U915 ( .A(n1325), .Y(n1326) );
  AND2X2 U916 ( .A(\mem<1><5> ), .B(n271), .Y(n1327) );
  INVX1 U917 ( .A(n1327), .Y(n1328) );
  AND2X2 U918 ( .A(\mem<1><6> ), .B(n271), .Y(n1329) );
  INVX1 U919 ( .A(n1329), .Y(n1330) );
  AND2X2 U920 ( .A(\mem<1><8> ), .B(n271), .Y(n1331) );
  INVX1 U921 ( .A(n1331), .Y(n1332) );
  AND2X2 U922 ( .A(\mem<1><9> ), .B(n271), .Y(n1333) );
  INVX1 U923 ( .A(n1333), .Y(n1334) );
  AND2X2 U924 ( .A(\mem<1><10> ), .B(n271), .Y(n1335) );
  INVX1 U925 ( .A(n1335), .Y(n1336) );
  AND2X2 U926 ( .A(\mem<1><11> ), .B(n271), .Y(n1337) );
  INVX1 U927 ( .A(n1337), .Y(n1338) );
  AND2X2 U928 ( .A(\mem<1><12> ), .B(n271), .Y(n1339) );
  INVX1 U929 ( .A(n1339), .Y(n1340) );
  AND2X2 U930 ( .A(\mem<1><13> ), .B(n271), .Y(n1341) );
  INVX1 U931 ( .A(n1341), .Y(n1342) );
  AND2X2 U932 ( .A(\mem<1><14> ), .B(n271), .Y(n1343) );
  INVX1 U933 ( .A(n1343), .Y(n1344) );
  AND2X2 U934 ( .A(\mem<0><0> ), .B(n206), .Y(n1345) );
  INVX1 U935 ( .A(n1345), .Y(n1346) );
  AND2X2 U936 ( .A(\mem<0><1> ), .B(n206), .Y(n1347) );
  INVX1 U937 ( .A(n1347), .Y(n1348) );
  AND2X2 U938 ( .A(\mem<0><2> ), .B(n206), .Y(n1349) );
  INVX1 U939 ( .A(n1349), .Y(n1350) );
  AND2X2 U940 ( .A(\mem<0><3> ), .B(n206), .Y(n1351) );
  INVX1 U941 ( .A(n1351), .Y(n1352) );
  AND2X2 U942 ( .A(\mem<0><4> ), .B(n206), .Y(n1353) );
  INVX1 U943 ( .A(n1353), .Y(n1354) );
  AND2X2 U944 ( .A(\mem<0><5> ), .B(n206), .Y(n1355) );
  INVX1 U945 ( .A(n1355), .Y(n1356) );
  AND2X2 U946 ( .A(\mem<0><6> ), .B(n206), .Y(n1357) );
  INVX1 U947 ( .A(n1357), .Y(n1358) );
  AND2X2 U948 ( .A(\mem<0><8> ), .B(n206), .Y(n1359) );
  INVX1 U949 ( .A(n1359), .Y(n1360) );
  AND2X2 U950 ( .A(\mem<0><9> ), .B(n206), .Y(n1361) );
  INVX1 U951 ( .A(n1361), .Y(n1362) );
  AND2X2 U952 ( .A(\mem<0><10> ), .B(n206), .Y(n1363) );
  INVX1 U953 ( .A(n1363), .Y(n1364) );
  AND2X2 U954 ( .A(\mem<0><11> ), .B(n206), .Y(n1365) );
  INVX1 U955 ( .A(n1365), .Y(n1366) );
  AND2X2 U956 ( .A(\mem<0><12> ), .B(n206), .Y(n1367) );
  INVX1 U957 ( .A(n1367), .Y(n1368) );
  AND2X2 U958 ( .A(\mem<0><13> ), .B(n206), .Y(n1369) );
  INVX1 U959 ( .A(n1369), .Y(n1370) );
  AND2X2 U960 ( .A(\mem<0><14> ), .B(n206), .Y(n1371) );
  INVX1 U961 ( .A(n1371), .Y(n1372) );
  BUFX2 U962 ( .A(n2137), .Y(n1373) );
  INVX1 U963 ( .A(n1373), .Y(n2248) );
  BUFX2 U964 ( .A(n2147), .Y(n1374) );
  INVX1 U965 ( .A(n1374), .Y(n2250) );
  BUFX2 U966 ( .A(n2157), .Y(n1375) );
  INVX1 U967 ( .A(n1375), .Y(n2251) );
  BUFX2 U968 ( .A(n2167), .Y(n1376) );
  INVX1 U969 ( .A(n1376), .Y(n2253) );
  BUFX2 U970 ( .A(n2177), .Y(n1377) );
  INVX1 U971 ( .A(n1377), .Y(n2255) );
  BUFX2 U972 ( .A(n2236), .Y(n1378) );
  INVX1 U973 ( .A(n1378), .Y(n2244) );
  BUFX2 U974 ( .A(n2245), .Y(n1379) );
  INVX1 U975 ( .A(n1379), .Y(n2257) );
  AND2X1 U976 ( .A(n2108), .B(n295), .Y(n1380) );
  AND2X1 U977 ( .A(n2114), .B(n296), .Y(n1381) );
  AND2X1 U978 ( .A(n2109), .B(n295), .Y(n1382) );
  AND2X1 U979 ( .A(n2115), .B(n296), .Y(n1383) );
  AND2X1 U980 ( .A(n1381), .B(n2258), .Y(n1384) );
  AND2X1 U981 ( .A(n2258), .B(n1383), .Y(n1385) );
  AND2X1 U982 ( .A(n2258), .B(n2244), .Y(n1386) );
  AND2X1 U983 ( .A(n2258), .B(n2257), .Y(n1387) );
  AND2X1 U984 ( .A(n1380), .B(n1381), .Y(n1388) );
  INVX1 U985 ( .A(n1388), .Y(n1389) );
  AND2X1 U986 ( .A(n1381), .B(n1382), .Y(n1390) );
  INVX1 U987 ( .A(n1390), .Y(n1391) );
  AND2X1 U988 ( .A(n1381), .B(n2248), .Y(n1392) );
  INVX1 U989 ( .A(n1392), .Y(n1393) );
  AND2X1 U990 ( .A(n1381), .B(n2250), .Y(n1394) );
  INVX1 U991 ( .A(n1394), .Y(n1395) );
  AND2X1 U992 ( .A(n1381), .B(n2251), .Y(n1396) );
  INVX1 U993 ( .A(n1396), .Y(n1397) );
  AND2X1 U994 ( .A(n1381), .B(n2253), .Y(n1398) );
  INVX1 U995 ( .A(n1398), .Y(n1399) );
  AND2X1 U996 ( .A(n1381), .B(n2255), .Y(n1400) );
  INVX1 U997 ( .A(n1400), .Y(n1401) );
  AND2X1 U998 ( .A(n1380), .B(n1383), .Y(n1402) );
  INVX1 U999 ( .A(n1402), .Y(n1403) );
  AND2X1 U1000 ( .A(n1382), .B(n1383), .Y(n1404) );
  INVX1 U1001 ( .A(n1404), .Y(n1405) );
  AND2X1 U1002 ( .A(n2248), .B(n1383), .Y(n1406) );
  INVX1 U1003 ( .A(n1406), .Y(n1407) );
  AND2X1 U1004 ( .A(n2250), .B(n1383), .Y(n1408) );
  INVX1 U1005 ( .A(n1408), .Y(n1409) );
  AND2X1 U1006 ( .A(n2251), .B(n1383), .Y(n1410) );
  INVX1 U1007 ( .A(n1410), .Y(n1411) );
  BUFX2 U1008 ( .A(n184), .Y(n2038) );
  AND2X1 U1009 ( .A(n2253), .B(n1383), .Y(n1412) );
  INVX1 U1010 ( .A(n1412), .Y(n1413) );
  AND2X1 U1011 ( .A(n2255), .B(n1383), .Y(n1414) );
  INVX1 U1012 ( .A(n1414), .Y(n1415) );
  AND2X1 U1013 ( .A(n1380), .B(n2244), .Y(n1416) );
  INVX1 U1014 ( .A(n1416), .Y(n1417) );
  AND2X1 U1015 ( .A(n1382), .B(n2244), .Y(n1418) );
  INVX1 U1016 ( .A(n1418), .Y(n1419) );
  AND2X1 U1017 ( .A(n2248), .B(n2244), .Y(n1420) );
  INVX1 U1018 ( .A(n1420), .Y(n1421) );
  AND2X1 U1019 ( .A(n2250), .B(n2244), .Y(n1422) );
  INVX1 U1020 ( .A(n1422), .Y(n1423) );
  AND2X1 U1021 ( .A(n2251), .B(n2244), .Y(n1424) );
  INVX1 U1022 ( .A(n1424), .Y(n1425) );
  AND2X1 U1023 ( .A(n2253), .B(n2244), .Y(n1426) );
  INVX1 U1024 ( .A(n1426), .Y(n1427) );
  AND2X1 U1025 ( .A(n2255), .B(n2244), .Y(n1428) );
  INVX1 U1026 ( .A(n1428), .Y(n1429) );
  AND2X1 U1027 ( .A(n1380), .B(n2257), .Y(n1430) );
  INVX1 U1028 ( .A(n1430), .Y(n1431) );
  AND2X1 U1029 ( .A(n1382), .B(n2257), .Y(n1432) );
  INVX1 U1030 ( .A(n1432), .Y(n1433) );
  AND2X1 U1031 ( .A(n2248), .B(n2257), .Y(n1434) );
  INVX1 U1032 ( .A(n1434), .Y(n1435) );
  AND2X1 U1033 ( .A(n2250), .B(n2257), .Y(n1436) );
  INVX1 U1034 ( .A(n1436), .Y(n1437) );
  AND2X1 U1035 ( .A(n2251), .B(n2257), .Y(n1438) );
  INVX1 U1036 ( .A(n1438), .Y(n1439) );
  AND2X1 U1037 ( .A(n2253), .B(n2257), .Y(n1440) );
  INVX1 U1038 ( .A(n1440), .Y(n1441) );
  AND2X1 U1039 ( .A(n2255), .B(n2257), .Y(n1442) );
  INVX1 U1040 ( .A(n1442), .Y(n1443) );
  AND2X1 U1041 ( .A(N21), .B(n2107), .Y(n1444) );
  AND2X2 U1042 ( .A(n1469), .B(n2107), .Y(n1470) );
  INVX1 U1043 ( .A(rst), .Y(n2107) );
  INVX1 U1044 ( .A(n233), .Y(n1445) );
  INVX1 U1045 ( .A(n233), .Y(n1446) );
  INVX1 U1046 ( .A(n233), .Y(n1447) );
  INVX1 U1047 ( .A(n233), .Y(n1448) );
  INVX1 U1048 ( .A(n233), .Y(n1449) );
  INVX1 U1049 ( .A(n233), .Y(n1450) );
  INVX1 U1050 ( .A(n274), .Y(n1451) );
  INVX1 U1051 ( .A(n274), .Y(n1452) );
  INVX1 U1052 ( .A(n274), .Y(n1453) );
  INVX1 U1053 ( .A(n1456), .Y(n1454) );
  INVX1 U1054 ( .A(n273), .Y(n1455) );
  INVX1 U1055 ( .A(n272), .Y(n1456) );
  INVX1 U1056 ( .A(n1455), .Y(n1457) );
  INVX1 U1057 ( .A(n1455), .Y(n1458) );
  INVX1 U1058 ( .A(n1456), .Y(n1459) );
  INVX1 U1059 ( .A(n1456), .Y(n1460) );
  INVX1 U1060 ( .A(n273), .Y(n1461) );
  INVX1 U1061 ( .A(n1461), .Y(n1462) );
  INVX1 U1062 ( .A(n1461), .Y(n1463) );
  INVX1 U1063 ( .A(n276), .Y(n1464) );
  INVX1 U1064 ( .A(n274), .Y(n1465) );
  INVX1 U1065 ( .A(n274), .Y(n1466) );
  INVX1 U1066 ( .A(n1464), .Y(n1467) );
  INVX1 U1067 ( .A(n1464), .Y(n1468) );
  INVX1 U1068 ( .A(n2107), .Y(n2106) );
  INVX1 U1069 ( .A(n2117), .Y(n2118) );
  INVX1 U1070 ( .A(n2117), .Y(n1471) );
  INVX1 U1071 ( .A(n2117), .Y(n1472) );
  INVX1 U1072 ( .A(N12), .Y(n2113) );
  MUX2X1 U1073 ( .B(n1474), .A(n1475), .S(n1978), .Y(n1473) );
  MUX2X1 U1074 ( .B(n1477), .A(n1478), .S(n1983), .Y(n1476) );
  MUX2X1 U1075 ( .B(n1480), .A(n1481), .S(n1977), .Y(n1479) );
  MUX2X1 U1076 ( .B(n1483), .A(n1484), .S(n1977), .Y(n1482) );
  MUX2X1 U1077 ( .B(n1486), .A(n1487), .S(n1972), .Y(n1485) );
  MUX2X1 U1078 ( .B(n1489), .A(n1490), .S(n1978), .Y(n1488) );
  MUX2X1 U1079 ( .B(n1492), .A(n1493), .S(n1978), .Y(n1491) );
  MUX2X1 U1080 ( .B(n1495), .A(n1496), .S(n1983), .Y(n1494) );
  MUX2X1 U1081 ( .B(n1498), .A(n1499), .S(n1977), .Y(n1497) );
  MUX2X1 U1082 ( .B(n1501), .A(n1502), .S(n1972), .Y(n1500) );
  MUX2X1 U1083 ( .B(n1504), .A(n1505), .S(n1977), .Y(n1503) );
  MUX2X1 U1084 ( .B(n1507), .A(n1508), .S(n1977), .Y(n1506) );
  MUX2X1 U1085 ( .B(n1510), .A(n1511), .S(n1977), .Y(n1509) );
  MUX2X1 U1086 ( .B(n1513), .A(n1514), .S(n1977), .Y(n1512) );
  MUX2X1 U1087 ( .B(n1516), .A(n1517), .S(n1972), .Y(n1515) );
  MUX2X1 U1088 ( .B(n1519), .A(n1520), .S(n1977), .Y(n1518) );
  MUX2X1 U1089 ( .B(n1522), .A(n1523), .S(n1977), .Y(n1521) );
  MUX2X1 U1090 ( .B(n1525), .A(n1526), .S(n1977), .Y(n1524) );
  MUX2X1 U1091 ( .B(n1528), .A(n1529), .S(n1977), .Y(n1527) );
  MUX2X1 U1092 ( .B(n1531), .A(n1532), .S(n1972), .Y(n1530) );
  MUX2X1 U1093 ( .B(n1534), .A(n1535), .S(n1977), .Y(n1533) );
  MUX2X1 U1094 ( .B(n1537), .A(n1538), .S(n1977), .Y(n1536) );
  MUX2X1 U1095 ( .B(n1540), .A(n1541), .S(n1977), .Y(n1539) );
  MUX2X1 U1096 ( .B(n1543), .A(n1544), .S(n1977), .Y(n1542) );
  MUX2X1 U1097 ( .B(n1546), .A(n1547), .S(n1972), .Y(n1545) );
  MUX2X1 U1098 ( .B(n1549), .A(n1550), .S(n1978), .Y(n1548) );
  MUX2X1 U1099 ( .B(n1552), .A(n1553), .S(n1978), .Y(n1551) );
  MUX2X1 U1100 ( .B(n1555), .A(n1556), .S(n1978), .Y(n1554) );
  MUX2X1 U1101 ( .B(n1558), .A(n1559), .S(n1978), .Y(n1557) );
  MUX2X1 U1102 ( .B(n1561), .A(n1562), .S(n1972), .Y(n1560) );
  MUX2X1 U1103 ( .B(n1564), .A(n1565), .S(n1978), .Y(n1563) );
  MUX2X1 U1104 ( .B(n1567), .A(n1568), .S(n1978), .Y(n1566) );
  MUX2X1 U1105 ( .B(n1570), .A(n1571), .S(n1978), .Y(n1569) );
  MUX2X1 U1106 ( .B(n1573), .A(n1574), .S(n1978), .Y(n1572) );
  MUX2X1 U1107 ( .B(n1576), .A(n1577), .S(n1972), .Y(n1575) );
  MUX2X1 U1108 ( .B(n1579), .A(n1580), .S(n1978), .Y(n1578) );
  MUX2X1 U1109 ( .B(n1582), .A(n1583), .S(n1978), .Y(n1581) );
  MUX2X1 U1110 ( .B(n1585), .A(n1586), .S(n1978), .Y(n1584) );
  MUX2X1 U1111 ( .B(n1588), .A(n1589), .S(n1978), .Y(n1587) );
  MUX2X1 U1112 ( .B(n1591), .A(n1592), .S(n1972), .Y(n1590) );
  MUX2X1 U1113 ( .B(n1594), .A(n1595), .S(n1979), .Y(n1593) );
  MUX2X1 U1114 ( .B(n1597), .A(n1598), .S(n1979), .Y(n1596) );
  MUX2X1 U1115 ( .B(n1600), .A(n1601), .S(n1979), .Y(n1599) );
  MUX2X1 U1116 ( .B(n1603), .A(n1604), .S(n1979), .Y(n1602) );
  MUX2X1 U1117 ( .B(n1606), .A(n1607), .S(n1972), .Y(n1605) );
  MUX2X1 U1118 ( .B(n1609), .A(n1610), .S(n1979), .Y(n1608) );
  MUX2X1 U1119 ( .B(n1612), .A(n1613), .S(n1979), .Y(n1611) );
  MUX2X1 U1120 ( .B(n1615), .A(n1616), .S(n1979), .Y(n1614) );
  MUX2X1 U1121 ( .B(n1618), .A(n1619), .S(n1979), .Y(n1617) );
  MUX2X1 U1122 ( .B(n1621), .A(n1622), .S(n1972), .Y(n1620) );
  MUX2X1 U1123 ( .B(n1624), .A(n1625), .S(n1979), .Y(n1623) );
  MUX2X1 U1124 ( .B(n1627), .A(n1628), .S(n1979), .Y(n1626) );
  MUX2X1 U1125 ( .B(n1630), .A(n1631), .S(n1979), .Y(n1629) );
  MUX2X1 U1126 ( .B(n1633), .A(n1634), .S(n1979), .Y(n1632) );
  MUX2X1 U1127 ( .B(n1636), .A(n1637), .S(n1972), .Y(n1635) );
  MUX2X1 U1128 ( .B(n1639), .A(n1640), .S(n1980), .Y(n1638) );
  MUX2X1 U1129 ( .B(n1642), .A(n1643), .S(n1980), .Y(n1641) );
  MUX2X1 U1130 ( .B(n1645), .A(n1646), .S(n1980), .Y(n1644) );
  MUX2X1 U1131 ( .B(n1648), .A(n1649), .S(n1980), .Y(n1647) );
  MUX2X1 U1132 ( .B(n1651), .A(n1652), .S(n1972), .Y(n1650) );
  MUX2X1 U1133 ( .B(n1654), .A(n1655), .S(n1980), .Y(n1653) );
  MUX2X1 U1134 ( .B(n1657), .A(n1658), .S(n1980), .Y(n1656) );
  MUX2X1 U1135 ( .B(n1660), .A(n1661), .S(n1980), .Y(n1659) );
  MUX2X1 U1136 ( .B(n1663), .A(n1664), .S(n1980), .Y(n1662) );
  MUX2X1 U1137 ( .B(n1666), .A(n1667), .S(n1971), .Y(n1665) );
  MUX2X1 U1138 ( .B(n1669), .A(n1670), .S(n1980), .Y(n1668) );
  MUX2X1 U1139 ( .B(n1672), .A(n1673), .S(n1980), .Y(n1671) );
  MUX2X1 U1140 ( .B(n1675), .A(n1676), .S(n1980), .Y(n1674) );
  MUX2X1 U1141 ( .B(n1678), .A(n1679), .S(n1980), .Y(n1677) );
  MUX2X1 U1142 ( .B(n1681), .A(n1682), .S(n1971), .Y(n1680) );
  MUX2X1 U1143 ( .B(n1684), .A(n1685), .S(n1981), .Y(n1683) );
  MUX2X1 U1144 ( .B(n1687), .A(n1688), .S(n1981), .Y(n1686) );
  MUX2X1 U1145 ( .B(n1690), .A(n1691), .S(n1981), .Y(n1689) );
  MUX2X1 U1146 ( .B(n1693), .A(n1694), .S(n1981), .Y(n1692) );
  MUX2X1 U1147 ( .B(n1696), .A(n1697), .S(n1971), .Y(n1695) );
  MUX2X1 U1148 ( .B(n1699), .A(n1700), .S(n1981), .Y(n1698) );
  MUX2X1 U1149 ( .B(n1702), .A(n1703), .S(n1981), .Y(n1701) );
  MUX2X1 U1150 ( .B(n1705), .A(n1706), .S(n1981), .Y(n1704) );
  MUX2X1 U1151 ( .B(n1708), .A(n1709), .S(n1981), .Y(n1707) );
  MUX2X1 U1152 ( .B(n1711), .A(n1712), .S(n1971), .Y(n1710) );
  MUX2X1 U1153 ( .B(n1714), .A(n1715), .S(n1981), .Y(n1713) );
  MUX2X1 U1154 ( .B(n1717), .A(n1718), .S(n1981), .Y(n1716) );
  MUX2X1 U1155 ( .B(n1720), .A(n1721), .S(n1981), .Y(n1719) );
  MUX2X1 U1156 ( .B(n1723), .A(n1724), .S(n1981), .Y(n1722) );
  MUX2X1 U1157 ( .B(n1726), .A(n1727), .S(n1971), .Y(n1725) );
  MUX2X1 U1158 ( .B(n1729), .A(n1730), .S(n1982), .Y(n1728) );
  MUX2X1 U1159 ( .B(n1732), .A(n1733), .S(n1982), .Y(n1731) );
  MUX2X1 U1160 ( .B(n1735), .A(n1736), .S(n1982), .Y(n1734) );
  MUX2X1 U1161 ( .B(n1738), .A(n1739), .S(n1982), .Y(n1737) );
  MUX2X1 U1162 ( .B(n1741), .A(n1742), .S(n1971), .Y(n1740) );
  MUX2X1 U1163 ( .B(n1744), .A(n1745), .S(n1982), .Y(n1743) );
  MUX2X1 U1164 ( .B(n1747), .A(n1748), .S(n1982), .Y(n1746) );
  MUX2X1 U1165 ( .B(n1750), .A(n1751), .S(n1982), .Y(n1749) );
  MUX2X1 U1166 ( .B(n1753), .A(n1754), .S(n1982), .Y(n1752) );
  MUX2X1 U1167 ( .B(n1756), .A(n1757), .S(n1971), .Y(n1755) );
  MUX2X1 U1168 ( .B(n1759), .A(n1760), .S(n1982), .Y(n1758) );
  MUX2X1 U1169 ( .B(n1762), .A(n1763), .S(n1982), .Y(n1761) );
  MUX2X1 U1170 ( .B(n1765), .A(n1766), .S(n1982), .Y(n1764) );
  MUX2X1 U1171 ( .B(n1768), .A(n1769), .S(n1982), .Y(n1767) );
  MUX2X1 U1172 ( .B(n1771), .A(n1772), .S(n1971), .Y(n1770) );
  MUX2X1 U1173 ( .B(n1774), .A(n1775), .S(n1982), .Y(n1773) );
  MUX2X1 U1174 ( .B(n1777), .A(n1778), .S(n1982), .Y(n1776) );
  MUX2X1 U1175 ( .B(n1780), .A(n1781), .S(n1982), .Y(n1779) );
  MUX2X1 U1177 ( .B(n1783), .A(n1784), .S(n1982), .Y(n1782) );
  MUX2X1 U1178 ( .B(n1786), .A(n1787), .S(n1971), .Y(n1785) );
  MUX2X1 U1179 ( .B(n1789), .A(n1790), .S(n1982), .Y(n1788) );
  MUX2X1 U1180 ( .B(n1792), .A(n1793), .S(n1982), .Y(n1791) );
  MUX2X1 U1181 ( .B(n1795), .A(n1796), .S(n1982), .Y(n1794) );
  MUX2X1 U1182 ( .B(n1798), .A(n1799), .S(n1982), .Y(n1797) );
  MUX2X1 U1183 ( .B(n1801), .A(n1802), .S(n1971), .Y(n1800) );
  MUX2X1 U1184 ( .B(n1804), .A(n1805), .S(n1982), .Y(n1803) );
  MUX2X1 U1185 ( .B(n1807), .A(n1808), .S(n1982), .Y(n1806) );
  MUX2X1 U1186 ( .B(n1810), .A(n1811), .S(n1982), .Y(n1809) );
  MUX2X1 U1187 ( .B(n1813), .A(n1814), .S(n1982), .Y(n1812) );
  MUX2X1 U1188 ( .B(n1816), .A(n1817), .S(n1971), .Y(n1815) );
  MUX2X1 U1189 ( .B(n1819), .A(n1820), .S(n1982), .Y(n1818) );
  MUX2X1 U1190 ( .B(n1822), .A(n1823), .S(n1982), .Y(n1821) );
  MUX2X1 U1191 ( .B(n1825), .A(n1826), .S(n1982), .Y(n1824) );
  MUX2X1 U1192 ( .B(n1828), .A(n1829), .S(n1982), .Y(n1827) );
  MUX2X1 U1193 ( .B(n1831), .A(n1832), .S(n1971), .Y(n1830) );
  MUX2X1 U1194 ( .B(n1834), .A(n1835), .S(n1982), .Y(n1833) );
  MUX2X1 U1195 ( .B(n1837), .A(n1838), .S(n1982), .Y(n1836) );
  MUX2X1 U1196 ( .B(n1840), .A(n1841), .S(n1982), .Y(n1839) );
  MUX2X1 U1197 ( .B(n1843), .A(n1844), .S(n1982), .Y(n1842) );
  MUX2X1 U1198 ( .B(n1846), .A(n1847), .S(n1970), .Y(n1845) );
  MUX2X1 U1199 ( .B(n1849), .A(n1850), .S(n1982), .Y(n1848) );
  MUX2X1 U1200 ( .B(n1852), .A(n1853), .S(n1982), .Y(n1851) );
  MUX2X1 U1201 ( .B(n1855), .A(n1856), .S(n1982), .Y(n1854) );
  MUX2X1 U1202 ( .B(n1858), .A(n1859), .S(n1982), .Y(n1857) );
  MUX2X1 U1203 ( .B(n1861), .A(n1862), .S(n1970), .Y(n1860) );
  MUX2X1 U1204 ( .B(n1864), .A(n1865), .S(n1983), .Y(n1863) );
  MUX2X1 U1205 ( .B(n1867), .A(n1868), .S(n1983), .Y(n1866) );
  MUX2X1 U1206 ( .B(n1870), .A(n1871), .S(n1983), .Y(n1869) );
  MUX2X1 U1207 ( .B(n1873), .A(n1874), .S(n1983), .Y(n1872) );
  MUX2X1 U1208 ( .B(n1876), .A(n1877), .S(n1970), .Y(n1875) );
  MUX2X1 U1209 ( .B(n1879), .A(n1880), .S(n1983), .Y(n1878) );
  MUX2X1 U1210 ( .B(n1882), .A(n1883), .S(n1983), .Y(n1881) );
  MUX2X1 U1211 ( .B(n1885), .A(n1886), .S(n1983), .Y(n1884) );
  MUX2X1 U1212 ( .B(n1888), .A(n1889), .S(n1983), .Y(n1887) );
  MUX2X1 U1213 ( .B(n1891), .A(n1892), .S(n1970), .Y(n1890) );
  MUX2X1 U1214 ( .B(n1894), .A(n1895), .S(n1983), .Y(n1893) );
  MUX2X1 U1215 ( .B(n1897), .A(n1898), .S(n1983), .Y(n1896) );
  MUX2X1 U1216 ( .B(n1900), .A(n1901), .S(n1983), .Y(n1899) );
  MUX2X1 U1217 ( .B(n1903), .A(n1904), .S(n1983), .Y(n1902) );
  MUX2X1 U1218 ( .B(n1906), .A(n1907), .S(n1970), .Y(n1905) );
  MUX2X1 U1219 ( .B(n1909), .A(n1910), .S(n1981), .Y(n1908) );
  MUX2X1 U1220 ( .B(n1912), .A(n1913), .S(n1979), .Y(n1911) );
  MUX2X1 U1221 ( .B(n1915), .A(n1916), .S(n1980), .Y(n1914) );
  MUX2X1 U1222 ( .B(n1918), .A(n1919), .S(n1981), .Y(n1917) );
  MUX2X1 U1223 ( .B(n1921), .A(n1922), .S(n1970), .Y(n1920) );
  MUX2X1 U1224 ( .B(n1924), .A(n1925), .S(n1981), .Y(n1923) );
  MUX2X1 U1225 ( .B(n1927), .A(n1928), .S(n1981), .Y(n1926) );
  MUX2X1 U1226 ( .B(n1930), .A(n1931), .S(n1979), .Y(n1929) );
  MUX2X1 U1227 ( .B(n1933), .A(n1934), .S(n1979), .Y(n1932) );
  MUX2X1 U1228 ( .B(n1936), .A(n1937), .S(n1970), .Y(n1935) );
  MUX2X1 U1229 ( .B(n1939), .A(n1940), .S(n1980), .Y(n1938) );
  MUX2X1 U1230 ( .B(n1942), .A(n1943), .S(n1981), .Y(n1941) );
  MUX2X1 U1231 ( .B(n1945), .A(n1946), .S(n1980), .Y(n1944) );
  MUX2X1 U1232 ( .B(n1948), .A(n1949), .S(n1979), .Y(n1947) );
  MUX2X1 U1233 ( .B(n1951), .A(n1952), .S(n1970), .Y(n1950) );
  MUX2X1 U1234 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1988), .Y(n1475) );
  MUX2X1 U1235 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1988), .Y(n1474) );
  MUX2X1 U1236 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1988), .Y(n1478) );
  MUX2X1 U1237 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1988), .Y(n1477) );
  MUX2X1 U1238 ( .B(n1476), .A(n1473), .S(n1974), .Y(n1487) );
  MUX2X1 U1239 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1989), .Y(n1481) );
  MUX2X1 U1240 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1989), .Y(n1480) );
  MUX2X1 U1241 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1989), .Y(n1484) );
  MUX2X1 U1242 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1989), .Y(n1483) );
  MUX2X1 U1243 ( .B(n1482), .A(n1479), .S(n1974), .Y(n1486) );
  MUX2X1 U1244 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1989), .Y(n1490) );
  MUX2X1 U1245 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1989), .Y(n1489) );
  MUX2X1 U1246 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1989), .Y(n1493) );
  MUX2X1 U1247 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1989), .Y(n1492) );
  MUX2X1 U1248 ( .B(n1491), .A(n1488), .S(n1974), .Y(n1502) );
  MUX2X1 U1249 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1989), .Y(n1496) );
  MUX2X1 U1250 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1989), .Y(n1495) );
  MUX2X1 U1251 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1989), .Y(n1499) );
  MUX2X1 U1252 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1989), .Y(n1498) );
  MUX2X1 U1253 ( .B(n1497), .A(n1494), .S(n1974), .Y(n1501) );
  MUX2X1 U1254 ( .B(n1500), .A(n1485), .S(n1969), .Y(n1953) );
  MUX2X1 U1255 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1990), .Y(n1505) );
  MUX2X1 U1256 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1990), .Y(n1504) );
  MUX2X1 U1257 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1990), .Y(n1508) );
  MUX2X1 U1258 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1990), .Y(n1507) );
  MUX2X1 U1259 ( .B(n1506), .A(n1503), .S(n1974), .Y(n1517) );
  MUX2X1 U1260 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1990), .Y(n1511) );
  MUX2X1 U1261 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1990), .Y(n1510) );
  MUX2X1 U1262 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1990), .Y(n1514) );
  MUX2X1 U1263 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1990), .Y(n1513) );
  MUX2X1 U1264 ( .B(n1512), .A(n1509), .S(n1974), .Y(n1516) );
  MUX2X1 U1265 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1990), .Y(n1520) );
  MUX2X1 U1266 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1990), .Y(n1519) );
  MUX2X1 U1267 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1990), .Y(n1523) );
  MUX2X1 U1268 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1990), .Y(n1522) );
  MUX2X1 U1269 ( .B(n1521), .A(n1518), .S(n1974), .Y(n1532) );
  MUX2X1 U1270 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1991), .Y(n1526) );
  MUX2X1 U1271 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1991), .Y(n1525) );
  MUX2X1 U1272 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1991), .Y(n1529) );
  MUX2X1 U1273 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1991), .Y(n1528) );
  MUX2X1 U1274 ( .B(n1527), .A(n1524), .S(n1974), .Y(n1531) );
  MUX2X1 U1275 ( .B(n1530), .A(n1515), .S(n1969), .Y(n1954) );
  MUX2X1 U1276 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1991), .Y(n1535) );
  MUX2X1 U1277 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1991), .Y(n1534) );
  MUX2X1 U1278 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1991), .Y(n1538) );
  MUX2X1 U1279 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1991), .Y(n1537) );
  MUX2X1 U1280 ( .B(n1536), .A(n1533), .S(n1974), .Y(n1547) );
  MUX2X1 U1281 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1991), .Y(n1541) );
  MUX2X1 U1282 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1991), .Y(n1540) );
  MUX2X1 U1283 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1991), .Y(n1544) );
  MUX2X1 U1284 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1991), .Y(n1543) );
  MUX2X1 U1285 ( .B(n1542), .A(n1539), .S(n1974), .Y(n1546) );
  MUX2X1 U1286 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1992), .Y(n1550) );
  MUX2X1 U1287 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1992), .Y(n1549) );
  MUX2X1 U1288 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1992), .Y(n1553) );
  MUX2X1 U1289 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1992), .Y(n1552) );
  MUX2X1 U1290 ( .B(n1551), .A(n1548), .S(n1974), .Y(n1562) );
  MUX2X1 U1291 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1992), .Y(n1556) );
  MUX2X1 U1292 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1992), .Y(n1555) );
  MUX2X1 U1293 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1992), .Y(n1559) );
  MUX2X1 U1294 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1992), .Y(n1558) );
  MUX2X1 U1295 ( .B(n1557), .A(n1554), .S(n1974), .Y(n1561) );
  MUX2X1 U1296 ( .B(n1560), .A(n1545), .S(n1969), .Y(n1955) );
  MUX2X1 U1297 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1992), .Y(n1565) );
  MUX2X1 U1298 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1992), .Y(n1564) );
  MUX2X1 U1299 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1992), .Y(n1568) );
  MUX2X1 U1300 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1992), .Y(n1567) );
  MUX2X1 U1301 ( .B(n1566), .A(n1563), .S(n1974), .Y(n1577) );
  MUX2X1 U1302 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1993), .Y(n1571) );
  MUX2X1 U1303 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1993), .Y(n1570) );
  MUX2X1 U1304 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1993), .Y(n1574) );
  MUX2X1 U1305 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1993), .Y(n1573) );
  MUX2X1 U1306 ( .B(n1572), .A(n1569), .S(n1974), .Y(n1576) );
  MUX2X1 U1307 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1993), .Y(n1580) );
  MUX2X1 U1308 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1993), .Y(n1579) );
  MUX2X1 U1309 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1993), .Y(n1583) );
  MUX2X1 U1310 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1993), .Y(n1582) );
  MUX2X1 U1311 ( .B(n1581), .A(n1578), .S(n2112), .Y(n1592) );
  MUX2X1 U1312 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1993), .Y(n1586) );
  MUX2X1 U1313 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1993), .Y(n1585) );
  MUX2X1 U1314 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1993), .Y(n1589) );
  MUX2X1 U1315 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1993), .Y(n1588) );
  MUX2X1 U1316 ( .B(n1587), .A(n1584), .S(n2112), .Y(n1591) );
  MUX2X1 U1317 ( .B(n1590), .A(n1575), .S(n1969), .Y(n1956) );
  MUX2X1 U1318 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1994), .Y(n1595) );
  MUX2X1 U1319 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1994), .Y(n1594) );
  MUX2X1 U1320 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1994), .Y(n1598) );
  MUX2X1 U1321 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1994), .Y(n1597) );
  MUX2X1 U1322 ( .B(n1596), .A(n1593), .S(n2112), .Y(n1607) );
  MUX2X1 U1323 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1994), .Y(n1601) );
  MUX2X1 U1324 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1994), .Y(n1600) );
  MUX2X1 U1325 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1994), .Y(n1604) );
  MUX2X1 U1326 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1994), .Y(n1603) );
  MUX2X1 U1327 ( .B(n1602), .A(n1599), .S(n2112), .Y(n1606) );
  MUX2X1 U1328 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1994), .Y(n1610) );
  MUX2X1 U1329 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1994), .Y(n1609) );
  MUX2X1 U1330 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1994), .Y(n1613) );
  MUX2X1 U1331 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1994), .Y(n1612) );
  MUX2X1 U1332 ( .B(n1611), .A(n1608), .S(n2112), .Y(n1622) );
  MUX2X1 U1333 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1995), .Y(n1616) );
  MUX2X1 U1334 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1995), .Y(n1615) );
  MUX2X1 U1335 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1995), .Y(n1619) );
  MUX2X1 U1336 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1995), .Y(n1618) );
  MUX2X1 U1337 ( .B(n1617), .A(n1614), .S(n2112), .Y(n1621) );
  MUX2X1 U1338 ( .B(n1620), .A(n1605), .S(n1969), .Y(n1957) );
  MUX2X1 U1339 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1995), .Y(n1625) );
  MUX2X1 U1340 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1995), .Y(n1624) );
  MUX2X1 U1341 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1995), .Y(n1628) );
  MUX2X1 U1342 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1995), .Y(n1627) );
  MUX2X1 U1343 ( .B(n1626), .A(n1623), .S(n2112), .Y(n1637) );
  MUX2X1 U1344 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1995), .Y(n1631) );
  MUX2X1 U1345 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1995), .Y(n1630) );
  MUX2X1 U1346 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1995), .Y(n1634) );
  MUX2X1 U1347 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1995), .Y(n1633) );
  MUX2X1 U1348 ( .B(n1632), .A(n1629), .S(n1974), .Y(n1636) );
  MUX2X1 U1349 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1996), .Y(n1640) );
  MUX2X1 U1350 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1996), .Y(n1639) );
  MUX2X1 U1351 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1996), .Y(n1643) );
  MUX2X1 U1352 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1996), .Y(n1642) );
  MUX2X1 U1353 ( .B(n1641), .A(n1638), .S(n2112), .Y(n1652) );
  MUX2X1 U1354 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1996), .Y(n1646) );
  MUX2X1 U1355 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1996), .Y(n1645) );
  MUX2X1 U1356 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1996), .Y(n1649) );
  MUX2X1 U1357 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1996), .Y(n1648) );
  MUX2X1 U1358 ( .B(n1647), .A(n1644), .S(n2112), .Y(n1651) );
  MUX2X1 U1359 ( .B(n1650), .A(n1635), .S(n1969), .Y(n1958) );
  MUX2X1 U1360 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1996), .Y(n1655) );
  MUX2X1 U1361 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1996), .Y(n1654) );
  MUX2X1 U1362 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1996), .Y(n1658) );
  MUX2X1 U1363 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1996), .Y(n1657) );
  MUX2X1 U1364 ( .B(n1656), .A(n1653), .S(n1974), .Y(n1667) );
  MUX2X1 U1365 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1997), .Y(n1661) );
  MUX2X1 U1366 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1997), .Y(n1660) );
  MUX2X1 U1367 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1997), .Y(n1664) );
  MUX2X1 U1368 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1997), .Y(n1663) );
  MUX2X1 U1369 ( .B(n1662), .A(n1659), .S(n1974), .Y(n1666) );
  MUX2X1 U1370 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1997), .Y(n1670) );
  MUX2X1 U1371 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1997), .Y(n1669) );
  MUX2X1 U1372 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1997), .Y(n1673) );
  MUX2X1 U1373 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1997), .Y(n1672) );
  MUX2X1 U1374 ( .B(n1671), .A(n1668), .S(n1974), .Y(n1682) );
  MUX2X1 U1375 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1997), .Y(n1676) );
  MUX2X1 U1376 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1997), .Y(n1675) );
  MUX2X1 U1377 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1997), .Y(n1679) );
  MUX2X1 U1378 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1997), .Y(n1678) );
  MUX2X1 U1379 ( .B(n1677), .A(n1674), .S(n1974), .Y(n1681) );
  MUX2X1 U1380 ( .B(n1680), .A(n1665), .S(n1969), .Y(n1959) );
  MUX2X1 U1381 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1998), .Y(n1685) );
  MUX2X1 U1382 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1998), .Y(n1684) );
  MUX2X1 U1383 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1998), .Y(n1688) );
  MUX2X1 U1384 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1998), .Y(n1687) );
  MUX2X1 U1385 ( .B(n1686), .A(n1683), .S(n1974), .Y(n1697) );
  MUX2X1 U1386 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1998), .Y(n1691) );
  MUX2X1 U1387 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1998), .Y(n1690) );
  MUX2X1 U1388 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1998), .Y(n1694) );
  MUX2X1 U1389 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1998), .Y(n1693) );
  MUX2X1 U1390 ( .B(n1692), .A(n1689), .S(n1974), .Y(n1696) );
  MUX2X1 U1391 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1998), .Y(n1700) );
  MUX2X1 U1392 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1998), .Y(n1699) );
  MUX2X1 U1393 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1998), .Y(n1703) );
  MUX2X1 U1394 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1998), .Y(n1702) );
  MUX2X1 U1395 ( .B(n1701), .A(n1698), .S(n1974), .Y(n1712) );
  MUX2X1 U1396 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1999), .Y(n1706) );
  MUX2X1 U1397 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1999), .Y(n1705) );
  MUX2X1 U1398 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1999), .Y(n1709) );
  MUX2X1 U1399 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1999), .Y(n1708) );
  MUX2X1 U1400 ( .B(n1707), .A(n1704), .S(n1974), .Y(n1711) );
  MUX2X1 U1401 ( .B(n1710), .A(n1695), .S(n1969), .Y(n1960) );
  MUX2X1 U1402 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1999), .Y(n1715) );
  MUX2X1 U1403 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1999), .Y(n1714) );
  MUX2X1 U1404 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1999), .Y(n1718) );
  MUX2X1 U1405 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1999), .Y(n1717) );
  MUX2X1 U1406 ( .B(n1716), .A(n1713), .S(n1974), .Y(n1727) );
  MUX2X1 U1407 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1999), .Y(n1721) );
  MUX2X1 U1408 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1999), .Y(n1720) );
  MUX2X1 U1409 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1999), .Y(n1724) );
  MUX2X1 U1410 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1999), .Y(n1723) );
  MUX2X1 U1411 ( .B(n1722), .A(n1719), .S(n1974), .Y(n1726) );
  MUX2X1 U1412 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n2000), .Y(n1730) );
  MUX2X1 U1413 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n2000), .Y(n1729) );
  MUX2X1 U1414 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n2000), .Y(n1733) );
  MUX2X1 U1415 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n2000), .Y(n1732) );
  MUX2X1 U1416 ( .B(n1731), .A(n1728), .S(n1974), .Y(n1742) );
  MUX2X1 U1417 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n2000), .Y(n1736) );
  MUX2X1 U1418 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n2000), .Y(n1735) );
  MUX2X1 U1419 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n2000), .Y(n1739) );
  MUX2X1 U1420 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n2000), .Y(n1738) );
  MUX2X1 U1421 ( .B(n1737), .A(n1734), .S(n1974), .Y(n1741) );
  MUX2X1 U1422 ( .B(n1740), .A(n1725), .S(n1969), .Y(n1961) );
  MUX2X1 U1423 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n2000), .Y(n1745) );
  MUX2X1 U1424 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n2000), .Y(n1744) );
  MUX2X1 U1425 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n2000), .Y(n1748) );
  MUX2X1 U1426 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n2000), .Y(n1747) );
  MUX2X1 U1427 ( .B(n1746), .A(n1743), .S(n1973), .Y(n1757) );
  MUX2X1 U1428 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n2001), .Y(n1751) );
  MUX2X1 U1429 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n2001), .Y(n1750) );
  MUX2X1 U1430 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n2001), .Y(n1754) );
  MUX2X1 U1431 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n2001), .Y(n1753) );
  MUX2X1 U1432 ( .B(n1752), .A(n1749), .S(n1973), .Y(n1756) );
  MUX2X1 U1433 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n2001), .Y(n1760) );
  MUX2X1 U1434 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n2001), .Y(n1759) );
  MUX2X1 U1435 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n2001), .Y(n1763) );
  MUX2X1 U1436 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n2001), .Y(n1762) );
  MUX2X1 U1437 ( .B(n1761), .A(n1758), .S(n1973), .Y(n1772) );
  MUX2X1 U1438 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n2001), .Y(n1766) );
  MUX2X1 U1439 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n2001), .Y(n1765) );
  MUX2X1 U1440 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n2001), .Y(n1769) );
  MUX2X1 U1441 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n2001), .Y(n1768) );
  MUX2X1 U1442 ( .B(n1767), .A(n1764), .S(n1973), .Y(n1771) );
  MUX2X1 U1443 ( .B(n1770), .A(n1755), .S(n1969), .Y(n1962) );
  MUX2X1 U1444 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n2002), .Y(n1775) );
  MUX2X1 U1445 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n2002), .Y(n1774) );
  MUX2X1 U1446 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n2002), .Y(n1778) );
  MUX2X1 U1447 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n2002), .Y(n1777) );
  MUX2X1 U1448 ( .B(n1776), .A(n1773), .S(n1973), .Y(n1787) );
  MUX2X1 U1449 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n2002), .Y(n1781) );
  MUX2X1 U1450 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n2002), .Y(n1780) );
  MUX2X1 U1451 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n2002), .Y(n1784) );
  MUX2X1 U1452 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n2002), .Y(n1783) );
  MUX2X1 U1453 ( .B(n1782), .A(n1779), .S(n1973), .Y(n1786) );
  MUX2X1 U1454 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n2002), .Y(n1790) );
  MUX2X1 U1455 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n2002), .Y(n1789) );
  MUX2X1 U1456 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n2002), .Y(n1793) );
  MUX2X1 U1457 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n2002), .Y(n1792) );
  MUX2X1 U1458 ( .B(n1791), .A(n1788), .S(n1973), .Y(n1802) );
  MUX2X1 U1459 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n2003), .Y(n1796) );
  MUX2X1 U1460 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n2003), .Y(n1795) );
  MUX2X1 U1461 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n2003), .Y(n1799) );
  MUX2X1 U1462 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n2003), .Y(n1798) );
  MUX2X1 U1463 ( .B(n1797), .A(n1794), .S(n1973), .Y(n1801) );
  MUX2X1 U1464 ( .B(n1800), .A(n1785), .S(n1969), .Y(n1963) );
  MUX2X1 U1465 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n2003), .Y(n1805) );
  MUX2X1 U1466 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n2003), .Y(n1804) );
  MUX2X1 U1467 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n2003), .Y(n1808) );
  MUX2X1 U1468 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n2003), .Y(n1807) );
  MUX2X1 U1469 ( .B(n1806), .A(n1803), .S(n1973), .Y(n1817) );
  MUX2X1 U1470 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n2003), .Y(n1811) );
  MUX2X1 U1471 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n2003), .Y(n1810) );
  MUX2X1 U1472 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n2003), .Y(n1814) );
  MUX2X1 U1473 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n2003), .Y(n1813) );
  MUX2X1 U1474 ( .B(n1812), .A(n1809), .S(n1973), .Y(n1816) );
  MUX2X1 U1475 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n2004), .Y(n1820) );
  MUX2X1 U1476 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n2004), .Y(n1819) );
  MUX2X1 U1477 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n2004), .Y(n1823) );
  MUX2X1 U1478 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n2004), .Y(n1822) );
  MUX2X1 U1479 ( .B(n1821), .A(n1818), .S(n1973), .Y(n1832) );
  MUX2X1 U1480 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n2004), .Y(n1826) );
  MUX2X1 U1481 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n2004), .Y(n1825) );
  MUX2X1 U1482 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n2004), .Y(n1829) );
  MUX2X1 U1483 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n2004), .Y(n1828) );
  MUX2X1 U1484 ( .B(n1827), .A(n1824), .S(n1973), .Y(n1831) );
  MUX2X1 U1485 ( .B(n1830), .A(n1815), .S(n1969), .Y(n1964) );
  MUX2X1 U1486 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n2004), .Y(n1835) );
  MUX2X1 U1487 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n2004), .Y(n1834) );
  MUX2X1 U1488 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n2004), .Y(n1838) );
  MUX2X1 U1489 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n2004), .Y(n1837) );
  MUX2X1 U1490 ( .B(n1836), .A(n1833), .S(n1973), .Y(n1847) );
  MUX2X1 U1491 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n2005), .Y(n1841) );
  MUX2X1 U1492 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n2005), .Y(n1840) );
  MUX2X1 U1493 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n2005), .Y(n1844) );
  MUX2X1 U1494 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n2005), .Y(n1843) );
  MUX2X1 U1495 ( .B(n1842), .A(n1839), .S(n1973), .Y(n1846) );
  MUX2X1 U1496 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n2005), .Y(n1850) );
  MUX2X1 U1497 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n2005), .Y(n1849) );
  MUX2X1 U1498 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n2005), .Y(n1853) );
  MUX2X1 U1499 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n2005), .Y(n1852) );
  MUX2X1 U1500 ( .B(n1851), .A(n1848), .S(n1973), .Y(n1862) );
  MUX2X1 U1501 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n2005), .Y(n1856) );
  MUX2X1 U1502 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n2005), .Y(n1855) );
  MUX2X1 U1503 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n2005), .Y(n1859) );
  MUX2X1 U1504 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n2005), .Y(n1858) );
  MUX2X1 U1505 ( .B(n1857), .A(n1854), .S(n1973), .Y(n1861) );
  MUX2X1 U1506 ( .B(n1860), .A(n1845), .S(n1969), .Y(n1965) );
  MUX2X1 U1507 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n2006), .Y(n1865) );
  MUX2X1 U1508 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n2006), .Y(n1864) );
  MUX2X1 U1509 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n2006), .Y(n1868) );
  MUX2X1 U1510 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n2006), .Y(n1867) );
  MUX2X1 U1511 ( .B(n1866), .A(n1863), .S(n1973), .Y(n1877) );
  MUX2X1 U1512 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n2006), .Y(n1871) );
  MUX2X1 U1513 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n2006), .Y(n1870) );
  MUX2X1 U1514 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n2006), .Y(n1874) );
  MUX2X1 U1515 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n2006), .Y(n1873) );
  MUX2X1 U1516 ( .B(n1872), .A(n1869), .S(n2112), .Y(n1876) );
  MUX2X1 U1517 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n2006), .Y(n1880) );
  MUX2X1 U1518 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n2006), .Y(n1879) );
  MUX2X1 U1519 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n2006), .Y(n1883) );
  MUX2X1 U1520 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n2006), .Y(n1882) );
  MUX2X1 U1521 ( .B(n1881), .A(n1878), .S(n1973), .Y(n1892) );
  MUX2X1 U1522 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n2007), .Y(n1886) );
  MUX2X1 U1523 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n2007), .Y(n1885) );
  MUX2X1 U1524 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n2007), .Y(n1889) );
  MUX2X1 U1525 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n2007), .Y(n1888) );
  MUX2X1 U1526 ( .B(n1887), .A(n1884), .S(n1973), .Y(n1891) );
  MUX2X1 U1527 ( .B(n1890), .A(n1875), .S(n1969), .Y(n1966) );
  MUX2X1 U1528 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n2007), .Y(n1895) );
  MUX2X1 U1529 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n2007), .Y(n1894) );
  MUX2X1 U1530 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n2007), .Y(n1898) );
  MUX2X1 U1531 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n2007), .Y(n1897) );
  MUX2X1 U1532 ( .B(n1896), .A(n1893), .S(n1973), .Y(n1907) );
  MUX2X1 U1533 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n2007), .Y(n1901) );
  MUX2X1 U1534 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n2007), .Y(n1900) );
  MUX2X1 U1535 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n2007), .Y(n1904) );
  MUX2X1 U1536 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n2007), .Y(n1903) );
  MUX2X1 U1537 ( .B(n1902), .A(n1899), .S(n1973), .Y(n1906) );
  MUX2X1 U1538 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n2008), .Y(n1910) );
  MUX2X1 U1539 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n2008), .Y(n1909) );
  MUX2X1 U1540 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n2008), .Y(n1913) );
  MUX2X1 U1541 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n2008), .Y(n1912) );
  MUX2X1 U1542 ( .B(n1911), .A(n1908), .S(n2112), .Y(n1922) );
  MUX2X1 U1543 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n2008), .Y(n1916) );
  MUX2X1 U1544 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n2008), .Y(n1915) );
  MUX2X1 U1545 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n2008), .Y(n1919) );
  MUX2X1 U1546 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n2008), .Y(n1918) );
  MUX2X1 U1547 ( .B(n1917), .A(n1914), .S(n1973), .Y(n1921) );
  MUX2X1 U1548 ( .B(n1920), .A(n1905), .S(n1969), .Y(n1967) );
  MUX2X1 U1549 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n2008), .Y(n1925) );
  MUX2X1 U1550 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n2008), .Y(n1924) );
  MUX2X1 U1551 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n2008), .Y(n1928) );
  MUX2X1 U1552 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n2008), .Y(n1927) );
  MUX2X1 U1553 ( .B(n1926), .A(n1923), .S(n1974), .Y(n1937) );
  MUX2X1 U1554 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n2009), .Y(n1931) );
  MUX2X1 U1555 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n2009), .Y(n1930) );
  MUX2X1 U1556 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n2009), .Y(n1934) );
  MUX2X1 U1557 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n2009), .Y(n1933) );
  MUX2X1 U1558 ( .B(n1932), .A(n1929), .S(n1973), .Y(n1936) );
  MUX2X1 U1559 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n2009), .Y(n1940) );
  MUX2X1 U1560 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n2009), .Y(n1939) );
  MUX2X1 U1561 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n2009), .Y(n1943) );
  MUX2X1 U1562 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n2009), .Y(n1942) );
  MUX2X1 U1563 ( .B(n1941), .A(n1938), .S(n1973), .Y(n1952) );
  MUX2X1 U1564 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n2009), .Y(n1946) );
  MUX2X1 U1565 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n2009), .Y(n1945) );
  MUX2X1 U1566 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n2009), .Y(n1949) );
  MUX2X1 U1567 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n2009), .Y(n1948) );
  MUX2X1 U1568 ( .B(n1947), .A(n1944), .S(n1973), .Y(n1951) );
  MUX2X1 U1569 ( .B(n1950), .A(n1935), .S(n1969), .Y(n1968) );
  INVX8 U1570 ( .A(n1984), .Y(n1982) );
  INVX8 U1571 ( .A(n2011), .Y(n1985) );
  INVX8 U1572 ( .A(n2012), .Y(n1986) );
  INVX8 U1573 ( .A(n2012), .Y(n1987) );
  INVX8 U1574 ( .A(n1987), .Y(n1988) );
  INVX8 U1575 ( .A(n1987), .Y(n1989) );
  INVX8 U1576 ( .A(n1987), .Y(n1990) );
  INVX8 U1577 ( .A(n1987), .Y(n1991) );
  INVX8 U1578 ( .A(n1987), .Y(n1992) );
  INVX8 U1579 ( .A(n1987), .Y(n1993) );
  INVX8 U1580 ( .A(n1987), .Y(n1994) );
  INVX8 U1581 ( .A(n1987), .Y(n1995) );
  INVX8 U1582 ( .A(n1987), .Y(n1996) );
  INVX8 U1583 ( .A(n1986), .Y(n1997) );
  INVX8 U1584 ( .A(n1986), .Y(n1998) );
  INVX8 U1585 ( .A(n1986), .Y(n1999) );
  INVX8 U1586 ( .A(n1986), .Y(n2000) );
  INVX8 U1587 ( .A(n1986), .Y(n2001) );
  INVX8 U1588 ( .A(n1986), .Y(n2002) );
  INVX8 U1589 ( .A(n2010), .Y(n2003) );
  INVX8 U1590 ( .A(n2010), .Y(n2004) );
  INVX8 U1591 ( .A(n1986), .Y(n2005) );
  INVX8 U1592 ( .A(n1985), .Y(n2006) );
  INVX8 U1593 ( .A(n1985), .Y(n2007) );
  INVX8 U1594 ( .A(n1985), .Y(n2008) );
  INVX8 U1595 ( .A(n1985), .Y(n2009) );
  INVX1 U1596 ( .A(N11), .Y(n2111) );
  INVX1 U1597 ( .A(N10), .Y(n2109) );
  INVX8 U1598 ( .A(n2077), .Y(n2074) );
  INVX8 U1599 ( .A(n2077), .Y(n2075) );
  INVX8 U1600 ( .A(n2077), .Y(n2076) );
  INVX8 U1601 ( .A(n291), .Y(n2077) );
  INVX8 U1602 ( .A(n277), .Y(n2078) );
  INVX8 U1603 ( .A(n277), .Y(n2079) );
  INVX8 U1604 ( .A(n278), .Y(n2080) );
  INVX8 U1605 ( .A(n278), .Y(n2081) );
  INVX8 U1606 ( .A(n279), .Y(n2082) );
  INVX8 U1607 ( .A(n279), .Y(n2083) );
  INVX8 U1608 ( .A(n280), .Y(n2084) );
  INVX8 U1609 ( .A(n280), .Y(n2085) );
  INVX8 U1610 ( .A(n281), .Y(n2086) );
  INVX8 U1611 ( .A(n281), .Y(n2087) );
  INVX8 U1612 ( .A(n282), .Y(n2088) );
  INVX8 U1613 ( .A(n282), .Y(n2089) );
  INVX8 U1614 ( .A(n283), .Y(n2090) );
  INVX8 U1615 ( .A(n283), .Y(n2091) );
  INVX8 U1616 ( .A(n284), .Y(n2092) );
  INVX8 U1617 ( .A(n284), .Y(n2093) );
  INVX8 U1618 ( .A(n285), .Y(n2094) );
  INVX8 U1619 ( .A(n285), .Y(n2095) );
  INVX8 U1620 ( .A(n286), .Y(n2096) );
  INVX8 U1621 ( .A(n286), .Y(n2097) );
  INVX8 U1622 ( .A(n287), .Y(n2098) );
  INVX8 U1623 ( .A(n287), .Y(n2099) );
  INVX8 U1624 ( .A(n288), .Y(n2100) );
  INVX8 U1625 ( .A(n288), .Y(n2101) );
  INVX8 U1626 ( .A(n289), .Y(n2102) );
  INVX8 U1627 ( .A(n289), .Y(n2103) );
  INVX8 U1628 ( .A(n290), .Y(n2104) );
  INVX8 U1629 ( .A(n290), .Y(n2105) );
  OR2X2 U1630 ( .A(write), .B(n2106), .Y(n2117) );
  AND2X2 U1631 ( .A(N32), .B(n1472), .Y(\data_out<0> ) );
  AND2X2 U1632 ( .A(n1472), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U1633 ( .A(N30), .B(n292), .Y(\data_out<2> ) );
  AND2X2 U1634 ( .A(N29), .B(n292), .Y(\data_out<3> ) );
  AND2X2 U1635 ( .A(n2118), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U1636 ( .A(N27), .B(n292), .Y(\data_out<5> ) );
  AND2X2 U1637 ( .A(n1470), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U1638 ( .A(N25), .B(n2118), .Y(\data_out<7> ) );
  AND2X2 U1639 ( .A(N24), .B(n292), .Y(\data_out<8> ) );
  AND2X2 U1640 ( .A(N23), .B(n1470), .Y(\data_out<9> ) );
  AND2X2 U1641 ( .A(N22), .B(n1471), .Y(\data_out<10> ) );
  AND2X2 U1642 ( .A(n1444), .B(n1469), .Y(\data_out<11> ) );
  AND2X2 U1643 ( .A(n1470), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U1644 ( .A(n1471), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U1645 ( .A(n2118), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U1646 ( .A(N17), .B(n1472), .Y(\data_out<15> ) );
  OAI21X1 U1647 ( .A(n2014), .B(n2078), .C(n2), .Y(n2772) );
  OAI21X1 U1648 ( .A(n2081), .B(n2013), .C(n4), .Y(n2771) );
  OAI21X1 U1649 ( .A(n2083), .B(n2013), .C(n6), .Y(n2770) );
  OAI21X1 U1650 ( .A(n2085), .B(n2013), .C(n8), .Y(n2769) );
  OAI21X1 U1651 ( .A(n2087), .B(n2013), .C(n10), .Y(n2768) );
  OAI21X1 U1652 ( .A(n2089), .B(n2013), .C(n12), .Y(n2767) );
  OAI21X1 U1653 ( .A(n2091), .B(n2013), .C(n14), .Y(n2766) );
  NAND2X1 U1654 ( .A(\mem<31><7> ), .B(n209), .Y(n2119) );
  OAI21X1 U1655 ( .A(n275), .B(n2013), .C(n2119), .Y(n2765) );
  NAND2X1 U1656 ( .A(\mem<31><8> ), .B(n209), .Y(n2120) );
  OAI21X1 U1657 ( .A(n2093), .B(n2013), .C(n2120), .Y(n2764) );
  NAND2X1 U1658 ( .A(\mem<31><9> ), .B(n209), .Y(n2121) );
  OAI21X1 U1659 ( .A(n2095), .B(n2014), .C(n2121), .Y(n2763) );
  NAND2X1 U1660 ( .A(\mem<31><10> ), .B(n209), .Y(n2122) );
  OAI21X1 U1661 ( .A(n2097), .B(n2014), .C(n2122), .Y(n2762) );
  NAND2X1 U1662 ( .A(\mem<31><11> ), .B(n209), .Y(n2123) );
  OAI21X1 U1663 ( .A(n2099), .B(n2014), .C(n2123), .Y(n2761) );
  NAND2X1 U1664 ( .A(\mem<31><12> ), .B(n209), .Y(n2124) );
  OAI21X1 U1665 ( .A(n2101), .B(n2014), .C(n2124), .Y(n2760) );
  NAND2X1 U1666 ( .A(\mem<31><13> ), .B(n209), .Y(n2125) );
  OAI21X1 U1667 ( .A(n2103), .B(n2014), .C(n2125), .Y(n2759) );
  NAND2X1 U1668 ( .A(\mem<31><14> ), .B(n209), .Y(n2126) );
  OAI21X1 U1669 ( .A(n2105), .B(n2014), .C(n2126), .Y(n2758) );
  NAND2X1 U1670 ( .A(\mem<31><15> ), .B(n209), .Y(n2127) );
  OAI21X1 U1671 ( .A(n1457), .B(n2014), .C(n2127), .Y(n2757) );
  NAND2X1 U1672 ( .A(\mem<30><0> ), .B(n211), .Y(n2128) );
  OAI21X1 U1673 ( .A(n2015), .B(n2078), .C(n2128), .Y(n2756) );
  NAND2X1 U1674 ( .A(\mem<30><1> ), .B(n211), .Y(n2129) );
  OAI21X1 U1675 ( .A(n2015), .B(n2081), .C(n2129), .Y(n2755) );
  NAND2X1 U1676 ( .A(\mem<30><2> ), .B(n211), .Y(n2130) );
  OAI21X1 U1677 ( .A(n2015), .B(n2083), .C(n2130), .Y(n2754) );
  NAND2X1 U1678 ( .A(\mem<30><3> ), .B(n211), .Y(n2131) );
  OAI21X1 U1679 ( .A(n2015), .B(n2085), .C(n2131), .Y(n2753) );
  NAND2X1 U1680 ( .A(\mem<30><4> ), .B(n211), .Y(n2132) );
  OAI21X1 U1681 ( .A(n2015), .B(n2087), .C(n2132), .Y(n2752) );
  NAND2X1 U1682 ( .A(\mem<30><5> ), .B(n211), .Y(n2133) );
  OAI21X1 U1683 ( .A(n2015), .B(n2089), .C(n2133), .Y(n2751) );
  NAND2X1 U1684 ( .A(\mem<30><6> ), .B(n211), .Y(n2134) );
  OAI21X1 U1685 ( .A(n2015), .B(n2091), .C(n2134), .Y(n2750) );
  NAND2X1 U1686 ( .A(\mem<30><7> ), .B(n211), .Y(n2135) );
  OAI21X1 U1687 ( .A(n2015), .B(n1446), .C(n2135), .Y(n2749) );
  OAI21X1 U1688 ( .A(n2016), .B(n2092), .C(n16), .Y(n2748) );
  OAI21X1 U1689 ( .A(n2016), .B(n2094), .C(n18), .Y(n2747) );
  OAI21X1 U1690 ( .A(n2016), .B(n2096), .C(n20), .Y(n2746) );
  OAI21X1 U1691 ( .A(n2016), .B(n2098), .C(n22), .Y(n2745) );
  OAI21X1 U1692 ( .A(n2016), .B(n2100), .C(n24), .Y(n2744) );
  OAI21X1 U1693 ( .A(n2016), .B(n2102), .C(n26), .Y(n2743) );
  OAI21X1 U1694 ( .A(n2016), .B(n2104), .C(n28), .Y(n2742) );
  NAND2X1 U1695 ( .A(\mem<30><15> ), .B(n211), .Y(n2136) );
  OAI21X1 U1696 ( .A(n2016), .B(n1462), .C(n2136), .Y(n2741) );
  NAND3X1 U1697 ( .A(n2108), .B(n2112), .C(n2111), .Y(n2137) );
  NAND2X1 U1698 ( .A(\mem<29><0> ), .B(n213), .Y(n2138) );
  OAI21X1 U1699 ( .A(n2017), .B(n2078), .C(n2138), .Y(n2740) );
  NAND2X1 U1700 ( .A(\mem<29><1> ), .B(n213), .Y(n2139) );
  OAI21X1 U1701 ( .A(n2017), .B(n2080), .C(n2139), .Y(n2739) );
  NAND2X1 U1702 ( .A(\mem<29><2> ), .B(n213), .Y(n2140) );
  OAI21X1 U1703 ( .A(n2017), .B(n2082), .C(n2140), .Y(n2738) );
  NAND2X1 U1704 ( .A(\mem<29><3> ), .B(n213), .Y(n2141) );
  OAI21X1 U1705 ( .A(n2017), .B(n2084), .C(n2141), .Y(n2737) );
  NAND2X1 U1706 ( .A(\mem<29><4> ), .B(n213), .Y(n2142) );
  OAI21X1 U1707 ( .A(n2017), .B(n2086), .C(n2142), .Y(n2736) );
  NAND2X1 U1708 ( .A(\mem<29><5> ), .B(n213), .Y(n2143) );
  OAI21X1 U1709 ( .A(n2017), .B(n2088), .C(n2143), .Y(n2735) );
  NAND2X1 U1710 ( .A(\mem<29><6> ), .B(n213), .Y(n2144) );
  OAI21X1 U1711 ( .A(n2017), .B(n2090), .C(n2144), .Y(n2734) );
  NAND2X1 U1712 ( .A(\mem<29><7> ), .B(n213), .Y(n2145) );
  OAI21X1 U1713 ( .A(n2017), .B(n1447), .C(n2145), .Y(n2733) );
  OAI21X1 U1714 ( .A(n2018), .B(n2093), .C(n30), .Y(n2732) );
  OAI21X1 U1715 ( .A(n2018), .B(n2095), .C(n32), .Y(n2731) );
  OAI21X1 U1716 ( .A(n2018), .B(n2097), .C(n34), .Y(n2730) );
  OAI21X1 U1717 ( .A(n2018), .B(n2099), .C(n36), .Y(n2729) );
  OAI21X1 U1718 ( .A(n2018), .B(n2101), .C(n38), .Y(n2728) );
  OAI21X1 U1719 ( .A(n2018), .B(n2103), .C(n40), .Y(n2727) );
  OAI21X1 U1720 ( .A(n2018), .B(n2105), .C(n42), .Y(n2726) );
  NAND2X1 U1721 ( .A(\mem<29><15> ), .B(n213), .Y(n2146) );
  OAI21X1 U1722 ( .A(n2018), .B(n1451), .C(n2146), .Y(n2725) );
  NAND3X1 U1723 ( .A(n2112), .B(n2111), .C(n2109), .Y(n2147) );
  NAND2X1 U1724 ( .A(\mem<28><0> ), .B(n216), .Y(n2148) );
  OAI21X1 U1725 ( .A(n2019), .B(n2078), .C(n2148), .Y(n2724) );
  NAND2X1 U1726 ( .A(\mem<28><1> ), .B(n216), .Y(n2149) );
  OAI21X1 U1727 ( .A(n2019), .B(n2081), .C(n2149), .Y(n2723) );
  NAND2X1 U1728 ( .A(\mem<28><2> ), .B(n216), .Y(n2150) );
  OAI21X1 U1729 ( .A(n2019), .B(n2083), .C(n2150), .Y(n2722) );
  NAND2X1 U1730 ( .A(\mem<28><3> ), .B(n216), .Y(n2151) );
  OAI21X1 U1731 ( .A(n2019), .B(n2085), .C(n2151), .Y(n2721) );
  NAND2X1 U1732 ( .A(\mem<28><4> ), .B(n216), .Y(n2152) );
  OAI21X1 U1733 ( .A(n2019), .B(n2087), .C(n2152), .Y(n2720) );
  NAND2X1 U1734 ( .A(\mem<28><5> ), .B(n216), .Y(n2153) );
  OAI21X1 U1735 ( .A(n2019), .B(n2089), .C(n2153), .Y(n2719) );
  NAND2X1 U1736 ( .A(\mem<28><6> ), .B(n216), .Y(n2154) );
  OAI21X1 U1737 ( .A(n2019), .B(n2091), .C(n2154), .Y(n2718) );
  NAND2X1 U1738 ( .A(\mem<28><7> ), .B(n216), .Y(n2155) );
  OAI21X1 U1739 ( .A(n2019), .B(n1448), .C(n2155), .Y(n2717) );
  OAI21X1 U1740 ( .A(n2020), .B(n2092), .C(n44), .Y(n2716) );
  OAI21X1 U1741 ( .A(n2020), .B(n2094), .C(n46), .Y(n2715) );
  OAI21X1 U1742 ( .A(n2020), .B(n2096), .C(n48), .Y(n2714) );
  OAI21X1 U1743 ( .A(n2020), .B(n2098), .C(n50), .Y(n2713) );
  OAI21X1 U1744 ( .A(n2020), .B(n2100), .C(n52), .Y(n2712) );
  OAI21X1 U1745 ( .A(n2020), .B(n2102), .C(n54), .Y(n2711) );
  OAI21X1 U1746 ( .A(n2020), .B(n2104), .C(n56), .Y(n2710) );
  NAND2X1 U1747 ( .A(\mem<28><15> ), .B(n216), .Y(n2156) );
  OAI21X1 U1748 ( .A(n2020), .B(n1452), .C(n2156), .Y(n2709) );
  NAND3X1 U1749 ( .A(n2108), .B(n2110), .C(n2113), .Y(n2157) );
  NAND2X1 U1750 ( .A(\mem<27><0> ), .B(n218), .Y(n2158) );
  OAI21X1 U1751 ( .A(n2021), .B(n2078), .C(n2158), .Y(n2708) );
  NAND2X1 U1752 ( .A(\mem<27><1> ), .B(n218), .Y(n2159) );
  OAI21X1 U1753 ( .A(n2021), .B(n2080), .C(n2159), .Y(n2707) );
  NAND2X1 U1754 ( .A(\mem<27><2> ), .B(n218), .Y(n2160) );
  OAI21X1 U1755 ( .A(n2021), .B(n2082), .C(n2160), .Y(n2706) );
  NAND2X1 U1756 ( .A(\mem<27><3> ), .B(n218), .Y(n2161) );
  OAI21X1 U1757 ( .A(n2021), .B(n2084), .C(n2161), .Y(n2705) );
  NAND2X1 U1758 ( .A(\mem<27><4> ), .B(n218), .Y(n2162) );
  OAI21X1 U1759 ( .A(n2021), .B(n2086), .C(n2162), .Y(n2704) );
  NAND2X1 U1760 ( .A(\mem<27><5> ), .B(n218), .Y(n2163) );
  OAI21X1 U1761 ( .A(n2021), .B(n2088), .C(n2163), .Y(n2703) );
  NAND2X1 U1762 ( .A(\mem<27><6> ), .B(n218), .Y(n2164) );
  OAI21X1 U1763 ( .A(n2021), .B(n2090), .C(n2164), .Y(n2702) );
  NAND2X1 U1764 ( .A(\mem<27><7> ), .B(n218), .Y(n2165) );
  OAI21X1 U1765 ( .A(n2021), .B(n1449), .C(n2165), .Y(n2701) );
  OAI21X1 U1766 ( .A(n2022), .B(n2093), .C(n58), .Y(n2700) );
  OAI21X1 U1767 ( .A(n2022), .B(n2095), .C(n60), .Y(n2699) );
  OAI21X1 U1768 ( .A(n2022), .B(n2097), .C(n62), .Y(n2698) );
  OAI21X1 U1769 ( .A(n2022), .B(n2099), .C(n64), .Y(n2697) );
  OAI21X1 U1770 ( .A(n2022), .B(n2101), .C(n66), .Y(n2696) );
  OAI21X1 U1771 ( .A(n2022), .B(n2103), .C(n68), .Y(n2695) );
  OAI21X1 U1772 ( .A(n2022), .B(n2105), .C(n70), .Y(n2694) );
  NAND2X1 U1773 ( .A(\mem<27><15> ), .B(n218), .Y(n2166) );
  OAI21X1 U1774 ( .A(n2022), .B(n1453), .C(n2166), .Y(n2693) );
  NAND3X1 U1775 ( .A(n2113), .B(n2110), .C(n2109), .Y(n2167) );
  NAND2X1 U1776 ( .A(\mem<26><0> ), .B(n220), .Y(n2168) );
  OAI21X1 U1777 ( .A(n2023), .B(n2078), .C(n2168), .Y(n2692) );
  NAND2X1 U1778 ( .A(\mem<26><1> ), .B(n220), .Y(n2169) );
  OAI21X1 U1779 ( .A(n2023), .B(n2081), .C(n2169), .Y(n2691) );
  NAND2X1 U1780 ( .A(\mem<26><2> ), .B(n220), .Y(n2170) );
  OAI21X1 U1781 ( .A(n2023), .B(n2083), .C(n2170), .Y(n2690) );
  NAND2X1 U1782 ( .A(\mem<26><3> ), .B(n220), .Y(n2171) );
  OAI21X1 U1783 ( .A(n2023), .B(n2085), .C(n2171), .Y(n2689) );
  NAND2X1 U1784 ( .A(\mem<26><4> ), .B(n220), .Y(n2172) );
  OAI21X1 U1785 ( .A(n2023), .B(n2087), .C(n2172), .Y(n2688) );
  NAND2X1 U1786 ( .A(\mem<26><5> ), .B(n220), .Y(n2173) );
  OAI21X1 U1787 ( .A(n2023), .B(n2089), .C(n2173), .Y(n2687) );
  NAND2X1 U1788 ( .A(\mem<26><6> ), .B(n220), .Y(n2174) );
  OAI21X1 U1789 ( .A(n2023), .B(n2091), .C(n2174), .Y(n2686) );
  NAND2X1 U1790 ( .A(\mem<26><7> ), .B(n220), .Y(n2175) );
  OAI21X1 U1791 ( .A(n2023), .B(n1450), .C(n2175), .Y(n2685) );
  OAI21X1 U1792 ( .A(n2024), .B(n2092), .C(n72), .Y(n2684) );
  OAI21X1 U1793 ( .A(n2024), .B(n2094), .C(n74), .Y(n2683) );
  OAI21X1 U1794 ( .A(n2024), .B(n2096), .C(n76), .Y(n2682) );
  OAI21X1 U1795 ( .A(n2024), .B(n2098), .C(n78), .Y(n2681) );
  OAI21X1 U1796 ( .A(n2024), .B(n2100), .C(n80), .Y(n2680) );
  OAI21X1 U1797 ( .A(n2024), .B(n2102), .C(n82), .Y(n2679) );
  OAI21X1 U1798 ( .A(n2024), .B(n2104), .C(n84), .Y(n2678) );
  NAND2X1 U1799 ( .A(\mem<26><15> ), .B(n220), .Y(n2176) );
  OAI21X1 U1800 ( .A(n2024), .B(n1452), .C(n2176), .Y(n2677) );
  NAND3X1 U1801 ( .A(n2108), .B(n2113), .C(n2111), .Y(n2177) );
  NAND2X1 U1802 ( .A(\mem<25><0> ), .B(n222), .Y(n2178) );
  OAI21X1 U1803 ( .A(n2025), .B(n2078), .C(n2178), .Y(n2676) );
  NAND2X1 U1804 ( .A(\mem<25><1> ), .B(n222), .Y(n2179) );
  OAI21X1 U1805 ( .A(n2025), .B(n2080), .C(n2179), .Y(n2675) );
  NAND2X1 U1806 ( .A(\mem<25><2> ), .B(n222), .Y(n2180) );
  OAI21X1 U1807 ( .A(n2025), .B(n2082), .C(n2180), .Y(n2674) );
  NAND2X1 U1808 ( .A(\mem<25><3> ), .B(n222), .Y(n2181) );
  OAI21X1 U1809 ( .A(n2025), .B(n2084), .C(n2181), .Y(n2673) );
  NAND2X1 U1810 ( .A(\mem<25><4> ), .B(n222), .Y(n2182) );
  OAI21X1 U1811 ( .A(n2025), .B(n2086), .C(n2182), .Y(n2672) );
  NAND2X1 U1812 ( .A(\mem<25><5> ), .B(n222), .Y(n2183) );
  OAI21X1 U1813 ( .A(n2025), .B(n2088), .C(n2183), .Y(n2671) );
  NAND2X1 U1814 ( .A(\mem<25><6> ), .B(n222), .Y(n2184) );
  OAI21X1 U1815 ( .A(n2025), .B(n2090), .C(n2184), .Y(n2670) );
  NAND2X1 U1816 ( .A(\mem<25><7> ), .B(n222), .Y(n2185) );
  OAI21X1 U1817 ( .A(n2025), .B(n1448), .C(n2185), .Y(n2669) );
  OAI21X1 U1818 ( .A(n2026), .B(n2093), .C(n86), .Y(n2668) );
  OAI21X1 U1819 ( .A(n2026), .B(n2095), .C(n88), .Y(n2667) );
  OAI21X1 U1820 ( .A(n2026), .B(n2097), .C(n90), .Y(n2666) );
  OAI21X1 U1821 ( .A(n2026), .B(n2099), .C(n92), .Y(n2665) );
  OAI21X1 U1822 ( .A(n2026), .B(n2101), .C(n94), .Y(n2664) );
  OAI21X1 U1823 ( .A(n2026), .B(n2103), .C(n96), .Y(n2663) );
  OAI21X1 U1824 ( .A(n2026), .B(n2105), .C(n98), .Y(n2662) );
  NAND2X1 U1825 ( .A(\mem<25><15> ), .B(n222), .Y(n2186) );
  OAI21X1 U1826 ( .A(n2026), .B(n1454), .C(n2186), .Y(n2661) );
  NOR3X1 U1827 ( .A(n2108), .B(n2110), .C(n2112), .Y(n2258) );
  NAND2X1 U1828 ( .A(\mem<24><0> ), .B(n224), .Y(n2187) );
  OAI21X1 U1829 ( .A(n2027), .B(n2078), .C(n2187), .Y(n2660) );
  NAND2X1 U1830 ( .A(\mem<24><1> ), .B(n224), .Y(n2188) );
  OAI21X1 U1831 ( .A(n2027), .B(n2080), .C(n2188), .Y(n2659) );
  NAND2X1 U1832 ( .A(\mem<24><2> ), .B(n224), .Y(n2189) );
  OAI21X1 U1833 ( .A(n2027), .B(n2082), .C(n2189), .Y(n2658) );
  NAND2X1 U1834 ( .A(\mem<24><3> ), .B(n224), .Y(n2190) );
  OAI21X1 U1835 ( .A(n2027), .B(n2084), .C(n2190), .Y(n2657) );
  NAND2X1 U1836 ( .A(\mem<24><4> ), .B(n224), .Y(n2191) );
  OAI21X1 U1837 ( .A(n2027), .B(n2086), .C(n2191), .Y(n2656) );
  NAND2X1 U1838 ( .A(\mem<24><5> ), .B(n224), .Y(n2192) );
  OAI21X1 U1839 ( .A(n2027), .B(n2088), .C(n2192), .Y(n2655) );
  NAND2X1 U1840 ( .A(\mem<24><6> ), .B(n224), .Y(n2193) );
  OAI21X1 U1841 ( .A(n2027), .B(n2090), .C(n2193), .Y(n2654) );
  NAND2X1 U1842 ( .A(\mem<24><7> ), .B(n224), .Y(n2194) );
  OAI21X1 U1843 ( .A(n2027), .B(n275), .C(n2194), .Y(n2653) );
  OAI21X1 U1844 ( .A(n2027), .B(n2092), .C(n100), .Y(n2652) );
  OAI21X1 U1845 ( .A(n2027), .B(n2094), .C(n102), .Y(n2651) );
  OAI21X1 U1846 ( .A(n2027), .B(n2096), .C(n104), .Y(n2650) );
  OAI21X1 U1847 ( .A(n2027), .B(n2098), .C(n106), .Y(n2649) );
  OAI21X1 U1848 ( .A(n2027), .B(n2100), .C(n108), .Y(n2648) );
  OAI21X1 U1849 ( .A(n2027), .B(n2102), .C(n110), .Y(n2647) );
  NAND2X1 U1850 ( .A(\mem<24><14> ), .B(n224), .Y(n2195) );
  OAI21X1 U1851 ( .A(n2027), .B(n2104), .C(n2195), .Y(n2646) );
  OAI21X1 U1852 ( .A(n2027), .B(n1465), .C(n112), .Y(n2645) );
  NAND2X1 U1853 ( .A(\mem<23><0> ), .B(n226), .Y(n2196) );
  OAI21X1 U1854 ( .A(n2028), .B(n2078), .C(n2196), .Y(n2644) );
  NAND2X1 U1855 ( .A(\mem<23><1> ), .B(n226), .Y(n2197) );
  OAI21X1 U1856 ( .A(n2028), .B(n2081), .C(n2197), .Y(n2643) );
  NAND2X1 U1857 ( .A(\mem<23><2> ), .B(n226), .Y(n2198) );
  OAI21X1 U1858 ( .A(n2028), .B(n2083), .C(n2198), .Y(n2642) );
  NAND2X1 U1859 ( .A(\mem<23><3> ), .B(n226), .Y(n2199) );
  OAI21X1 U1860 ( .A(n2028), .B(n2085), .C(n2199), .Y(n2641) );
  NAND2X1 U1861 ( .A(\mem<23><4> ), .B(n226), .Y(n2200) );
  OAI21X1 U1862 ( .A(n2028), .B(n2087), .C(n2200), .Y(n2640) );
  NAND2X1 U1863 ( .A(\mem<23><5> ), .B(n226), .Y(n2201) );
  OAI21X1 U1864 ( .A(n2028), .B(n2089), .C(n2201), .Y(n2639) );
  NAND2X1 U1865 ( .A(\mem<23><6> ), .B(n226), .Y(n2202) );
  OAI21X1 U1866 ( .A(n2028), .B(n2091), .C(n2202), .Y(n2638) );
  NAND2X1 U1867 ( .A(\mem<23><7> ), .B(n226), .Y(n2203) );
  OAI21X1 U1868 ( .A(n2028), .B(n1449), .C(n2203), .Y(n2637) );
  OAI21X1 U1869 ( .A(n2029), .B(n2093), .C(n114), .Y(n2636) );
  OAI21X1 U1870 ( .A(n2029), .B(n2095), .C(n116), .Y(n2635) );
  OAI21X1 U1871 ( .A(n2029), .B(n2097), .C(n118), .Y(n2634) );
  OAI21X1 U1872 ( .A(n2029), .B(n2099), .C(n120), .Y(n2633) );
  OAI21X1 U1873 ( .A(n2029), .B(n2101), .C(n122), .Y(n2632) );
  OAI21X1 U1874 ( .A(n2029), .B(n2103), .C(n124), .Y(n2631) );
  OAI21X1 U1875 ( .A(n2029), .B(n2105), .C(n126), .Y(n2630) );
  NAND2X1 U1876 ( .A(\mem<23><15> ), .B(n226), .Y(n2204) );
  OAI21X1 U1877 ( .A(n2029), .B(n1465), .C(n2204), .Y(n2629) );
  NAND2X1 U1878 ( .A(\mem<22><0> ), .B(n228), .Y(n2205) );
  OAI21X1 U1879 ( .A(n2030), .B(n2078), .C(n2205), .Y(n2628) );
  NAND2X1 U1880 ( .A(\mem<22><1> ), .B(n228), .Y(n2206) );
  OAI21X1 U1881 ( .A(n2030), .B(n2081), .C(n2206), .Y(n2627) );
  NAND2X1 U1882 ( .A(\mem<22><2> ), .B(n228), .Y(n2207) );
  OAI21X1 U1883 ( .A(n2030), .B(n2083), .C(n2207), .Y(n2626) );
  NAND2X1 U1884 ( .A(\mem<22><3> ), .B(n228), .Y(n2208) );
  OAI21X1 U1885 ( .A(n2030), .B(n2085), .C(n2208), .Y(n2625) );
  NAND2X1 U1886 ( .A(\mem<22><4> ), .B(n228), .Y(n2209) );
  OAI21X1 U1887 ( .A(n2030), .B(n2087), .C(n2209), .Y(n2624) );
  NAND2X1 U1888 ( .A(\mem<22><5> ), .B(n228), .Y(n2210) );
  OAI21X1 U1889 ( .A(n2030), .B(n2089), .C(n2210), .Y(n2623) );
  NAND2X1 U1890 ( .A(\mem<22><6> ), .B(n228), .Y(n2211) );
  OAI21X1 U1891 ( .A(n2030), .B(n2091), .C(n2211), .Y(n2622) );
  NAND2X1 U1892 ( .A(\mem<22><7> ), .B(n228), .Y(n2212) );
  OAI21X1 U1893 ( .A(n2030), .B(n1448), .C(n2212), .Y(n2621) );
  OAI21X1 U1894 ( .A(n2031), .B(n2093), .C(n128), .Y(n2620) );
  OAI21X1 U1895 ( .A(n2031), .B(n2095), .C(n130), .Y(n2619) );
  OAI21X1 U1896 ( .A(n2031), .B(n2097), .C(n132), .Y(n2618) );
  OAI21X1 U1897 ( .A(n2031), .B(n2099), .C(n134), .Y(n2617) );
  OAI21X1 U1898 ( .A(n2031), .B(n2101), .C(n136), .Y(n2616) );
  OAI21X1 U1899 ( .A(n2031), .B(n2103), .C(n138), .Y(n2615) );
  OAI21X1 U1900 ( .A(n2031), .B(n2105), .C(n140), .Y(n2614) );
  NAND2X1 U1901 ( .A(\mem<22><15> ), .B(n228), .Y(n2213) );
  OAI21X1 U1902 ( .A(n2031), .B(n1466), .C(n2213), .Y(n2613) );
  NAND2X1 U1903 ( .A(\mem<21><0> ), .B(n230), .Y(n2214) );
  OAI21X1 U1904 ( .A(n2032), .B(n2078), .C(n2214), .Y(n2612) );
  NAND2X1 U1905 ( .A(\mem<21><1> ), .B(n230), .Y(n2215) );
  OAI21X1 U1906 ( .A(n2032), .B(n2081), .C(n2215), .Y(n2611) );
  NAND2X1 U1907 ( .A(\mem<21><2> ), .B(n230), .Y(n2216) );
  OAI21X1 U1908 ( .A(n2032), .B(n2083), .C(n2216), .Y(n2610) );
  NAND2X1 U1909 ( .A(\mem<21><3> ), .B(n230), .Y(n2217) );
  OAI21X1 U1910 ( .A(n2032), .B(n2085), .C(n2217), .Y(n2609) );
  NAND2X1 U1911 ( .A(\mem<21><4> ), .B(n230), .Y(n2218) );
  OAI21X1 U1912 ( .A(n2032), .B(n2087), .C(n2218), .Y(n2608) );
  NAND2X1 U1913 ( .A(\mem<21><5> ), .B(n230), .Y(n2219) );
  OAI21X1 U1914 ( .A(n2032), .B(n2089), .C(n2219), .Y(n2607) );
  NAND2X1 U1915 ( .A(\mem<21><6> ), .B(n230), .Y(n2220) );
  OAI21X1 U1916 ( .A(n2032), .B(n2091), .C(n2220), .Y(n2606) );
  NAND2X1 U1917 ( .A(\mem<21><7> ), .B(n230), .Y(n2221) );
  OAI21X1 U1918 ( .A(n2032), .B(n1445), .C(n2221), .Y(n2605) );
  OAI21X1 U1919 ( .A(n2033), .B(n2093), .C(n142), .Y(n2604) );
  OAI21X1 U1920 ( .A(n2033), .B(n2095), .C(n144), .Y(n2603) );
  OAI21X1 U1921 ( .A(n2033), .B(n2097), .C(n146), .Y(n2602) );
  OAI21X1 U1922 ( .A(n2033), .B(n2099), .C(n148), .Y(n2601) );
  OAI21X1 U1923 ( .A(n2033), .B(n2101), .C(n150), .Y(n2600) );
  OAI21X1 U1924 ( .A(n2033), .B(n2103), .C(n152), .Y(n2599) );
  OAI21X1 U1925 ( .A(n2033), .B(n2105), .C(n154), .Y(n2598) );
  NAND2X1 U1926 ( .A(\mem<21><15> ), .B(n230), .Y(n2222) );
  OAI21X1 U1927 ( .A(n2033), .B(n1467), .C(n2222), .Y(n2597) );
  NAND2X1 U1928 ( .A(\mem<20><0> ), .B(n232), .Y(n2223) );
  OAI21X1 U1929 ( .A(n2034), .B(n2078), .C(n2223), .Y(n2596) );
  NAND2X1 U1930 ( .A(\mem<20><1> ), .B(n232), .Y(n2224) );
  OAI21X1 U1931 ( .A(n2034), .B(n2081), .C(n2224), .Y(n2595) );
  NAND2X1 U1932 ( .A(\mem<20><2> ), .B(n232), .Y(n2225) );
  OAI21X1 U1933 ( .A(n2034), .B(n2083), .C(n2225), .Y(n2594) );
  NAND2X1 U1934 ( .A(\mem<20><3> ), .B(n232), .Y(n2226) );
  OAI21X1 U1935 ( .A(n2034), .B(n2085), .C(n2226), .Y(n2593) );
  NAND2X1 U1936 ( .A(\mem<20><4> ), .B(n232), .Y(n2227) );
  OAI21X1 U1937 ( .A(n2034), .B(n2087), .C(n2227), .Y(n2592) );
  NAND2X1 U1938 ( .A(\mem<20><5> ), .B(n232), .Y(n2228) );
  OAI21X1 U1939 ( .A(n2034), .B(n2089), .C(n2228), .Y(n2591) );
  NAND2X1 U1940 ( .A(\mem<20><6> ), .B(n232), .Y(n2229) );
  OAI21X1 U1941 ( .A(n2034), .B(n2091), .C(n2229), .Y(n2590) );
  NAND2X1 U1942 ( .A(\mem<20><7> ), .B(n232), .Y(n2230) );
  OAI21X1 U1943 ( .A(n2034), .B(n1447), .C(n2230), .Y(n2589) );
  OAI21X1 U1944 ( .A(n2035), .B(n2093), .C(n156), .Y(n2588) );
  OAI21X1 U1945 ( .A(n2035), .B(n2095), .C(n158), .Y(n2587) );
  OAI21X1 U1946 ( .A(n2035), .B(n2097), .C(n160), .Y(n2586) );
  OAI21X1 U1947 ( .A(n2035), .B(n2099), .C(n162), .Y(n2585) );
  OAI21X1 U1948 ( .A(n2035), .B(n2101), .C(n164), .Y(n2584) );
  OAI21X1 U1949 ( .A(n2035), .B(n2103), .C(n166), .Y(n2583) );
  OAI21X1 U1950 ( .A(n2035), .B(n2105), .C(n168), .Y(n2582) );
  NAND2X1 U1951 ( .A(\mem<20><15> ), .B(n232), .Y(n2231) );
  OAI21X1 U1952 ( .A(n2035), .B(n1468), .C(n2231), .Y(n2581) );
  OAI21X1 U1953 ( .A(n2036), .B(n2079), .C(n298), .Y(n2580) );
  OAI21X1 U1954 ( .A(n2036), .B(n2081), .C(n300), .Y(n2579) );
  OAI21X1 U1955 ( .A(n2036), .B(n2083), .C(n302), .Y(n2578) );
  OAI21X1 U1956 ( .A(n2036), .B(n2085), .C(n304), .Y(n2577) );
  OAI21X1 U1957 ( .A(n2036), .B(n2087), .C(n306), .Y(n2576) );
  OAI21X1 U1958 ( .A(n2036), .B(n2089), .C(n308), .Y(n2575) );
  OAI21X1 U1959 ( .A(n2036), .B(n2091), .C(n310), .Y(n2574) );
  OAI21X1 U1960 ( .A(n2036), .B(n1446), .C(n235), .Y(n2573) );
  OAI21X1 U1961 ( .A(n2037), .B(n2093), .C(n312), .Y(n2572) );
  OAI21X1 U1962 ( .A(n2037), .B(n2095), .C(n314), .Y(n2571) );
  OAI21X1 U1963 ( .A(n2037), .B(n2097), .C(n316), .Y(n2570) );
  OAI21X1 U1964 ( .A(n2037), .B(n2099), .C(n318), .Y(n2569) );
  OAI21X1 U1965 ( .A(n2037), .B(n2101), .C(n320), .Y(n2568) );
  OAI21X1 U1966 ( .A(n2037), .B(n2103), .C(n322), .Y(n2567) );
  OAI21X1 U1967 ( .A(n2037), .B(n2105), .C(n324), .Y(n2566) );
  OAI21X1 U1968 ( .A(n2037), .B(n1451), .C(n237), .Y(n2565) );
  OAI21X1 U1969 ( .A(n2039), .B(n2079), .C(n326), .Y(n2564) );
  OAI21X1 U1970 ( .A(n2039), .B(n2081), .C(n328), .Y(n2563) );
  OAI21X1 U1971 ( .A(n2039), .B(n2083), .C(n330), .Y(n2562) );
  OAI21X1 U1972 ( .A(n2039), .B(n2085), .C(n332), .Y(n2561) );
  OAI21X1 U1973 ( .A(n2039), .B(n2087), .C(n334), .Y(n2560) );
  OAI21X1 U1974 ( .A(n2039), .B(n2089), .C(n336), .Y(n2559) );
  OAI21X1 U1975 ( .A(n2039), .B(n2091), .C(n338), .Y(n2558) );
  NAND2X1 U1976 ( .A(\mem<18><7> ), .B(n186), .Y(n2232) );
  OAI21X1 U1977 ( .A(n2039), .B(n207), .C(n2232), .Y(n2557) );
  OAI21X1 U1978 ( .A(n2040), .B(n2093), .C(n340), .Y(n2556) );
  OAI21X1 U1979 ( .A(n2040), .B(n2095), .C(n342), .Y(n2555) );
  OAI21X1 U1980 ( .A(n2040), .B(n2097), .C(n344), .Y(n2554) );
  OAI21X1 U1981 ( .A(n2040), .B(n2099), .C(n346), .Y(n2553) );
  OAI21X1 U1982 ( .A(n2040), .B(n2101), .C(n348), .Y(n2552) );
  OAI21X1 U1983 ( .A(n2040), .B(n2103), .C(n350), .Y(n2551) );
  OAI21X1 U1984 ( .A(n2040), .B(n2105), .C(n352), .Y(n2550) );
  OAI21X1 U1985 ( .A(n2040), .B(n276), .C(n354), .Y(n2549) );
  OAI21X1 U1986 ( .A(n2041), .B(n2079), .C(n356), .Y(n2548) );
  OAI21X1 U1987 ( .A(n2041), .B(n2081), .C(n358), .Y(n2547) );
  OAI21X1 U1988 ( .A(n2041), .B(n2083), .C(n360), .Y(n2546) );
  OAI21X1 U1989 ( .A(n2041), .B(n2085), .C(n362), .Y(n2545) );
  OAI21X1 U1990 ( .A(n2041), .B(n2087), .C(n364), .Y(n2544) );
  OAI21X1 U1991 ( .A(n2041), .B(n2089), .C(n366), .Y(n2543) );
  OAI21X1 U1992 ( .A(n2041), .B(n2091), .C(n368), .Y(n2542) );
  NAND2X1 U1993 ( .A(\mem<17><7> ), .B(n188), .Y(n2233) );
  OAI21X1 U1994 ( .A(n2041), .B(n1445), .C(n2233), .Y(n2541) );
  OAI21X1 U1995 ( .A(n2042), .B(n2093), .C(n370), .Y(n2540) );
  OAI21X1 U1996 ( .A(n2042), .B(n2095), .C(n372), .Y(n2539) );
  OAI21X1 U1997 ( .A(n2042), .B(n2097), .C(n374), .Y(n2538) );
  OAI21X1 U1998 ( .A(n2042), .B(n2099), .C(n376), .Y(n2537) );
  OAI21X1 U1999 ( .A(n2042), .B(n2101), .C(n378), .Y(n2536) );
  OAI21X1 U2000 ( .A(n2042), .B(n2103), .C(n380), .Y(n2535) );
  OAI21X1 U2001 ( .A(n2042), .B(n2105), .C(n382), .Y(n2534) );
  OAI21X1 U2002 ( .A(n2042), .B(n1463), .C(n384), .Y(n2533) );
  OAI21X1 U2003 ( .A(n2043), .B(n2079), .C(n386), .Y(n2532) );
  OAI21X1 U2004 ( .A(n2043), .B(n2081), .C(n388), .Y(n2531) );
  OAI21X1 U2005 ( .A(n2043), .B(n2083), .C(n390), .Y(n2530) );
  OAI21X1 U2006 ( .A(n2043), .B(n2085), .C(n392), .Y(n2529) );
  OAI21X1 U2007 ( .A(n2043), .B(n2087), .C(n394), .Y(n2528) );
  OAI21X1 U2008 ( .A(n2043), .B(n2089), .C(n396), .Y(n2527) );
  OAI21X1 U2009 ( .A(n2043), .B(n2091), .C(n398), .Y(n2526) );
  NAND2X1 U2010 ( .A(\mem<16><7> ), .B(n190), .Y(n2234) );
  OAI21X1 U2011 ( .A(n2043), .B(n1450), .C(n2234), .Y(n2525) );
  OAI21X1 U2012 ( .A(n2043), .B(n2093), .C(n400), .Y(n2524) );
  OAI21X1 U2013 ( .A(n2043), .B(n2095), .C(n402), .Y(n2523) );
  OAI21X1 U2014 ( .A(n2043), .B(n2097), .C(n404), .Y(n2522) );
  OAI21X1 U2015 ( .A(n2043), .B(n2099), .C(n406), .Y(n2521) );
  OAI21X1 U2016 ( .A(n2043), .B(n2101), .C(n408), .Y(n2520) );
  OAI21X1 U2017 ( .A(n2043), .B(n2103), .C(n410), .Y(n2519) );
  OAI21X1 U2018 ( .A(n2043), .B(n2105), .C(n412), .Y(n2518) );
  NAND2X1 U2019 ( .A(\mem<16><15> ), .B(n190), .Y(n2235) );
  OAI21X1 U2020 ( .A(n2043), .B(n1459), .C(n2235), .Y(n2517) );
  NAND3X1 U2021 ( .A(n2114), .B(n2773), .C(n2116), .Y(n2236) );
  OAI21X1 U2022 ( .A(n2044), .B(n2079), .C(n414), .Y(n2516) );
  OAI21X1 U2023 ( .A(n2044), .B(n2081), .C(n416), .Y(n2515) );
  OAI21X1 U2024 ( .A(n2044), .B(n2083), .C(n418), .Y(n2514) );
  OAI21X1 U2025 ( .A(n2044), .B(n2085), .C(n420), .Y(n2513) );
  OAI21X1 U2026 ( .A(n2044), .B(n2087), .C(n422), .Y(n2512) );
  OAI21X1 U2027 ( .A(n2044), .B(n2089), .C(n424), .Y(n2511) );
  OAI21X1 U2028 ( .A(n2044), .B(n2091), .C(n426), .Y(n2510) );
  NAND2X1 U2029 ( .A(\mem<15><7> ), .B(n192), .Y(n2237) );
  OAI21X1 U2030 ( .A(n2044), .B(n207), .C(n2237), .Y(n2509) );
  OAI21X1 U2031 ( .A(n2045), .B(n2093), .C(n428), .Y(n2508) );
  OAI21X1 U2032 ( .A(n2045), .B(n2095), .C(n430), .Y(n2507) );
  OAI21X1 U2033 ( .A(n2045), .B(n2097), .C(n432), .Y(n2506) );
  OAI21X1 U2034 ( .A(n2045), .B(n2099), .C(n434), .Y(n2505) );
  OAI21X1 U2035 ( .A(n2045), .B(n2101), .C(n436), .Y(n2504) );
  OAI21X1 U2036 ( .A(n2045), .B(n2103), .C(n438), .Y(n2503) );
  OAI21X1 U2037 ( .A(n2045), .B(n2105), .C(n440), .Y(n2502) );
  OAI21X1 U2038 ( .A(n2045), .B(n1458), .C(n239), .Y(n2501) );
  OAI21X1 U2039 ( .A(n2046), .B(n2079), .C(n442), .Y(n2500) );
  OAI21X1 U2040 ( .A(n2046), .B(n2081), .C(n444), .Y(n2499) );
  OAI21X1 U2041 ( .A(n2046), .B(n2083), .C(n446), .Y(n2498) );
  OAI21X1 U2042 ( .A(n2046), .B(n2085), .C(n448), .Y(n2497) );
  OAI21X1 U2043 ( .A(n2046), .B(n2087), .C(n450), .Y(n2496) );
  OAI21X1 U2044 ( .A(n2046), .B(n2089), .C(n452), .Y(n2495) );
  OAI21X1 U2045 ( .A(n2046), .B(n2091), .C(n454), .Y(n2494) );
  NAND2X1 U2046 ( .A(\mem<14><7> ), .B(n194), .Y(n2238) );
  OAI21X1 U2047 ( .A(n2046), .B(n1446), .C(n2238), .Y(n2493) );
  OAI21X1 U2048 ( .A(n2047), .B(n2093), .C(n456), .Y(n2492) );
  OAI21X1 U2049 ( .A(n2047), .B(n2095), .C(n458), .Y(n2491) );
  OAI21X1 U2050 ( .A(n2047), .B(n2097), .C(n460), .Y(n2490) );
  OAI21X1 U2051 ( .A(n2047), .B(n2099), .C(n462), .Y(n2489) );
  OAI21X1 U2052 ( .A(n2047), .B(n2101), .C(n464), .Y(n2488) );
  OAI21X1 U2053 ( .A(n2047), .B(n2103), .C(n466), .Y(n2487) );
  OAI21X1 U2054 ( .A(n2047), .B(n2105), .C(n468), .Y(n2486) );
  OAI21X1 U2055 ( .A(n2047), .B(n1459), .C(n241), .Y(n2485) );
  OAI21X1 U2056 ( .A(n2048), .B(n2079), .C(n470), .Y(n2484) );
  OAI21X1 U2057 ( .A(n2048), .B(n2081), .C(n472), .Y(n2483) );
  OAI21X1 U2058 ( .A(n2048), .B(n2083), .C(n474), .Y(n2482) );
  OAI21X1 U2059 ( .A(n2048), .B(n2085), .C(n476), .Y(n2481) );
  OAI21X1 U2060 ( .A(n2048), .B(n2087), .C(n478), .Y(n2480) );
  OAI21X1 U2061 ( .A(n2048), .B(n2089), .C(n480), .Y(n2479) );
  OAI21X1 U2062 ( .A(n2048), .B(n2091), .C(n482), .Y(n2478) );
  NAND2X1 U2063 ( .A(\mem<13><7> ), .B(n196), .Y(n2239) );
  OAI21X1 U2064 ( .A(n2048), .B(n1447), .C(n2239), .Y(n2477) );
  OAI21X1 U2065 ( .A(n2049), .B(n2093), .C(n484), .Y(n2476) );
  OAI21X1 U2066 ( .A(n2049), .B(n2095), .C(n486), .Y(n2475) );
  OAI21X1 U2067 ( .A(n2049), .B(n2097), .C(n488), .Y(n2474) );
  OAI21X1 U2068 ( .A(n2049), .B(n2099), .C(n490), .Y(n2473) );
  OAI21X1 U2069 ( .A(n2049), .B(n2101), .C(n492), .Y(n2472) );
  OAI21X1 U2070 ( .A(n2049), .B(n2103), .C(n494), .Y(n2471) );
  OAI21X1 U2071 ( .A(n2049), .B(n2105), .C(n496), .Y(n2470) );
  OAI21X1 U2072 ( .A(n2049), .B(n1460), .C(n243), .Y(n2469) );
  OAI21X1 U2073 ( .A(n2050), .B(n2079), .C(n498), .Y(n2468) );
  OAI21X1 U2074 ( .A(n2050), .B(n2081), .C(n500), .Y(n2467) );
  OAI21X1 U2075 ( .A(n2050), .B(n2083), .C(n502), .Y(n2466) );
  OAI21X1 U2076 ( .A(n2050), .B(n2085), .C(n504), .Y(n2465) );
  OAI21X1 U2077 ( .A(n2050), .B(n2087), .C(n506), .Y(n2464) );
  OAI21X1 U2078 ( .A(n2050), .B(n2089), .C(n508), .Y(n2463) );
  OAI21X1 U2079 ( .A(n2050), .B(n2091), .C(n510), .Y(n2462) );
  NAND2X1 U2080 ( .A(\mem<12><7> ), .B(n198), .Y(n2240) );
  OAI21X1 U2081 ( .A(n2050), .B(n1446), .C(n2240), .Y(n2461) );
  OAI21X1 U2082 ( .A(n2051), .B(n2093), .C(n512), .Y(n2460) );
  OAI21X1 U2083 ( .A(n2051), .B(n2095), .C(n514), .Y(n2459) );
  OAI21X1 U2084 ( .A(n2051), .B(n2097), .C(n516), .Y(n2458) );
  OAI21X1 U2085 ( .A(n2051), .B(n2099), .C(n518), .Y(n2457) );
  OAI21X1 U2086 ( .A(n2051), .B(n2101), .C(n520), .Y(n2456) );
  OAI21X1 U2087 ( .A(n2051), .B(n2103), .C(n522), .Y(n2455) );
  OAI21X1 U2088 ( .A(n2051), .B(n2105), .C(n524), .Y(n2454) );
  OAI21X1 U2089 ( .A(n2051), .B(n1465), .C(n245), .Y(n2453) );
  OAI21X1 U2090 ( .A(n2052), .B(n2079), .C(n526), .Y(n2452) );
  OAI21X1 U2091 ( .A(n2052), .B(n2080), .C(n528), .Y(n2451) );
  OAI21X1 U2092 ( .A(n2052), .B(n2082), .C(n530), .Y(n2450) );
  OAI21X1 U2093 ( .A(n2052), .B(n2084), .C(n532), .Y(n2449) );
  OAI21X1 U2094 ( .A(n2052), .B(n2086), .C(n534), .Y(n2448) );
  OAI21X1 U2095 ( .A(n2052), .B(n2088), .C(n536), .Y(n2447) );
  OAI21X1 U2096 ( .A(n2052), .B(n2090), .C(n538), .Y(n2446) );
  NAND2X1 U2097 ( .A(\mem<11><7> ), .B(n200), .Y(n2241) );
  OAI21X1 U2098 ( .A(n2052), .B(n1449), .C(n2241), .Y(n2445) );
  OAI21X1 U2099 ( .A(n2053), .B(n2092), .C(n540), .Y(n2444) );
  OAI21X1 U2100 ( .A(n2053), .B(n2094), .C(n542), .Y(n2443) );
  OAI21X1 U2101 ( .A(n2053), .B(n2096), .C(n544), .Y(n2442) );
  OAI21X1 U2102 ( .A(n2053), .B(n2098), .C(n546), .Y(n2441) );
  OAI21X1 U2103 ( .A(n2053), .B(n2100), .C(n548), .Y(n2440) );
  OAI21X1 U2104 ( .A(n2053), .B(n2102), .C(n550), .Y(n2439) );
  OAI21X1 U2105 ( .A(n2053), .B(n2104), .C(n552), .Y(n2438) );
  OAI21X1 U2106 ( .A(n2053), .B(n1462), .C(n247), .Y(n2437) );
  OAI21X1 U2107 ( .A(n2054), .B(n2079), .C(n554), .Y(n2436) );
  OAI21X1 U2108 ( .A(n2054), .B(n2080), .C(n556), .Y(n2435) );
  OAI21X1 U2109 ( .A(n2054), .B(n2082), .C(n558), .Y(n2434) );
  OAI21X1 U2110 ( .A(n2054), .B(n2084), .C(n560), .Y(n2433) );
  OAI21X1 U2111 ( .A(n2054), .B(n2086), .C(n562), .Y(n2432) );
  OAI21X1 U2112 ( .A(n2054), .B(n2088), .C(n564), .Y(n2431) );
  OAI21X1 U2113 ( .A(n2054), .B(n2090), .C(n566), .Y(n2430) );
  NAND2X1 U2114 ( .A(\mem<10><7> ), .B(n202), .Y(n2242) );
  OAI21X1 U2115 ( .A(n2054), .B(n207), .C(n2242), .Y(n2429) );
  OAI21X1 U2116 ( .A(n2055), .B(n2092), .C(n568), .Y(n2428) );
  OAI21X1 U2117 ( .A(n2055), .B(n2094), .C(n570), .Y(n2427) );
  OAI21X1 U2118 ( .A(n2055), .B(n2096), .C(n572), .Y(n2426) );
  OAI21X1 U2119 ( .A(n2055), .B(n2098), .C(n574), .Y(n2425) );
  OAI21X1 U2120 ( .A(n2055), .B(n2100), .C(n576), .Y(n2424) );
  OAI21X1 U2121 ( .A(n2055), .B(n2102), .C(n578), .Y(n2423) );
  OAI21X1 U2122 ( .A(n2055), .B(n2104), .C(n580), .Y(n2422) );
  OAI21X1 U2123 ( .A(n2055), .B(n1451), .C(n249), .Y(n2421) );
  OAI21X1 U2124 ( .A(n2056), .B(n2079), .C(n582), .Y(n2420) );
  OAI21X1 U2125 ( .A(n2056), .B(n2080), .C(n584), .Y(n2419) );
  OAI21X1 U2126 ( .A(n2056), .B(n2082), .C(n586), .Y(n2418) );
  OAI21X1 U2127 ( .A(n2056), .B(n2084), .C(n588), .Y(n2417) );
  OAI21X1 U2128 ( .A(n2056), .B(n2086), .C(n590), .Y(n2416) );
  OAI21X1 U2129 ( .A(n2056), .B(n2088), .C(n592), .Y(n2415) );
  OAI21X1 U2130 ( .A(n2056), .B(n2090), .C(n594), .Y(n2414) );
  NAND2X1 U2131 ( .A(\mem<9><7> ), .B(n204), .Y(n2243) );
  OAI21X1 U2132 ( .A(n2056), .B(n1448), .C(n2243), .Y(n2413) );
  OAI21X1 U2133 ( .A(n2057), .B(n2092), .C(n596), .Y(n2412) );
  OAI21X1 U2134 ( .A(n2057), .B(n2094), .C(n598), .Y(n2411) );
  OAI21X1 U2135 ( .A(n2057), .B(n2096), .C(n600), .Y(n2410) );
  OAI21X1 U2136 ( .A(n2057), .B(n2098), .C(n602), .Y(n2409) );
  OAI21X1 U2137 ( .A(n2057), .B(n2100), .C(n604), .Y(n2408) );
  OAI21X1 U2138 ( .A(n2057), .B(n2102), .C(n606), .Y(n2407) );
  OAI21X1 U2139 ( .A(n2057), .B(n2104), .C(n608), .Y(n2406) );
  OAI21X1 U2140 ( .A(n2057), .B(n1463), .C(n251), .Y(n2405) );
  OAI21X1 U2141 ( .A(n2058), .B(n2079), .C(n610), .Y(n2404) );
  OAI21X1 U2142 ( .A(n2058), .B(n2080), .C(n612), .Y(n2403) );
  OAI21X1 U2143 ( .A(n2058), .B(n2082), .C(n614), .Y(n2402) );
  OAI21X1 U2144 ( .A(n2058), .B(n2084), .C(n616), .Y(n2401) );
  OAI21X1 U2145 ( .A(n2058), .B(n2086), .C(n618), .Y(n2400) );
  OAI21X1 U2146 ( .A(n2058), .B(n2088), .C(n620), .Y(n2399) );
  OAI21X1 U2147 ( .A(n2058), .B(n2090), .C(n622), .Y(n2398) );
  OAI21X1 U2148 ( .A(n2058), .B(n1445), .C(n253), .Y(n2397) );
  OAI21X1 U2149 ( .A(n2058), .B(n2092), .C(n624), .Y(n2396) );
  OAI21X1 U2150 ( .A(n2058), .B(n2094), .C(n626), .Y(n2395) );
  OAI21X1 U2151 ( .A(n2058), .B(n2096), .C(n628), .Y(n2394) );
  OAI21X1 U2152 ( .A(n2058), .B(n2098), .C(n630), .Y(n2393) );
  OAI21X1 U2153 ( .A(n2058), .B(n2100), .C(n632), .Y(n2392) );
  OAI21X1 U2154 ( .A(n2058), .B(n2102), .C(n634), .Y(n2391) );
  OAI21X1 U2155 ( .A(n2058), .B(n2104), .C(n636), .Y(n2390) );
  OAI21X1 U2156 ( .A(n2058), .B(n1460), .C(n255), .Y(n2389) );
  NAND3X1 U2157 ( .A(n2115), .B(n2773), .C(n2116), .Y(n2245) );
  OAI21X1 U2158 ( .A(n2059), .B(n2078), .C(n638), .Y(n2388) );
  OAI21X1 U2159 ( .A(n2059), .B(n2080), .C(n640), .Y(n2387) );
  OAI21X1 U2160 ( .A(n2059), .B(n2082), .C(n642), .Y(n2386) );
  OAI21X1 U2161 ( .A(n2059), .B(n2084), .C(n644), .Y(n2385) );
  OAI21X1 U2162 ( .A(n2059), .B(n2086), .C(n646), .Y(n2384) );
  OAI21X1 U2163 ( .A(n2059), .B(n2088), .C(n648), .Y(n2383) );
  OAI21X1 U2164 ( .A(n2059), .B(n2090), .C(n650), .Y(n2382) );
  OAI21X1 U2165 ( .A(n2059), .B(n1449), .C(n170), .Y(n2381) );
  OAI21X1 U2166 ( .A(n2060), .B(n2092), .C(n1164), .Y(n2380) );
  OAI21X1 U2167 ( .A(n2060), .B(n2094), .C(n1166), .Y(n2379) );
  OAI21X1 U2168 ( .A(n2060), .B(n2096), .C(n1168), .Y(n2378) );
  OAI21X1 U2169 ( .A(n2060), .B(n2098), .C(n1170), .Y(n2377) );
  OAI21X1 U2170 ( .A(n2060), .B(n2100), .C(n1172), .Y(n2376) );
  OAI21X1 U2171 ( .A(n2060), .B(n2102), .C(n1174), .Y(n2375) );
  OAI21X1 U2172 ( .A(n2060), .B(n2104), .C(n1176), .Y(n2374) );
  NAND2X1 U2173 ( .A(\mem<7><15> ), .B(n259), .Y(n2246) );
  OAI21X1 U2174 ( .A(n2060), .B(n1452), .C(n2246), .Y(n2373) );
  OAI21X1 U2175 ( .A(n2061), .B(n2079), .C(n1178), .Y(n2372) );
  OAI21X1 U2176 ( .A(n2061), .B(n2080), .C(n1180), .Y(n2371) );
  OAI21X1 U2177 ( .A(n2061), .B(n2082), .C(n1182), .Y(n2370) );
  OAI21X1 U2178 ( .A(n2061), .B(n2084), .C(n1184), .Y(n2369) );
  OAI21X1 U2179 ( .A(n2061), .B(n2086), .C(n1186), .Y(n2368) );
  OAI21X1 U2180 ( .A(n2061), .B(n2088), .C(n1188), .Y(n2367) );
  OAI21X1 U2181 ( .A(n2061), .B(n2090), .C(n1190), .Y(n2366) );
  OAI21X1 U2182 ( .A(n2061), .B(n1450), .C(n172), .Y(n2365) );
  OAI21X1 U2183 ( .A(n2062), .B(n2092), .C(n1192), .Y(n2364) );
  OAI21X1 U2184 ( .A(n2062), .B(n2094), .C(n1194), .Y(n2363) );
  OAI21X1 U2185 ( .A(n2062), .B(n2096), .C(n1196), .Y(n2362) );
  OAI21X1 U2186 ( .A(n2062), .B(n2098), .C(n1198), .Y(n2361) );
  OAI21X1 U2187 ( .A(n2062), .B(n2100), .C(n1200), .Y(n2360) );
  OAI21X1 U2188 ( .A(n2062), .B(n2102), .C(n1202), .Y(n2359) );
  OAI21X1 U2189 ( .A(n2062), .B(n2104), .C(n1204), .Y(n2358) );
  NAND2X1 U2190 ( .A(\mem<6><15> ), .B(n261), .Y(n2247) );
  OAI21X1 U2191 ( .A(n2062), .B(n1453), .C(n2247), .Y(n2357) );
  OAI21X1 U2192 ( .A(n2063), .B(n2078), .C(n1206), .Y(n2356) );
  OAI21X1 U2193 ( .A(n2063), .B(n2080), .C(n1208), .Y(n2355) );
  OAI21X1 U2194 ( .A(n2063), .B(n2082), .C(n1210), .Y(n2354) );
  OAI21X1 U2195 ( .A(n2063), .B(n2084), .C(n1212), .Y(n2353) );
  OAI21X1 U2196 ( .A(n2063), .B(n2086), .C(n1214), .Y(n2352) );
  OAI21X1 U2197 ( .A(n2063), .B(n2088), .C(n1216), .Y(n2351) );
  OAI21X1 U2198 ( .A(n2063), .B(n2090), .C(n1218), .Y(n2350) );
  OAI21X1 U2199 ( .A(n2063), .B(n1450), .C(n174), .Y(n2349) );
  OAI21X1 U2200 ( .A(n2064), .B(n2092), .C(n1220), .Y(n2348) );
  OAI21X1 U2201 ( .A(n2064), .B(n2094), .C(n1222), .Y(n2347) );
  OAI21X1 U2202 ( .A(n2064), .B(n2096), .C(n1224), .Y(n2346) );
  OAI21X1 U2203 ( .A(n2064), .B(n2098), .C(n1226), .Y(n2345) );
  OAI21X1 U2204 ( .A(n2064), .B(n2100), .C(n1228), .Y(n2344) );
  OAI21X1 U2205 ( .A(n2064), .B(n2102), .C(n1230), .Y(n2343) );
  OAI21X1 U2206 ( .A(n2064), .B(n2104), .C(n1232), .Y(n2342) );
  NAND2X1 U2207 ( .A(\mem<5><15> ), .B(n263), .Y(n2249) );
  OAI21X1 U2208 ( .A(n2064), .B(n1453), .C(n2249), .Y(n2341) );
  OAI21X1 U2209 ( .A(n2065), .B(n2079), .C(n1234), .Y(n2340) );
  OAI21X1 U2210 ( .A(n2065), .B(n2080), .C(n1236), .Y(n2339) );
  OAI21X1 U2211 ( .A(n2065), .B(n2082), .C(n1238), .Y(n2338) );
  OAI21X1 U2212 ( .A(n2065), .B(n2084), .C(n1240), .Y(n2337) );
  OAI21X1 U2213 ( .A(n2065), .B(n2086), .C(n1242), .Y(n2336) );
  OAI21X1 U2214 ( .A(n2065), .B(n2088), .C(n1244), .Y(n2335) );
  OAI21X1 U2215 ( .A(n2065), .B(n2090), .C(n1246), .Y(n2334) );
  OAI21X1 U2216 ( .A(n2065), .B(n275), .C(n176), .Y(n2333) );
  OAI21X1 U2217 ( .A(n2066), .B(n2092), .C(n1248), .Y(n2332) );
  OAI21X1 U2218 ( .A(n2066), .B(n2094), .C(n1250), .Y(n2331) );
  OAI21X1 U2219 ( .A(n2066), .B(n2096), .C(n1252), .Y(n2330) );
  OAI21X1 U2220 ( .A(n2066), .B(n2098), .C(n1254), .Y(n2329) );
  OAI21X1 U2221 ( .A(n2066), .B(n2100), .C(n1256), .Y(n2328) );
  OAI21X1 U2222 ( .A(n2066), .B(n2102), .C(n1258), .Y(n2327) );
  OAI21X1 U2223 ( .A(n2066), .B(n2104), .C(n1260), .Y(n2326) );
  OAI21X1 U2224 ( .A(n2066), .B(n1454), .C(n294), .Y(n2325) );
  OAI21X1 U2225 ( .A(n2067), .B(n2078), .C(n1262), .Y(n2324) );
  OAI21X1 U2226 ( .A(n2067), .B(n2080), .C(n1264), .Y(n2323) );
  OAI21X1 U2227 ( .A(n2067), .B(n2082), .C(n1266), .Y(n2322) );
  OAI21X1 U2228 ( .A(n2067), .B(n2084), .C(n1268), .Y(n2321) );
  OAI21X1 U2229 ( .A(n2067), .B(n2086), .C(n1270), .Y(n2320) );
  OAI21X1 U2230 ( .A(n2067), .B(n2088), .C(n1272), .Y(n2319) );
  OAI21X1 U2231 ( .A(n2067), .B(n2090), .C(n1274), .Y(n2318) );
  OAI21X1 U2232 ( .A(n2067), .B(n207), .C(n178), .Y(n2317) );
  OAI21X1 U2233 ( .A(n2068), .B(n2092), .C(n1276), .Y(n2316) );
  OAI21X1 U2234 ( .A(n2068), .B(n2094), .C(n1278), .Y(n2315) );
  OAI21X1 U2235 ( .A(n2068), .B(n2096), .C(n1280), .Y(n2314) );
  OAI21X1 U2236 ( .A(n2068), .B(n2098), .C(n1282), .Y(n2313) );
  OAI21X1 U2237 ( .A(n2068), .B(n2100), .C(n1284), .Y(n2312) );
  OAI21X1 U2238 ( .A(n2068), .B(n2102), .C(n1286), .Y(n2311) );
  OAI21X1 U2239 ( .A(n2068), .B(n2104), .C(n1288), .Y(n2310) );
  NAND2X1 U2240 ( .A(\mem<3><15> ), .B(n267), .Y(n2252) );
  OAI21X1 U2241 ( .A(n2068), .B(n1466), .C(n2252), .Y(n2309) );
  OAI21X1 U2242 ( .A(n2069), .B(n2079), .C(n1290), .Y(n2308) );
  OAI21X1 U2243 ( .A(n2069), .B(n2080), .C(n1292), .Y(n2307) );
  OAI21X1 U2244 ( .A(n2069), .B(n2082), .C(n1294), .Y(n2306) );
  OAI21X1 U2245 ( .A(n2069), .B(n2084), .C(n1296), .Y(n2305) );
  OAI21X1 U2246 ( .A(n2069), .B(n2086), .C(n1298), .Y(n2304) );
  OAI21X1 U2247 ( .A(n2069), .B(n2088), .C(n1300), .Y(n2303) );
  OAI21X1 U2248 ( .A(n2069), .B(n2090), .C(n1302), .Y(n2302) );
  OAI21X1 U2249 ( .A(n2069), .B(n1445), .C(n180), .Y(n2301) );
  OAI21X1 U2250 ( .A(n2070), .B(n2092), .C(n1304), .Y(n2300) );
  OAI21X1 U2251 ( .A(n2070), .B(n2094), .C(n1306), .Y(n2299) );
  OAI21X1 U2252 ( .A(n2070), .B(n2096), .C(n1308), .Y(n2298) );
  OAI21X1 U2253 ( .A(n2070), .B(n2098), .C(n1310), .Y(n2297) );
  OAI21X1 U2254 ( .A(n2070), .B(n2100), .C(n1312), .Y(n2296) );
  OAI21X1 U2255 ( .A(n2070), .B(n2102), .C(n1314), .Y(n2295) );
  OAI21X1 U2256 ( .A(n2070), .B(n2104), .C(n1316), .Y(n2294) );
  NAND2X1 U2257 ( .A(\mem<2><15> ), .B(n269), .Y(n2254) );
  OAI21X1 U2258 ( .A(n2070), .B(n1457), .C(n2254), .Y(n2293) );
  OAI21X1 U2259 ( .A(n2071), .B(n2079), .C(n1318), .Y(n2292) );
  OAI21X1 U2260 ( .A(n2071), .B(n2080), .C(n1320), .Y(n2291) );
  OAI21X1 U2261 ( .A(n2071), .B(n2082), .C(n1322), .Y(n2290) );
  OAI21X1 U2262 ( .A(n2071), .B(n2084), .C(n1324), .Y(n2289) );
  OAI21X1 U2263 ( .A(n2071), .B(n2086), .C(n1326), .Y(n2288) );
  OAI21X1 U2264 ( .A(n2071), .B(n2088), .C(n1328), .Y(n2287) );
  OAI21X1 U2265 ( .A(n2071), .B(n2090), .C(n1330), .Y(n2286) );
  OAI21X1 U2266 ( .A(n2071), .B(n1447), .C(n182), .Y(n2285) );
  OAI21X1 U2267 ( .A(n2072), .B(n2092), .C(n1332), .Y(n2284) );
  OAI21X1 U2268 ( .A(n2072), .B(n2094), .C(n1334), .Y(n2283) );
  OAI21X1 U2269 ( .A(n2072), .B(n2096), .C(n1336), .Y(n2282) );
  OAI21X1 U2270 ( .A(n2072), .B(n2098), .C(n1338), .Y(n2281) );
  OAI21X1 U2271 ( .A(n2072), .B(n2100), .C(n1340), .Y(n2280) );
  OAI21X1 U2272 ( .A(n2072), .B(n2102), .C(n1342), .Y(n2279) );
  OAI21X1 U2273 ( .A(n2072), .B(n2104), .C(n1344), .Y(n2278) );
  NAND2X1 U2274 ( .A(\mem<1><15> ), .B(n271), .Y(n2256) );
  OAI21X1 U2275 ( .A(n2072), .B(n1458), .C(n2256), .Y(n2277) );
  OAI21X1 U2276 ( .A(n2073), .B(n2078), .C(n1346), .Y(n2276) );
  OAI21X1 U2277 ( .A(n2073), .B(n2080), .C(n1348), .Y(n2275) );
  OAI21X1 U2278 ( .A(n2073), .B(n2082), .C(n1350), .Y(n2274) );
  OAI21X1 U2279 ( .A(n2073), .B(n2084), .C(n1352), .Y(n2273) );
  OAI21X1 U2280 ( .A(n2073), .B(n2086), .C(n1354), .Y(n2272) );
  OAI21X1 U2281 ( .A(n2073), .B(n2088), .C(n1356), .Y(n2271) );
  OAI21X1 U2282 ( .A(n2073), .B(n2090), .C(n1358), .Y(n2270) );
  NAND2X1 U2283 ( .A(\mem<0><7> ), .B(n206), .Y(n2259) );
  OAI21X1 U2284 ( .A(n2073), .B(n275), .C(n2259), .Y(n2269) );
  OAI21X1 U2285 ( .A(n2073), .B(n2092), .C(n1360), .Y(n2268) );
  OAI21X1 U2286 ( .A(n2073), .B(n2094), .C(n1362), .Y(n2267) );
  OAI21X1 U2287 ( .A(n2073), .B(n2096), .C(n1364), .Y(n2266) );
  OAI21X1 U2288 ( .A(n2073), .B(n2098), .C(n1366), .Y(n2265) );
  OAI21X1 U2289 ( .A(n2073), .B(n2100), .C(n1368), .Y(n2264) );
  OAI21X1 U2290 ( .A(n2073), .B(n2102), .C(n1370), .Y(n2263) );
  OAI21X1 U2291 ( .A(n2073), .B(n2104), .C(n1372), .Y(n2262) );
  NAND2X1 U2292 ( .A(\mem<0><15> ), .B(n206), .Y(n2260) );
  OAI21X1 U2293 ( .A(n2073), .B(n1466), .C(n2260), .Y(n2261) );
endmodule


module memc_Size5_0 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , N17, N18, N19, N20, N21, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n58, n59, n60, n61, n62, n63,
         n64, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79,
         n80, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n106, n107, n108, n109,
         n110, n111, n112, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n287, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n847), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n848), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n849), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n850), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n851), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n852), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n853), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n854), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n855), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n856), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n857), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n858), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n859), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n860), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n861), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n862), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n863), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n864), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n865), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n866), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n867), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n868), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n869), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n870), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n871), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n872), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n873), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n874), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n875), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n876), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n877), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n878), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n879), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n880), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n881), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n882), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n883), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n884), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n885), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n886), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n887), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n888), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n889), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n890), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n891), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n892), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n893), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n894), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n895), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n896), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n897), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n898), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n899), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n900), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n901), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n902), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n903), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n904), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n905), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n906), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n907), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n908), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n909), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n910), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n911), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n912), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n913), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n914), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n915), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n916), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n917), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n918), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n919), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n920), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n921), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n922), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n923), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n924), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n925), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n926), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n927), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n928), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n929), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n930), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n931), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n932), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n933), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n934), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n935), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n936), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n937), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n938), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n939), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n940), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n941), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n942), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n943), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n944), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n945), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n946), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n947), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n948), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n949), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n950), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n951), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n952), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n953), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n954), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n955), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n956), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n957), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n958), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n959), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n960), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n961), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n962), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n963), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n964), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n965), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n966), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n967), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n968), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n969), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n970), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n971), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n972), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n973), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n974), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n975), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n976), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n977), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n978), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n979), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n980), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n981), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n982), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n983), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n984), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n985), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n986), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n987), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n988), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n989), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n990), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n991), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n992), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n993), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n994), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n995), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n996), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n997), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n998), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n999), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1000), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1001), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1002), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1003), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1004), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1005), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1006), .CLK(clk), .Q(\mem<31><0> ) );
  OAI21X1 U50 ( .A(n579), .B(n831), .C(n497), .Y(n1006) );
  OAI21X1 U52 ( .A(n579), .B(n829), .C(n495), .Y(n1005) );
  OAI21X1 U54 ( .A(n579), .B(n827), .C(n493), .Y(n1004) );
  OAI21X1 U56 ( .A(n579), .B(n825), .C(n491), .Y(n1003) );
  OAI21X1 U58 ( .A(n579), .B(n823), .C(n489), .Y(n1002) );
  OAI21X1 U62 ( .A(n831), .B(n642), .C(n487), .Y(n1001) );
  OAI21X1 U64 ( .A(n829), .B(n642), .C(n485), .Y(n1000) );
  OAI21X1 U66 ( .A(n827), .B(n642), .C(n483), .Y(n999) );
  OAI21X1 U68 ( .A(n825), .B(n642), .C(n481), .Y(n998) );
  OAI21X1 U70 ( .A(n823), .B(n642), .C(n479), .Y(n997) );
  OAI21X1 U74 ( .A(n831), .B(n640), .C(n477), .Y(n996) );
  OAI21X1 U76 ( .A(n829), .B(n640), .C(n475), .Y(n995) );
  OAI21X1 U78 ( .A(n827), .B(n640), .C(n473), .Y(n994) );
  OAI21X1 U80 ( .A(n825), .B(n640), .C(n471), .Y(n993) );
  OAI21X1 U82 ( .A(n823), .B(n640), .C(n469), .Y(n992) );
  OAI21X1 U86 ( .A(n831), .B(n638), .C(n467), .Y(n991) );
  OAI21X1 U88 ( .A(n829), .B(n638), .C(n465), .Y(n990) );
  OAI21X1 U90 ( .A(n827), .B(n638), .C(n463), .Y(n989) );
  OAI21X1 U92 ( .A(n825), .B(n638), .C(n461), .Y(n988) );
  OAI21X1 U94 ( .A(n823), .B(n638), .C(n459), .Y(n987) );
  OAI21X1 U98 ( .A(n831), .B(n636), .C(n457), .Y(n986) );
  OAI21X1 U100 ( .A(n829), .B(n636), .C(n455), .Y(n985) );
  OAI21X1 U102 ( .A(n827), .B(n636), .C(n453), .Y(n984) );
  OAI21X1 U104 ( .A(n825), .B(n636), .C(n451), .Y(n983) );
  OAI21X1 U106 ( .A(n823), .B(n636), .C(n449), .Y(n982) );
  OAI21X1 U110 ( .A(n831), .B(n634), .C(n287), .Y(n981) );
  OAI21X1 U112 ( .A(n829), .B(n634), .C(n284), .Y(n980) );
  OAI21X1 U114 ( .A(n827), .B(n634), .C(n282), .Y(n979) );
  OAI21X1 U116 ( .A(n825), .B(n634), .C(n280), .Y(n978) );
  OAI21X1 U118 ( .A(n823), .B(n634), .C(n278), .Y(n977) );
  OAI21X1 U122 ( .A(n831), .B(n632), .C(n276), .Y(n976) );
  OAI21X1 U124 ( .A(n829), .B(n632), .C(n274), .Y(n975) );
  OAI21X1 U126 ( .A(n827), .B(n632), .C(n272), .Y(n974) );
  OAI21X1 U128 ( .A(n825), .B(n632), .C(n270), .Y(n973) );
  OAI21X1 U130 ( .A(n823), .B(n632), .C(n268), .Y(n972) );
  OAI21X1 U134 ( .A(n831), .B(n630), .C(n266), .Y(n971) );
  OAI21X1 U136 ( .A(n829), .B(n630), .C(n264), .Y(n970) );
  OAI21X1 U138 ( .A(n827), .B(n630), .C(n262), .Y(n969) );
  OAI21X1 U140 ( .A(n825), .B(n630), .C(n260), .Y(n968) );
  OAI21X1 U142 ( .A(n823), .B(n630), .C(n258), .Y(n967) );
  NAND3X1 U146 ( .A(N13), .B(n1010), .C(n841), .Y(n1011) );
  OAI21X1 U147 ( .A(n831), .B(n628), .C(n256), .Y(n966) );
  OAI21X1 U149 ( .A(n829), .B(n628), .C(n254), .Y(n965) );
  OAI21X1 U151 ( .A(n827), .B(n628), .C(n252), .Y(n964) );
  OAI21X1 U153 ( .A(n825), .B(n628), .C(n250), .Y(n963) );
  OAI21X1 U155 ( .A(n823), .B(n628), .C(n248), .Y(n962) );
  OAI21X1 U159 ( .A(n831), .B(n625), .C(n246), .Y(n961) );
  OAI21X1 U161 ( .A(n829), .B(n625), .C(n244), .Y(n960) );
  OAI21X1 U163 ( .A(n827), .B(n625), .C(n242), .Y(n959) );
  OAI21X1 U165 ( .A(n825), .B(n625), .C(n240), .Y(n958) );
  OAI21X1 U167 ( .A(n823), .B(n625), .C(n238), .Y(n957) );
  OAI21X1 U171 ( .A(n831), .B(n624), .C(n236), .Y(n956) );
  OAI21X1 U173 ( .A(n829), .B(n624), .C(n234), .Y(n955) );
  OAI21X1 U175 ( .A(n827), .B(n624), .C(n232), .Y(n954) );
  OAI21X1 U177 ( .A(n825), .B(n624), .C(n230), .Y(n953) );
  OAI21X1 U179 ( .A(n823), .B(n624), .C(n227), .Y(n952) );
  OAI21X1 U183 ( .A(n831), .B(n621), .C(n225), .Y(n951) );
  OAI21X1 U185 ( .A(n829), .B(n621), .C(n223), .Y(n950) );
  OAI21X1 U187 ( .A(n827), .B(n621), .C(n221), .Y(n949) );
  OAI21X1 U189 ( .A(n825), .B(n621), .C(n219), .Y(n948) );
  OAI21X1 U191 ( .A(n823), .B(n621), .C(n217), .Y(n947) );
  OAI21X1 U195 ( .A(n831), .B(n620), .C(n215), .Y(n946) );
  OAI21X1 U197 ( .A(n829), .B(n620), .C(n213), .Y(n945) );
  OAI21X1 U199 ( .A(n827), .B(n620), .C(n211), .Y(n944) );
  OAI21X1 U201 ( .A(n825), .B(n620), .C(n209), .Y(n943) );
  OAI21X1 U203 ( .A(n823), .B(n620), .C(n207), .Y(n942) );
  OAI21X1 U207 ( .A(n832), .B(n617), .C(n205), .Y(n941) );
  OAI21X1 U209 ( .A(n830), .B(n617), .C(n203), .Y(n940) );
  OAI21X1 U211 ( .A(n828), .B(n617), .C(n201), .Y(n939) );
  OAI21X1 U213 ( .A(n826), .B(n617), .C(n199), .Y(n938) );
  OAI21X1 U215 ( .A(n824), .B(n617), .C(n197), .Y(n937) );
  OAI21X1 U219 ( .A(n832), .B(n616), .C(n195), .Y(n936) );
  OAI21X1 U221 ( .A(n830), .B(n616), .C(n193), .Y(n935) );
  OAI21X1 U223 ( .A(n828), .B(n616), .C(n191), .Y(n934) );
  OAI21X1 U225 ( .A(n826), .B(n616), .C(n189), .Y(n933) );
  OAI21X1 U227 ( .A(n824), .B(n616), .C(n187), .Y(n932) );
  OAI21X1 U231 ( .A(n832), .B(n614), .C(n185), .Y(n931) );
  OAI21X1 U233 ( .A(n830), .B(n614), .C(n183), .Y(n930) );
  OAI21X1 U235 ( .A(n828), .B(n614), .C(n181), .Y(n929) );
  OAI21X1 U237 ( .A(n826), .B(n614), .C(n179), .Y(n928) );
  OAI21X1 U239 ( .A(n824), .B(n614), .C(n177), .Y(n927) );
  NAND3X1 U243 ( .A(n1010), .B(n840), .C(n841), .Y(n1009) );
  OAI21X1 U244 ( .A(n832), .B(n612), .C(n175), .Y(n926) );
  OAI21X1 U246 ( .A(n830), .B(n612), .C(n173), .Y(n925) );
  OAI21X1 U248 ( .A(n828), .B(n612), .C(n170), .Y(n924) );
  OAI21X1 U250 ( .A(n826), .B(n612), .C(n168), .Y(n923) );
  OAI21X1 U252 ( .A(n824), .B(n612), .C(n166), .Y(n922) );
  OAI21X1 U256 ( .A(n832), .B(n610), .C(n164), .Y(n921) );
  OAI21X1 U258 ( .A(n830), .B(n610), .C(n162), .Y(n920) );
  OAI21X1 U260 ( .A(n828), .B(n610), .C(n160), .Y(n919) );
  OAI21X1 U262 ( .A(n826), .B(n610), .C(n158), .Y(n918) );
  OAI21X1 U264 ( .A(n824), .B(n610), .C(n156), .Y(n917) );
  OAI21X1 U268 ( .A(n832), .B(n608), .C(n154), .Y(n916) );
  OAI21X1 U270 ( .A(n830), .B(n608), .C(n152), .Y(n915) );
  OAI21X1 U272 ( .A(n828), .B(n608), .C(n150), .Y(n914) );
  OAI21X1 U274 ( .A(n826), .B(n608), .C(n148), .Y(n913) );
  OAI21X1 U276 ( .A(n824), .B(n608), .C(n146), .Y(n912) );
  OAI21X1 U280 ( .A(n832), .B(n606), .C(n144), .Y(n911) );
  OAI21X1 U282 ( .A(n830), .B(n606), .C(n142), .Y(n910) );
  OAI21X1 U284 ( .A(n828), .B(n606), .C(n140), .Y(n909) );
  OAI21X1 U286 ( .A(n826), .B(n606), .C(n138), .Y(n908) );
  OAI21X1 U288 ( .A(n824), .B(n606), .C(n136), .Y(n907) );
  OAI21X1 U292 ( .A(n832), .B(n604), .C(n134), .Y(n906) );
  OAI21X1 U294 ( .A(n830), .B(n604), .C(n132), .Y(n905) );
  OAI21X1 U296 ( .A(n828), .B(n604), .C(n130), .Y(n904) );
  OAI21X1 U298 ( .A(n826), .B(n604), .C(n128), .Y(n903) );
  OAI21X1 U300 ( .A(n824), .B(n604), .C(n126), .Y(n902) );
  OAI21X1 U304 ( .A(n832), .B(n602), .C(n124), .Y(n901) );
  OAI21X1 U306 ( .A(n830), .B(n602), .C(n122), .Y(n900) );
  OAI21X1 U308 ( .A(n828), .B(n602), .C(n120), .Y(n899) );
  OAI21X1 U310 ( .A(n826), .B(n602), .C(n118), .Y(n898) );
  OAI21X1 U312 ( .A(n824), .B(n602), .C(n116), .Y(n897) );
  OAI21X1 U316 ( .A(n832), .B(n600), .C(n111), .Y(n896) );
  OAI21X1 U318 ( .A(n830), .B(n600), .C(n109), .Y(n895) );
  OAI21X1 U320 ( .A(n828), .B(n600), .C(n107), .Y(n894) );
  OAI21X1 U322 ( .A(n826), .B(n600), .C(n104), .Y(n893) );
  OAI21X1 U324 ( .A(n824), .B(n600), .C(n102), .Y(n892) );
  OAI21X1 U328 ( .A(n832), .B(n598), .C(n100), .Y(n891) );
  OAI21X1 U330 ( .A(n830), .B(n598), .C(n98), .Y(n890) );
  OAI21X1 U332 ( .A(n828), .B(n598), .C(n95), .Y(n889) );
  OAI21X1 U334 ( .A(n826), .B(n598), .C(n93), .Y(n888) );
  OAI21X1 U336 ( .A(n824), .B(n598), .C(n91), .Y(n887) );
  NAND3X1 U340 ( .A(n1010), .B(n842), .C(N13), .Y(n1008) );
  OAI21X1 U341 ( .A(n832), .B(n596), .C(n88), .Y(n886) );
  OAI21X1 U343 ( .A(n830), .B(n596), .C(n86), .Y(n885) );
  OAI21X1 U345 ( .A(n828), .B(n596), .C(n84), .Y(n884) );
  OAI21X1 U347 ( .A(n826), .B(n596), .C(n82), .Y(n883) );
  OAI21X1 U349 ( .A(n824), .B(n596), .C(n79), .Y(n882) );
  NOR3X1 U353 ( .A(n837), .B(n822), .C(n839), .Y(n1019) );
  OAI21X1 U354 ( .A(n832), .B(n594), .C(n77), .Y(n881) );
  OAI21X1 U356 ( .A(n830), .B(n594), .C(n75), .Y(n880) );
  OAI21X1 U358 ( .A(n828), .B(n594), .C(n72), .Y(n879) );
  OAI21X1 U360 ( .A(n826), .B(n594), .C(n70), .Y(n878) );
  OAI21X1 U362 ( .A(n824), .B(n594), .C(n68), .Y(n877) );
  NOR3X1 U366 ( .A(n837), .B(n821), .C(n839), .Y(n1018) );
  OAI21X1 U367 ( .A(n831), .B(n592), .C(n66), .Y(n876) );
  OAI21X1 U369 ( .A(n829), .B(n592), .C(n63), .Y(n875) );
  OAI21X1 U371 ( .A(n827), .B(n592), .C(n61), .Y(n874) );
  OAI21X1 U373 ( .A(n825), .B(n592), .C(n59), .Y(n873) );
  OAI21X1 U375 ( .A(n823), .B(n592), .C(n55), .Y(n872) );
  NOR3X1 U379 ( .A(n822), .B(n836), .C(n839), .Y(n1017) );
  OAI21X1 U380 ( .A(n832), .B(n590), .C(n53), .Y(n871) );
  OAI21X1 U382 ( .A(n830), .B(n590), .C(n51), .Y(n870) );
  OAI21X1 U384 ( .A(n828), .B(n590), .C(n49), .Y(n869) );
  OAI21X1 U386 ( .A(n826), .B(n590), .C(n47), .Y(n868) );
  OAI21X1 U388 ( .A(n824), .B(n590), .C(n45), .Y(n867) );
  NOR3X1 U392 ( .A(n821), .B(n836), .C(n839), .Y(n1016) );
  OAI21X1 U393 ( .A(n831), .B(n588), .C(n43), .Y(n866) );
  OAI21X1 U395 ( .A(n829), .B(n588), .C(n41), .Y(n865) );
  OAI21X1 U397 ( .A(n827), .B(n588), .C(n39), .Y(n864) );
  OAI21X1 U399 ( .A(n825), .B(n588), .C(n37), .Y(n863) );
  OAI21X1 U401 ( .A(n823), .B(n588), .C(n35), .Y(n862) );
  NOR3X1 U405 ( .A(n822), .B(n838), .C(n837), .Y(n1015) );
  OAI21X1 U406 ( .A(n832), .B(n586), .C(n33), .Y(n861) );
  OAI21X1 U408 ( .A(n830), .B(n586), .C(n31), .Y(n860) );
  OAI21X1 U410 ( .A(n828), .B(n586), .C(n29), .Y(n859) );
  OAI21X1 U412 ( .A(n826), .B(n586), .C(n27), .Y(n858) );
  OAI21X1 U414 ( .A(n824), .B(n586), .C(n25), .Y(n857) );
  NOR3X1 U418 ( .A(n821), .B(n838), .C(n837), .Y(n1014) );
  OAI21X1 U419 ( .A(n831), .B(n584), .C(n23), .Y(n856) );
  OAI21X1 U421 ( .A(n829), .B(n584), .C(n21), .Y(n855) );
  OAI21X1 U423 ( .A(n827), .B(n584), .C(n19), .Y(n854) );
  OAI21X1 U425 ( .A(n825), .B(n584), .C(n17), .Y(n853) );
  OAI21X1 U427 ( .A(n823), .B(n584), .C(n15), .Y(n852) );
  NOR3X1 U431 ( .A(n836), .B(n838), .C(n822), .Y(n1013) );
  OAI21X1 U432 ( .A(n832), .B(n582), .C(n13), .Y(n851) );
  OAI21X1 U435 ( .A(n830), .B(n582), .C(n11), .Y(n850) );
  OAI21X1 U438 ( .A(n828), .B(n582), .C(n9), .Y(n849) );
  OAI21X1 U441 ( .A(n826), .B(n582), .C(n7), .Y(n848) );
  OAI21X1 U444 ( .A(n824), .B(n582), .C(n5), .Y(n847) );
  NOR3X1 U448 ( .A(n836), .B(n838), .C(n821), .Y(n1012) );
  NAND3X1 U449 ( .A(n840), .B(n842), .C(n1010), .Y(n1007) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n1010) );
  AND2X1 U2 ( .A(n646), .B(n833), .Y(n1020) );
  INVX1 U3 ( .A(rst), .Y(n833) );
  INVX1 U4 ( .A(n510), .Y(n824) );
  INVX1 U5 ( .A(n510), .Y(n823) );
  INVX1 U6 ( .A(n511), .Y(n826) );
  INVX1 U7 ( .A(n511), .Y(n825) );
  INVX1 U8 ( .A(n512), .Y(n828) );
  INVX1 U9 ( .A(n512), .Y(n827) );
  INVX1 U10 ( .A(n513), .Y(n830) );
  INVX1 U11 ( .A(n513), .Y(n829) );
  INVX1 U12 ( .A(n514), .Y(n832) );
  INVX1 U13 ( .A(n514), .Y(n831) );
  INVX2 U14 ( .A(n839), .Y(n838) );
  INVX8 U15 ( .A(N12), .Y(n839) );
  INVX1 U16 ( .A(N13), .Y(n840) );
  MUX2X1 U17 ( .B(n783), .A(n781), .S(n838), .Y(n794) );
  MUX2X1 U18 ( .B(n794), .A(n793), .S(n800), .Y(n792) );
  MUX2X1 U19 ( .B(n754), .A(n752), .S(n838), .Y(n765) );
  OR2X2 U20 ( .A(write), .B(rst), .Y(n1) );
  AND2X2 U21 ( .A(n500), .B(n501), .Y(n2) );
  AND2X2 U22 ( .A(n644), .B(n645), .Y(n3) );
  AND2X2 U23 ( .A(\mem<0><4> ), .B(n516), .Y(n4) );
  INVX1 U24 ( .A(n4), .Y(n5) );
  AND2X2 U25 ( .A(\mem<0><3> ), .B(n516), .Y(n6) );
  INVX1 U26 ( .A(n6), .Y(n7) );
  AND2X2 U27 ( .A(\mem<0><2> ), .B(n516), .Y(n8) );
  INVX1 U28 ( .A(n8), .Y(n9) );
  AND2X2 U29 ( .A(\mem<0><1> ), .B(n516), .Y(n10) );
  INVX1 U30 ( .A(n10), .Y(n11) );
  AND2X2 U31 ( .A(\mem<0><0> ), .B(n516), .Y(n12) );
  INVX1 U32 ( .A(n12), .Y(n13) );
  AND2X2 U33 ( .A(\mem<1><4> ), .B(n518), .Y(n14) );
  INVX1 U34 ( .A(n14), .Y(n15) );
  AND2X2 U35 ( .A(\mem<1><3> ), .B(n518), .Y(n16) );
  INVX1 U36 ( .A(n16), .Y(n17) );
  AND2X2 U37 ( .A(\mem<1><2> ), .B(n518), .Y(n18) );
  INVX1 U38 ( .A(n18), .Y(n19) );
  AND2X2 U39 ( .A(\mem<1><1> ), .B(n518), .Y(n20) );
  INVX1 U40 ( .A(n20), .Y(n21) );
  AND2X2 U41 ( .A(\mem<1><0> ), .B(n518), .Y(n22) );
  INVX1 U42 ( .A(n22), .Y(n23) );
  AND2X2 U43 ( .A(\mem<2><4> ), .B(n520), .Y(n24) );
  INVX1 U44 ( .A(n24), .Y(n25) );
  AND2X2 U45 ( .A(\mem<2><3> ), .B(n520), .Y(n26) );
  INVX1 U46 ( .A(n26), .Y(n27) );
  AND2X2 U47 ( .A(\mem<2><2> ), .B(n520), .Y(n28) );
  INVX1 U48 ( .A(n28), .Y(n29) );
  AND2X2 U49 ( .A(\mem<2><1> ), .B(n520), .Y(n30) );
  INVX1 U51 ( .A(n30), .Y(n31) );
  AND2X2 U53 ( .A(\mem<2><0> ), .B(n520), .Y(n32) );
  INVX1 U55 ( .A(n32), .Y(n33) );
  AND2X2 U57 ( .A(\mem<3><4> ), .B(n522), .Y(n34) );
  INVX1 U59 ( .A(n34), .Y(n35) );
  AND2X2 U60 ( .A(\mem<3><3> ), .B(n522), .Y(n36) );
  INVX1 U61 ( .A(n36), .Y(n37) );
  AND2X2 U63 ( .A(\mem<3><2> ), .B(n522), .Y(n38) );
  INVX1 U65 ( .A(n38), .Y(n39) );
  AND2X2 U67 ( .A(\mem<3><1> ), .B(n522), .Y(n40) );
  INVX1 U69 ( .A(n40), .Y(n41) );
  AND2X2 U71 ( .A(\mem<3><0> ), .B(n522), .Y(n42) );
  INVX1 U72 ( .A(n42), .Y(n43) );
  AND2X2 U73 ( .A(\mem<4><4> ), .B(n524), .Y(n44) );
  INVX1 U75 ( .A(n44), .Y(n45) );
  AND2X2 U77 ( .A(\mem<4><3> ), .B(n524), .Y(n46) );
  INVX1 U79 ( .A(n46), .Y(n47) );
  AND2X2 U81 ( .A(\mem<4><2> ), .B(n524), .Y(n48) );
  INVX1 U83 ( .A(n48), .Y(n49) );
  AND2X2 U84 ( .A(\mem<4><1> ), .B(n524), .Y(n50) );
  INVX1 U85 ( .A(n50), .Y(n51) );
  AND2X2 U87 ( .A(\mem<4><0> ), .B(n524), .Y(n52) );
  INVX1 U89 ( .A(n52), .Y(n53) );
  AND2X2 U91 ( .A(\mem<5><4> ), .B(n526), .Y(n54) );
  INVX1 U93 ( .A(n54), .Y(n55) );
  AND2X2 U95 ( .A(\mem<5><3> ), .B(n526), .Y(n58) );
  INVX1 U96 ( .A(n58), .Y(n59) );
  AND2X2 U97 ( .A(\mem<5><2> ), .B(n526), .Y(n60) );
  INVX1 U99 ( .A(n60), .Y(n61) );
  AND2X2 U101 ( .A(\mem<5><1> ), .B(n526), .Y(n62) );
  INVX1 U103 ( .A(n62), .Y(n63) );
  AND2X2 U105 ( .A(\mem<5><0> ), .B(n526), .Y(n64) );
  INVX1 U107 ( .A(n64), .Y(n66) );
  AND2X2 U108 ( .A(\mem<6><4> ), .B(n528), .Y(n67) );
  INVX1 U109 ( .A(n67), .Y(n68) );
  AND2X2 U111 ( .A(\mem<6><3> ), .B(n528), .Y(n69) );
  INVX1 U113 ( .A(n69), .Y(n70) );
  AND2X2 U115 ( .A(\mem<6><2> ), .B(n528), .Y(n71) );
  INVX1 U117 ( .A(n71), .Y(n72) );
  AND2X2 U119 ( .A(\mem<6><1> ), .B(n528), .Y(n74) );
  INVX1 U120 ( .A(n74), .Y(n75) );
  AND2X2 U121 ( .A(\mem<6><0> ), .B(n528), .Y(n76) );
  INVX1 U123 ( .A(n76), .Y(n77) );
  AND2X2 U125 ( .A(\mem<7><4> ), .B(n530), .Y(n78) );
  INVX1 U127 ( .A(n78), .Y(n79) );
  AND2X2 U129 ( .A(\mem<7><3> ), .B(n530), .Y(n80) );
  INVX1 U131 ( .A(n80), .Y(n82) );
  AND2X2 U132 ( .A(\mem<7><2> ), .B(n530), .Y(n83) );
  INVX1 U133 ( .A(n83), .Y(n84) );
  AND2X2 U135 ( .A(\mem<7><1> ), .B(n530), .Y(n85) );
  INVX1 U137 ( .A(n85), .Y(n86) );
  AND2X2 U139 ( .A(\mem<7><0> ), .B(n530), .Y(n87) );
  INVX1 U141 ( .A(n87), .Y(n88) );
  AND2X2 U143 ( .A(\mem<8><4> ), .B(n532), .Y(n90) );
  INVX1 U144 ( .A(n90), .Y(n91) );
  AND2X2 U145 ( .A(\mem<8><3> ), .B(n532), .Y(n92) );
  INVX1 U148 ( .A(n92), .Y(n93) );
  AND2X2 U150 ( .A(\mem<8><2> ), .B(n532), .Y(n94) );
  INVX1 U152 ( .A(n94), .Y(n95) );
  AND2X2 U154 ( .A(\mem<8><1> ), .B(n532), .Y(n96) );
  INVX1 U156 ( .A(n96), .Y(n98) );
  AND2X2 U157 ( .A(\mem<8><0> ), .B(n532), .Y(n99) );
  INVX1 U158 ( .A(n99), .Y(n100) );
  AND2X2 U160 ( .A(\mem<9><4> ), .B(n534), .Y(n101) );
  INVX1 U162 ( .A(n101), .Y(n102) );
  AND2X2 U164 ( .A(\mem<9><3> ), .B(n534), .Y(n103) );
  INVX1 U166 ( .A(n103), .Y(n104) );
  AND2X2 U168 ( .A(\mem<9><2> ), .B(n534), .Y(n106) );
  INVX1 U169 ( .A(n106), .Y(n107) );
  AND2X2 U170 ( .A(\mem<9><1> ), .B(n534), .Y(n108) );
  INVX1 U172 ( .A(n108), .Y(n109) );
  AND2X2 U174 ( .A(\mem<9><0> ), .B(n534), .Y(n110) );
  INVX1 U176 ( .A(n110), .Y(n111) );
  AND2X2 U178 ( .A(\mem<10><4> ), .B(n536), .Y(n112) );
  INVX1 U180 ( .A(n112), .Y(n116) );
  AND2X2 U181 ( .A(\mem<10><3> ), .B(n536), .Y(n117) );
  INVX1 U182 ( .A(n117), .Y(n118) );
  AND2X2 U184 ( .A(\mem<10><2> ), .B(n536), .Y(n119) );
  INVX1 U186 ( .A(n119), .Y(n120) );
  AND2X2 U188 ( .A(\mem<10><1> ), .B(n536), .Y(n121) );
  INVX1 U190 ( .A(n121), .Y(n122) );
  AND2X2 U192 ( .A(\mem<10><0> ), .B(n536), .Y(n123) );
  INVX1 U193 ( .A(n123), .Y(n124) );
  AND2X2 U194 ( .A(\mem<11><4> ), .B(n538), .Y(n125) );
  INVX1 U196 ( .A(n125), .Y(n126) );
  AND2X2 U198 ( .A(\mem<11><3> ), .B(n538), .Y(n127) );
  INVX1 U200 ( .A(n127), .Y(n128) );
  AND2X2 U202 ( .A(\mem<11><2> ), .B(n538), .Y(n129) );
  INVX1 U204 ( .A(n129), .Y(n130) );
  AND2X2 U205 ( .A(\mem<11><1> ), .B(n538), .Y(n131) );
  INVX1 U206 ( .A(n131), .Y(n132) );
  AND2X2 U208 ( .A(\mem<11><0> ), .B(n538), .Y(n133) );
  INVX1 U210 ( .A(n133), .Y(n134) );
  AND2X2 U212 ( .A(\mem<12><4> ), .B(n540), .Y(n135) );
  INVX1 U214 ( .A(n135), .Y(n136) );
  AND2X2 U216 ( .A(\mem<12><3> ), .B(n540), .Y(n137) );
  INVX1 U217 ( .A(n137), .Y(n138) );
  AND2X2 U218 ( .A(\mem<12><2> ), .B(n540), .Y(n139) );
  INVX1 U220 ( .A(n139), .Y(n140) );
  AND2X2 U222 ( .A(\mem<12><1> ), .B(n540), .Y(n141) );
  INVX1 U224 ( .A(n141), .Y(n142) );
  AND2X2 U226 ( .A(\mem<12><0> ), .B(n540), .Y(n143) );
  INVX1 U228 ( .A(n143), .Y(n144) );
  AND2X2 U229 ( .A(\mem<13><4> ), .B(n542), .Y(n145) );
  INVX1 U230 ( .A(n145), .Y(n146) );
  AND2X2 U232 ( .A(\mem<13><3> ), .B(n542), .Y(n147) );
  INVX1 U234 ( .A(n147), .Y(n148) );
  AND2X2 U236 ( .A(\mem<13><2> ), .B(n542), .Y(n149) );
  INVX1 U238 ( .A(n149), .Y(n150) );
  AND2X2 U240 ( .A(\mem<13><1> ), .B(n542), .Y(n151) );
  INVX1 U241 ( .A(n151), .Y(n152) );
  AND2X2 U242 ( .A(\mem<13><0> ), .B(n542), .Y(n153) );
  INVX1 U245 ( .A(n153), .Y(n154) );
  AND2X2 U247 ( .A(\mem<14><4> ), .B(n544), .Y(n155) );
  INVX1 U249 ( .A(n155), .Y(n156) );
  AND2X2 U251 ( .A(\mem<14><3> ), .B(n544), .Y(n157) );
  INVX1 U253 ( .A(n157), .Y(n158) );
  AND2X2 U254 ( .A(\mem<14><2> ), .B(n544), .Y(n159) );
  INVX1 U255 ( .A(n159), .Y(n160) );
  AND2X2 U257 ( .A(\mem<14><1> ), .B(n544), .Y(n161) );
  INVX1 U259 ( .A(n161), .Y(n162) );
  AND2X2 U261 ( .A(\mem<14><0> ), .B(n544), .Y(n163) );
  INVX1 U263 ( .A(n163), .Y(n164) );
  AND2X2 U265 ( .A(\mem<15><4> ), .B(n546), .Y(n165) );
  INVX1 U266 ( .A(n165), .Y(n166) );
  AND2X2 U267 ( .A(\mem<15><3> ), .B(n546), .Y(n167) );
  INVX1 U269 ( .A(n167), .Y(n168) );
  AND2X2 U271 ( .A(\mem<15><2> ), .B(n546), .Y(n169) );
  INVX1 U273 ( .A(n169), .Y(n170) );
  AND2X2 U275 ( .A(\mem<15><1> ), .B(n546), .Y(n171) );
  INVX1 U277 ( .A(n171), .Y(n173) );
  AND2X2 U278 ( .A(\mem<15><0> ), .B(n546), .Y(n174) );
  INVX1 U279 ( .A(n174), .Y(n175) );
  AND2X2 U281 ( .A(\mem<16><4> ), .B(n548), .Y(n176) );
  INVX1 U283 ( .A(n176), .Y(n177) );
  AND2X2 U285 ( .A(\mem<16><3> ), .B(n548), .Y(n178) );
  INVX1 U287 ( .A(n178), .Y(n179) );
  AND2X2 U289 ( .A(\mem<16><2> ), .B(n548), .Y(n180) );
  INVX1 U290 ( .A(n180), .Y(n181) );
  AND2X2 U291 ( .A(\mem<16><1> ), .B(n548), .Y(n182) );
  INVX1 U293 ( .A(n182), .Y(n183) );
  AND2X2 U295 ( .A(\mem<16><0> ), .B(n548), .Y(n184) );
  INVX1 U297 ( .A(n184), .Y(n185) );
  AND2X2 U299 ( .A(\mem<17><4> ), .B(n550), .Y(n186) );
  INVX1 U301 ( .A(n186), .Y(n187) );
  AND2X2 U302 ( .A(\mem<17><3> ), .B(n550), .Y(n188) );
  INVX1 U303 ( .A(n188), .Y(n189) );
  AND2X2 U305 ( .A(\mem<17><2> ), .B(n550), .Y(n190) );
  INVX1 U307 ( .A(n190), .Y(n191) );
  AND2X2 U309 ( .A(\mem<17><1> ), .B(n550), .Y(n192) );
  INVX1 U311 ( .A(n192), .Y(n193) );
  AND2X2 U313 ( .A(\mem<17><0> ), .B(n550), .Y(n194) );
  INVX1 U314 ( .A(n194), .Y(n195) );
  AND2X2 U315 ( .A(\mem<18><4> ), .B(n552), .Y(n196) );
  INVX1 U317 ( .A(n196), .Y(n197) );
  AND2X2 U319 ( .A(\mem<18><3> ), .B(n552), .Y(n198) );
  INVX1 U321 ( .A(n198), .Y(n199) );
  AND2X2 U323 ( .A(\mem<18><2> ), .B(n552), .Y(n200) );
  INVX1 U325 ( .A(n200), .Y(n201) );
  AND2X2 U326 ( .A(\mem<18><1> ), .B(n552), .Y(n202) );
  INVX1 U327 ( .A(n202), .Y(n203) );
  AND2X2 U329 ( .A(\mem<18><0> ), .B(n552), .Y(n204) );
  INVX1 U331 ( .A(n204), .Y(n205) );
  AND2X2 U333 ( .A(\mem<19><4> ), .B(n554), .Y(n206) );
  INVX1 U335 ( .A(n206), .Y(n207) );
  AND2X2 U337 ( .A(\mem<19><3> ), .B(n554), .Y(n208) );
  INVX1 U338 ( .A(n208), .Y(n209) );
  AND2X2 U339 ( .A(\mem<19><2> ), .B(n554), .Y(n210) );
  INVX1 U342 ( .A(n210), .Y(n211) );
  AND2X2 U344 ( .A(\mem<19><1> ), .B(n554), .Y(n212) );
  INVX1 U346 ( .A(n212), .Y(n213) );
  AND2X2 U348 ( .A(\mem<19><0> ), .B(n554), .Y(n214) );
  INVX1 U350 ( .A(n214), .Y(n215) );
  AND2X2 U351 ( .A(\mem<20><4> ), .B(n556), .Y(n216) );
  INVX1 U352 ( .A(n216), .Y(n217) );
  AND2X2 U355 ( .A(\mem<20><3> ), .B(n556), .Y(n218) );
  INVX1 U357 ( .A(n218), .Y(n219) );
  AND2X2 U359 ( .A(\mem<20><2> ), .B(n556), .Y(n220) );
  INVX1 U361 ( .A(n220), .Y(n221) );
  AND2X2 U363 ( .A(\mem<20><1> ), .B(n556), .Y(n222) );
  INVX1 U364 ( .A(n222), .Y(n223) );
  AND2X2 U365 ( .A(\mem<20><0> ), .B(n556), .Y(n224) );
  INVX1 U368 ( .A(n224), .Y(n225) );
  AND2X2 U370 ( .A(\mem<21><4> ), .B(n558), .Y(n226) );
  INVX1 U372 ( .A(n226), .Y(n227) );
  AND2X2 U374 ( .A(\mem<21><3> ), .B(n558), .Y(n228) );
  INVX1 U376 ( .A(n228), .Y(n230) );
  AND2X2 U377 ( .A(\mem<21><2> ), .B(n558), .Y(n231) );
  INVX1 U378 ( .A(n231), .Y(n232) );
  AND2X2 U381 ( .A(\mem<21><1> ), .B(n558), .Y(n233) );
  INVX1 U383 ( .A(n233), .Y(n234) );
  AND2X2 U385 ( .A(\mem<21><0> ), .B(n558), .Y(n235) );
  INVX1 U387 ( .A(n235), .Y(n236) );
  AND2X2 U389 ( .A(\mem<22><4> ), .B(n560), .Y(n237) );
  INVX1 U390 ( .A(n237), .Y(n238) );
  AND2X2 U391 ( .A(\mem<22><3> ), .B(n560), .Y(n239) );
  INVX1 U394 ( .A(n239), .Y(n240) );
  AND2X2 U396 ( .A(\mem<22><2> ), .B(n560), .Y(n241) );
  INVX1 U398 ( .A(n241), .Y(n242) );
  AND2X2 U400 ( .A(\mem<22><1> ), .B(n560), .Y(n243) );
  INVX1 U402 ( .A(n243), .Y(n244) );
  AND2X2 U403 ( .A(\mem<22><0> ), .B(n560), .Y(n245) );
  INVX1 U404 ( .A(n245), .Y(n246) );
  AND2X2 U407 ( .A(\mem<23><4> ), .B(n562), .Y(n247) );
  INVX1 U409 ( .A(n247), .Y(n248) );
  AND2X2 U411 ( .A(\mem<23><3> ), .B(n562), .Y(n249) );
  INVX1 U413 ( .A(n249), .Y(n250) );
  AND2X2 U415 ( .A(\mem<23><2> ), .B(n562), .Y(n251) );
  INVX1 U416 ( .A(n251), .Y(n252) );
  AND2X2 U417 ( .A(\mem<23><1> ), .B(n562), .Y(n253) );
  INVX1 U420 ( .A(n253), .Y(n254) );
  AND2X2 U422 ( .A(\mem<23><0> ), .B(n562), .Y(n255) );
  INVX1 U424 ( .A(n255), .Y(n256) );
  AND2X2 U426 ( .A(\mem<24><4> ), .B(n564), .Y(n257) );
  INVX1 U428 ( .A(n257), .Y(n258) );
  AND2X2 U429 ( .A(\mem<24><3> ), .B(n564), .Y(n259) );
  INVX1 U430 ( .A(n259), .Y(n260) );
  AND2X2 U433 ( .A(\mem<24><2> ), .B(n564), .Y(n261) );
  INVX1 U434 ( .A(n261), .Y(n262) );
  AND2X2 U436 ( .A(\mem<24><1> ), .B(n564), .Y(n263) );
  INVX1 U437 ( .A(n263), .Y(n264) );
  AND2X2 U439 ( .A(\mem<24><0> ), .B(n564), .Y(n265) );
  INVX1 U440 ( .A(n265), .Y(n266) );
  AND2X2 U442 ( .A(\mem<25><4> ), .B(n566), .Y(n267) );
  INVX1 U443 ( .A(n267), .Y(n268) );
  AND2X2 U445 ( .A(\mem<25><3> ), .B(n566), .Y(n269) );
  INVX1 U446 ( .A(n269), .Y(n270) );
  AND2X2 U447 ( .A(\mem<25><2> ), .B(n566), .Y(n271) );
  INVX1 U451 ( .A(n271), .Y(n272) );
  AND2X2 U452 ( .A(\mem<25><1> ), .B(n566), .Y(n273) );
  INVX1 U453 ( .A(n273), .Y(n274) );
  AND2X2 U454 ( .A(\mem<25><0> ), .B(n566), .Y(n275) );
  INVX1 U455 ( .A(n275), .Y(n276) );
  AND2X2 U456 ( .A(\mem<26><4> ), .B(n568), .Y(n277) );
  INVX1 U457 ( .A(n277), .Y(n278) );
  AND2X2 U458 ( .A(\mem<26><3> ), .B(n568), .Y(n279) );
  INVX1 U459 ( .A(n279), .Y(n280) );
  AND2X2 U460 ( .A(\mem<26><2> ), .B(n568), .Y(n281) );
  INVX1 U461 ( .A(n281), .Y(n282) );
  AND2X2 U462 ( .A(\mem<26><1> ), .B(n568), .Y(n283) );
  INVX1 U463 ( .A(n283), .Y(n284) );
  AND2X2 U464 ( .A(\mem<26><0> ), .B(n568), .Y(n285) );
  INVX1 U465 ( .A(n285), .Y(n287) );
  AND2X2 U466 ( .A(\mem<27><4> ), .B(n570), .Y(n448) );
  INVX1 U467 ( .A(n448), .Y(n449) );
  AND2X2 U468 ( .A(\mem<27><3> ), .B(n570), .Y(n450) );
  INVX1 U469 ( .A(n450), .Y(n451) );
  AND2X2 U470 ( .A(\mem<27><2> ), .B(n570), .Y(n452) );
  INVX1 U471 ( .A(n452), .Y(n453) );
  AND2X2 U472 ( .A(\mem<27><1> ), .B(n570), .Y(n454) );
  INVX1 U473 ( .A(n454), .Y(n455) );
  AND2X2 U474 ( .A(\mem<27><0> ), .B(n570), .Y(n456) );
  INVX1 U475 ( .A(n456), .Y(n457) );
  AND2X2 U476 ( .A(\mem<28><4> ), .B(n572), .Y(n458) );
  INVX1 U477 ( .A(n458), .Y(n459) );
  AND2X2 U478 ( .A(\mem<28><3> ), .B(n572), .Y(n460) );
  INVX1 U479 ( .A(n460), .Y(n461) );
  AND2X2 U480 ( .A(\mem<28><2> ), .B(n572), .Y(n462) );
  INVX1 U481 ( .A(n462), .Y(n463) );
  AND2X2 U482 ( .A(\mem<28><1> ), .B(n572), .Y(n464) );
  INVX1 U483 ( .A(n464), .Y(n465) );
  AND2X2 U484 ( .A(\mem<28><0> ), .B(n572), .Y(n466) );
  INVX1 U485 ( .A(n466), .Y(n467) );
  AND2X2 U486 ( .A(\mem<29><4> ), .B(n574), .Y(n468) );
  INVX1 U487 ( .A(n468), .Y(n469) );
  AND2X2 U488 ( .A(\mem<29><3> ), .B(n574), .Y(n470) );
  INVX1 U489 ( .A(n470), .Y(n471) );
  AND2X2 U490 ( .A(\mem<29><2> ), .B(n574), .Y(n472) );
  INVX1 U491 ( .A(n472), .Y(n473) );
  AND2X2 U492 ( .A(\mem<29><1> ), .B(n574), .Y(n474) );
  INVX1 U493 ( .A(n474), .Y(n475) );
  AND2X2 U494 ( .A(\mem<29><0> ), .B(n574), .Y(n476) );
  INVX1 U495 ( .A(n476), .Y(n477) );
  AND2X2 U496 ( .A(\mem<30><4> ), .B(n576), .Y(n478) );
  INVX1 U497 ( .A(n478), .Y(n479) );
  AND2X2 U498 ( .A(\mem<30><3> ), .B(n576), .Y(n480) );
  INVX1 U499 ( .A(n480), .Y(n481) );
  AND2X2 U500 ( .A(\mem<30><2> ), .B(n576), .Y(n482) );
  INVX1 U501 ( .A(n482), .Y(n483) );
  AND2X2 U502 ( .A(\mem<30><1> ), .B(n576), .Y(n484) );
  INVX1 U503 ( .A(n484), .Y(n485) );
  AND2X2 U504 ( .A(\mem<30><0> ), .B(n576), .Y(n486) );
  INVX1 U505 ( .A(n486), .Y(n487) );
  AND2X2 U506 ( .A(\mem<31><4> ), .B(n578), .Y(n488) );
  INVX1 U507 ( .A(n488), .Y(n489) );
  AND2X2 U508 ( .A(\mem<31><3> ), .B(n578), .Y(n490) );
  INVX1 U509 ( .A(n490), .Y(n491) );
  AND2X2 U510 ( .A(\mem<31><2> ), .B(n578), .Y(n492) );
  INVX1 U511 ( .A(n492), .Y(n493) );
  AND2X2 U512 ( .A(\mem<31><1> ), .B(n578), .Y(n494) );
  INVX1 U513 ( .A(n494), .Y(n495) );
  AND2X2 U514 ( .A(\mem<31><0> ), .B(n578), .Y(n496) );
  INVX1 U515 ( .A(n496), .Y(n497) );
  OR2X2 U516 ( .A(write), .B(rst), .Y(n498) );
  MUX2X1 U517 ( .B(n694), .A(n693), .S(n805), .Y(n692) );
  INVX4 U518 ( .A(n834), .Y(n810) );
  MUX2X1 U519 ( .B(\mem<11><1> ), .A(\mem<10><1> ), .S(n811), .Y(n697) );
  INVX2 U520 ( .A(n836), .Y(n804) );
  MUX2X1 U521 ( .B(n676), .A(n675), .S(n800), .Y(n674) );
  NAND2X1 U522 ( .A(\mem<14><4> ), .B(n499), .Y(n500) );
  NAND2X1 U523 ( .A(\mem<15><4> ), .B(n814), .Y(n501) );
  INVX1 U524 ( .A(n813), .Y(n499) );
  INVX1 U525 ( .A(n1), .Y(n502) );
  INVX1 U526 ( .A(n1), .Y(n503) );
  BUFX2 U527 ( .A(n1007), .Y(n504) );
  INVX1 U528 ( .A(n504), .Y(n843) );
  BUFX2 U529 ( .A(n1008), .Y(n505) );
  INVX1 U530 ( .A(n505), .Y(n844) );
  BUFX2 U531 ( .A(n1009), .Y(n506) );
  INVX1 U532 ( .A(n506), .Y(n845) );
  BUFX2 U533 ( .A(n1011), .Y(n507) );
  INVX1 U534 ( .A(n507), .Y(n846) );
  INVX1 U535 ( .A(n1), .Y(n508) );
  INVX1 U536 ( .A(n498), .Y(n509) );
  AND2X1 U537 ( .A(\data_in<4> ), .B(n1020), .Y(n510) );
  AND2X1 U538 ( .A(\data_in<3> ), .B(n1020), .Y(n511) );
  AND2X1 U539 ( .A(\data_in<2> ), .B(n1020), .Y(n512) );
  AND2X1 U540 ( .A(\data_in<1> ), .B(n1020), .Y(n513) );
  AND2X1 U541 ( .A(\data_in<0> ), .B(n1020), .Y(n514) );
  AND2X1 U542 ( .A(n581), .B(n1020), .Y(n515) );
  INVX1 U543 ( .A(n515), .Y(n516) );
  AND2X1 U544 ( .A(n583), .B(n1020), .Y(n517) );
  INVX1 U545 ( .A(n517), .Y(n518) );
  AND2X1 U546 ( .A(n585), .B(n1020), .Y(n519) );
  INVX1 U547 ( .A(n519), .Y(n520) );
  AND2X1 U548 ( .A(n587), .B(n1020), .Y(n521) );
  INVX1 U549 ( .A(n521), .Y(n522) );
  AND2X1 U550 ( .A(n589), .B(n1020), .Y(n523) );
  INVX1 U551 ( .A(n523), .Y(n524) );
  AND2X1 U552 ( .A(n591), .B(n1020), .Y(n525) );
  INVX1 U553 ( .A(n525), .Y(n526) );
  AND2X1 U554 ( .A(n593), .B(n1020), .Y(n527) );
  INVX1 U555 ( .A(n527), .Y(n528) );
  AND2X1 U556 ( .A(n595), .B(n1020), .Y(n529) );
  INVX1 U557 ( .A(n529), .Y(n530) );
  AND2X1 U558 ( .A(n597), .B(n1020), .Y(n531) );
  INVX1 U559 ( .A(n531), .Y(n532) );
  AND2X1 U560 ( .A(n599), .B(n1020), .Y(n533) );
  INVX1 U561 ( .A(n533), .Y(n534) );
  AND2X1 U562 ( .A(n601), .B(n1020), .Y(n535) );
  INVX1 U563 ( .A(n535), .Y(n536) );
  AND2X1 U564 ( .A(n603), .B(n1020), .Y(n537) );
  INVX1 U565 ( .A(n537), .Y(n538) );
  AND2X1 U566 ( .A(n605), .B(n1020), .Y(n539) );
  INVX1 U567 ( .A(n539), .Y(n540) );
  AND2X1 U568 ( .A(n607), .B(n1020), .Y(n541) );
  INVX1 U569 ( .A(n541), .Y(n542) );
  AND2X1 U570 ( .A(n609), .B(n1020), .Y(n543) );
  INVX1 U571 ( .A(n543), .Y(n544) );
  AND2X1 U572 ( .A(n611), .B(n1020), .Y(n545) );
  INVX1 U573 ( .A(n545), .Y(n546) );
  AND2X1 U574 ( .A(n613), .B(n1020), .Y(n547) );
  INVX1 U575 ( .A(n547), .Y(n548) );
  AND2X1 U576 ( .A(n615), .B(n1020), .Y(n549) );
  INVX1 U577 ( .A(n549), .Y(n550) );
  AND2X1 U578 ( .A(n618), .B(n1020), .Y(n551) );
  INVX1 U579 ( .A(n551), .Y(n552) );
  AND2X1 U580 ( .A(n619), .B(n1020), .Y(n553) );
  INVX1 U581 ( .A(n553), .Y(n554) );
  AND2X1 U582 ( .A(n622), .B(n1020), .Y(n555) );
  INVX1 U583 ( .A(n555), .Y(n556) );
  AND2X1 U584 ( .A(n623), .B(n1020), .Y(n557) );
  INVX1 U585 ( .A(n557), .Y(n558) );
  AND2X1 U586 ( .A(n626), .B(n1020), .Y(n559) );
  INVX1 U587 ( .A(n559), .Y(n560) );
  AND2X1 U588 ( .A(n627), .B(n1020), .Y(n561) );
  INVX1 U589 ( .A(n561), .Y(n562) );
  AND2X1 U590 ( .A(n629), .B(n1020), .Y(n563) );
  INVX1 U591 ( .A(n563), .Y(n564) );
  AND2X1 U592 ( .A(n631), .B(n1020), .Y(n565) );
  INVX1 U593 ( .A(n565), .Y(n566) );
  AND2X1 U594 ( .A(n633), .B(n1020), .Y(n567) );
  INVX1 U595 ( .A(n567), .Y(n568) );
  AND2X1 U596 ( .A(n635), .B(n1020), .Y(n569) );
  INVX1 U597 ( .A(n569), .Y(n570) );
  AND2X1 U598 ( .A(n637), .B(n1020), .Y(n571) );
  INVX1 U599 ( .A(n571), .Y(n572) );
  AND2X1 U600 ( .A(n639), .B(n1020), .Y(n573) );
  INVX1 U601 ( .A(n573), .Y(n574) );
  AND2X1 U602 ( .A(n641), .B(n1020), .Y(n575) );
  INVX1 U603 ( .A(n575), .Y(n576) );
  AND2X1 U604 ( .A(n580), .B(n1020), .Y(n577) );
  INVX1 U605 ( .A(n577), .Y(n578) );
  INVX1 U606 ( .A(n580), .Y(n579) );
  AND2X1 U607 ( .A(n1019), .B(n846), .Y(n580) );
  AND2X1 U608 ( .A(n843), .B(n1012), .Y(n581) );
  INVX1 U609 ( .A(n581), .Y(n582) );
  AND2X1 U610 ( .A(n843), .B(n1013), .Y(n583) );
  INVX1 U611 ( .A(n583), .Y(n584) );
  AND2X1 U612 ( .A(n843), .B(n1014), .Y(n585) );
  INVX1 U613 ( .A(n585), .Y(n586) );
  AND2X1 U614 ( .A(n843), .B(n1015), .Y(n587) );
  INVX1 U615 ( .A(n587), .Y(n588) );
  AND2X1 U616 ( .A(n843), .B(n1016), .Y(n589) );
  INVX1 U617 ( .A(n589), .Y(n590) );
  AND2X1 U618 ( .A(n843), .B(n1017), .Y(n591) );
  INVX1 U619 ( .A(n591), .Y(n592) );
  AND2X1 U620 ( .A(n843), .B(n1018), .Y(n593) );
  INVX1 U621 ( .A(n593), .Y(n594) );
  AND2X1 U622 ( .A(n843), .B(n1019), .Y(n595) );
  INVX1 U623 ( .A(n595), .Y(n596) );
  AND2X1 U624 ( .A(n844), .B(n1012), .Y(n597) );
  INVX1 U625 ( .A(n597), .Y(n598) );
  AND2X1 U626 ( .A(n844), .B(n1013), .Y(n599) );
  INVX1 U627 ( .A(n599), .Y(n600) );
  AND2X1 U628 ( .A(n844), .B(n1014), .Y(n601) );
  INVX1 U629 ( .A(n601), .Y(n602) );
  AND2X1 U630 ( .A(n844), .B(n1015), .Y(n603) );
  INVX1 U631 ( .A(n603), .Y(n604) );
  AND2X1 U632 ( .A(n844), .B(n1016), .Y(n605) );
  INVX1 U633 ( .A(n605), .Y(n606) );
  AND2X1 U634 ( .A(n844), .B(n1017), .Y(n607) );
  INVX1 U635 ( .A(n607), .Y(n608) );
  AND2X1 U636 ( .A(n844), .B(n1018), .Y(n609) );
  INVX1 U637 ( .A(n609), .Y(n610) );
  AND2X1 U638 ( .A(n844), .B(n1019), .Y(n611) );
  INVX1 U639 ( .A(n611), .Y(n612) );
  AND2X1 U640 ( .A(n845), .B(n1012), .Y(n613) );
  INVX1 U641 ( .A(n613), .Y(n614) );
  AND2X1 U642 ( .A(n845), .B(n1013), .Y(n615) );
  INVX1 U643 ( .A(n615), .Y(n616) );
  INVX1 U644 ( .A(n618), .Y(n617) );
  AND2X1 U645 ( .A(n845), .B(n1014), .Y(n618) );
  AND2X1 U646 ( .A(n845), .B(n1015), .Y(n619) );
  INVX1 U647 ( .A(n619), .Y(n620) );
  INVX1 U648 ( .A(n622), .Y(n621) );
  AND2X1 U649 ( .A(n845), .B(n1016), .Y(n622) );
  AND2X1 U650 ( .A(n845), .B(n1017), .Y(n623) );
  INVX1 U651 ( .A(n623), .Y(n624) );
  INVX1 U652 ( .A(n626), .Y(n625) );
  AND2X1 U653 ( .A(n845), .B(n1018), .Y(n626) );
  AND2X1 U654 ( .A(n845), .B(n1019), .Y(n627) );
  INVX1 U655 ( .A(n627), .Y(n628) );
  AND2X1 U656 ( .A(n1012), .B(n846), .Y(n629) );
  INVX1 U657 ( .A(n629), .Y(n630) );
  AND2X1 U658 ( .A(n1013), .B(n846), .Y(n631) );
  INVX1 U659 ( .A(n631), .Y(n632) );
  AND2X1 U660 ( .A(n1014), .B(n846), .Y(n633) );
  INVX1 U661 ( .A(n633), .Y(n634) );
  AND2X1 U662 ( .A(n1015), .B(n846), .Y(n635) );
  INVX1 U663 ( .A(n635), .Y(n636) );
  AND2X1 U664 ( .A(n1016), .B(n846), .Y(n637) );
  INVX1 U665 ( .A(n637), .Y(n638) );
  AND2X1 U666 ( .A(n1017), .B(n846), .Y(n639) );
  INVX1 U667 ( .A(n639), .Y(n640) );
  AND2X1 U668 ( .A(n1018), .B(n846), .Y(n641) );
  INVX1 U669 ( .A(n641), .Y(n642) );
  INVX4 U670 ( .A(n839), .Y(n802) );
  INVX8 U671 ( .A(n805), .Y(n808) );
  INVX8 U672 ( .A(n835), .Y(n834) );
  MUX2X1 U673 ( .B(n737), .A(n740), .S(n839), .Y(n751) );
  NAND2X1 U674 ( .A(\mem<14><3> ), .B(n643), .Y(n644) );
  NAND2X1 U675 ( .A(\mem<15><3> ), .B(n815), .Y(n645) );
  INVX1 U676 ( .A(n813), .Y(n643) );
  MUX2X1 U677 ( .B(\mem<9><3> ), .A(\mem<8><3> ), .S(n812), .Y(n755) );
  INVX4 U678 ( .A(N11), .Y(n837) );
  MUX2X1 U679 ( .B(n756), .A(n755), .S(n805), .Y(n754) );
  BUFX2 U680 ( .A(write), .Y(n646) );
  INVX1 U681 ( .A(n795), .Y(N21) );
  INVX1 U682 ( .A(n796), .Y(N20) );
  MUX2X1 U683 ( .B(n648), .A(n649), .S(n809), .Y(n647) );
  MUX2X1 U684 ( .B(n651), .A(n652), .S(n809), .Y(n650) );
  MUX2X1 U685 ( .B(n654), .A(n655), .S(n809), .Y(n653) );
  MUX2X1 U686 ( .B(n657), .A(n658), .S(n809), .Y(n656) );
  MUX2X1 U687 ( .B(n660), .A(n661), .S(n801), .Y(n659) );
  MUX2X1 U688 ( .B(n663), .A(n664), .S(n809), .Y(n662) );
  MUX2X1 U689 ( .B(n666), .A(n667), .S(n809), .Y(n665) );
  MUX2X1 U690 ( .B(n669), .A(n670), .S(n809), .Y(n668) );
  MUX2X1 U691 ( .B(n672), .A(n673), .S(n809), .Y(n671) );
  MUX2X1 U692 ( .B(n678), .A(n679), .S(n809), .Y(n677) );
  MUX2X1 U693 ( .B(n681), .A(n682), .S(n809), .Y(n680) );
  MUX2X1 U694 ( .B(n684), .A(n685), .S(n809), .Y(n683) );
  MUX2X1 U695 ( .B(n687), .A(n688), .S(n809), .Y(n686) );
  MUX2X1 U696 ( .B(n690), .A(n691), .S(n801), .Y(n689) );
  MUX2X1 U697 ( .B(n696), .A(n697), .S(n807), .Y(n695) );
  MUX2X1 U698 ( .B(n699), .A(n700), .S(n807), .Y(n698) );
  MUX2X1 U699 ( .B(n702), .A(n703), .S(n806), .Y(n701) );
  MUX2X1 U700 ( .B(n705), .A(n706), .S(n801), .Y(n704) );
  MUX2X1 U701 ( .B(n708), .A(n709), .S(n806), .Y(n707) );
  MUX2X1 U702 ( .B(n711), .A(n712), .S(n807), .Y(n710) );
  MUX2X1 U703 ( .B(n714), .A(n715), .S(n806), .Y(n713) );
  MUX2X1 U704 ( .B(n717), .A(n718), .S(n806), .Y(n716) );
  MUX2X1 U705 ( .B(n720), .A(n721), .S(n801), .Y(n719) );
  MUX2X1 U706 ( .B(n723), .A(n724), .S(n806), .Y(n722) );
  MUX2X1 U707 ( .B(n726), .A(n727), .S(n808), .Y(n725) );
  MUX2X1 U708 ( .B(n729), .A(n730), .S(n807), .Y(n728) );
  MUX2X1 U709 ( .B(n732), .A(n733), .S(n808), .Y(n731) );
  MUX2X1 U710 ( .B(n735), .A(n736), .S(n801), .Y(n734) );
  MUX2X1 U711 ( .B(n738), .A(n739), .S(n807), .Y(n737) );
  MUX2X1 U712 ( .B(n741), .A(n742), .S(n806), .Y(n740) );
  MUX2X1 U713 ( .B(n744), .A(n745), .S(n807), .Y(n743) );
  MUX2X1 U714 ( .B(n747), .A(n748), .S(n807), .Y(n746) );
  MUX2X1 U715 ( .B(n750), .A(n751), .S(n801), .Y(n749) );
  MUX2X1 U716 ( .B(n753), .A(n3), .S(n807), .Y(n752) );
  MUX2X1 U717 ( .B(n758), .A(n759), .S(n806), .Y(n757) );
  MUX2X1 U718 ( .B(n761), .A(n762), .S(n808), .Y(n760) );
  MUX2X1 U719 ( .B(n764), .A(n765), .S(n801), .Y(n763) );
  MUX2X1 U720 ( .B(n767), .A(n768), .S(n806), .Y(n766) );
  MUX2X1 U721 ( .B(n770), .A(n771), .S(n806), .Y(n769) );
  MUX2X1 U722 ( .B(n773), .A(n774), .S(n807), .Y(n772) );
  MUX2X1 U723 ( .B(n776), .A(n777), .S(n806), .Y(n775) );
  MUX2X1 U724 ( .B(n779), .A(n780), .S(n801), .Y(n778) );
  MUX2X1 U725 ( .B(n782), .A(n2), .S(n807), .Y(n781) );
  MUX2X1 U726 ( .B(n784), .A(n785), .S(n808), .Y(n783) );
  MUX2X1 U727 ( .B(n787), .A(n788), .S(n807), .Y(n786) );
  MUX2X1 U728 ( .B(n790), .A(n791), .S(n808), .Y(n789) );
  MUX2X1 U729 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n819), .Y(n649) );
  MUX2X1 U730 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n819), .Y(n648) );
  MUX2X1 U731 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n819), .Y(n652) );
  MUX2X1 U732 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n819), .Y(n651) );
  MUX2X1 U733 ( .B(n650), .A(n647), .S(n803), .Y(n661) );
  MUX2X1 U734 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n819), .Y(n655) );
  MUX2X1 U735 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n819), .Y(n654) );
  MUX2X1 U736 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n819), .Y(n658) );
  MUX2X1 U737 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n819), .Y(n657) );
  MUX2X1 U738 ( .B(n656), .A(n653), .S(n803), .Y(n660) );
  MUX2X1 U739 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n819), .Y(n664) );
  MUX2X1 U740 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n819), .Y(n663) );
  MUX2X1 U741 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n819), .Y(n667) );
  MUX2X1 U742 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n819), .Y(n666) );
  MUX2X1 U743 ( .B(n665), .A(n662), .S(n803), .Y(n676) );
  MUX2X1 U744 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n818), .Y(n670) );
  MUX2X1 U745 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n818), .Y(n669) );
  MUX2X1 U746 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n816), .Y(n673) );
  MUX2X1 U747 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n818), .Y(n672) );
  MUX2X1 U748 ( .B(n671), .A(n668), .S(n803), .Y(n675) );
  MUX2X1 U749 ( .B(n674), .A(n659), .S(n841), .Y(n795) );
  MUX2X1 U750 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n817), .Y(n679) );
  MUX2X1 U751 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n817), .Y(n678) );
  MUX2X1 U752 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n817), .Y(n682) );
  MUX2X1 U753 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n817), .Y(n681) );
  MUX2X1 U754 ( .B(n680), .A(n677), .S(n803), .Y(n691) );
  MUX2X1 U755 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n818), .Y(n685) );
  MUX2X1 U756 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n816), .Y(n684) );
  MUX2X1 U757 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n818), .Y(n688) );
  MUX2X1 U758 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n817), .Y(n687) );
  MUX2X1 U759 ( .B(n686), .A(n683), .S(n803), .Y(n690) );
  MUX2X1 U760 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n818), .Y(n694) );
  MUX2X1 U761 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n817), .Y(n693) );
  MUX2X1 U762 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n816), .Y(n696) );
  MUX2X1 U763 ( .B(n695), .A(n692), .S(n803), .Y(n706) );
  MUX2X1 U764 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n818), .Y(n700) );
  MUX2X1 U765 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n818), .Y(n699) );
  MUX2X1 U766 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n816), .Y(n703) );
  MUX2X1 U767 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n816), .Y(n702) );
  MUX2X1 U768 ( .B(n701), .A(n698), .S(n803), .Y(n705) );
  MUX2X1 U769 ( .B(n704), .A(n689), .S(n841), .Y(n796) );
  MUX2X1 U770 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n817), .Y(n709) );
  MUX2X1 U771 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n817), .Y(n708) );
  MUX2X1 U772 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n817), .Y(n712) );
  MUX2X1 U773 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n817), .Y(n711) );
  MUX2X1 U774 ( .B(n710), .A(n707), .S(n803), .Y(n721) );
  MUX2X1 U775 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n818), .Y(n715) );
  MUX2X1 U776 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n817), .Y(n714) );
  MUX2X1 U777 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n818), .Y(n718) );
  MUX2X1 U778 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n818), .Y(n717) );
  MUX2X1 U779 ( .B(n716), .A(n713), .S(n803), .Y(n720) );
  MUX2X1 U780 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n818), .Y(n724) );
  MUX2X1 U781 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n817), .Y(n723) );
  MUX2X1 U782 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n816), .Y(n727) );
  MUX2X1 U783 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n816), .Y(n726) );
  MUX2X1 U784 ( .B(n725), .A(n722), .S(n803), .Y(n736) );
  MUX2X1 U785 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n818), .Y(n730) );
  MUX2X1 U786 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n817), .Y(n729) );
  MUX2X1 U787 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n816), .Y(n733) );
  MUX2X1 U788 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n820), .Y(n732) );
  MUX2X1 U789 ( .B(n731), .A(n728), .S(n803), .Y(n735) );
  MUX2X1 U790 ( .B(n734), .A(n719), .S(n841), .Y(n797) );
  MUX2X1 U791 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n814), .Y(n739) );
  MUX2X1 U792 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n814), .Y(n738) );
  MUX2X1 U793 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n814), .Y(n742) );
  MUX2X1 U794 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n814), .Y(n741) );
  MUX2X1 U795 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n815), .Y(n745) );
  MUX2X1 U796 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n815), .Y(n744) );
  MUX2X1 U797 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n814), .Y(n748) );
  MUX2X1 U798 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n814), .Y(n747) );
  MUX2X1 U799 ( .B(n746), .A(n743), .S(n802), .Y(n750) );
  MUX2X1 U800 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n813), .Y(n753) );
  MUX2X1 U801 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n815), .Y(n756) );
  MUX2X1 U802 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n814), .Y(n759) );
  MUX2X1 U803 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n815), .Y(n758) );
  MUX2X1 U804 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n813), .Y(n762) );
  MUX2X1 U805 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n815), .Y(n761) );
  MUX2X1 U806 ( .B(n760), .A(n757), .S(n802), .Y(n764) );
  MUX2X1 U807 ( .B(n763), .A(n749), .S(n841), .Y(n798) );
  MUX2X1 U808 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n815), .Y(n768) );
  MUX2X1 U809 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n814), .Y(n767) );
  MUX2X1 U810 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n814), .Y(n771) );
  MUX2X1 U811 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n815), .Y(n770) );
  MUX2X1 U812 ( .B(n769), .A(n766), .S(n802), .Y(n780) );
  MUX2X1 U813 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n815), .Y(n774) );
  MUX2X1 U814 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n815), .Y(n773) );
  MUX2X1 U815 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n815), .Y(n777) );
  MUX2X1 U816 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n815), .Y(n776) );
  MUX2X1 U817 ( .B(n775), .A(n772), .S(n802), .Y(n779) );
  MUX2X1 U818 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n813), .Y(n782) );
  MUX2X1 U819 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n814), .Y(n785) );
  MUX2X1 U820 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n814), .Y(n784) );
  MUX2X1 U821 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n814), .Y(n788) );
  MUX2X1 U822 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n815), .Y(n787) );
  MUX2X1 U823 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n813), .Y(n791) );
  MUX2X1 U824 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n813), .Y(n790) );
  MUX2X1 U825 ( .B(n789), .A(n786), .S(n802), .Y(n793) );
  MUX2X1 U826 ( .B(n792), .A(n778), .S(n841), .Y(n799) );
  INVX8 U827 ( .A(N13), .Y(n800) );
  INVX8 U828 ( .A(n800), .Y(n801) );
  INVX8 U829 ( .A(n839), .Y(n803) );
  INVX8 U830 ( .A(n836), .Y(n805) );
  INVX8 U831 ( .A(n805), .Y(n806) );
  INVX8 U832 ( .A(n805), .Y(n807) );
  INVX8 U833 ( .A(n804), .Y(n809) );
  INVX8 U834 ( .A(n834), .Y(n811) );
  INVX8 U835 ( .A(n834), .Y(n812) );
  INVX8 U836 ( .A(n812), .Y(n813) );
  INVX8 U837 ( .A(n812), .Y(n814) );
  INVX8 U838 ( .A(n812), .Y(n815) );
  INVX8 U839 ( .A(n811), .Y(n816) );
  INVX8 U840 ( .A(n811), .Y(n817) );
  INVX8 U841 ( .A(n811), .Y(n818) );
  INVX8 U842 ( .A(n810), .Y(n819) );
  INVX1 U843 ( .A(n798), .Y(N18) );
  INVX1 U844 ( .A(n810), .Y(n820) );
  INVX1 U845 ( .A(n797), .Y(N19) );
  INVX1 U846 ( .A(n799), .Y(N17) );
  INVX2 U847 ( .A(N10), .Y(n835) );
  INVX1 U848 ( .A(n499), .Y(n821) );
  INVX1 U849 ( .A(n821), .Y(n822) );
  INVX8 U850 ( .A(n837), .Y(n836) );
  INVX8 U851 ( .A(n842), .Y(n841) );
  INVX8 U852 ( .A(N14), .Y(n842) );
  AND2X2 U853 ( .A(n509), .B(N21), .Y(\data_out<0> ) );
  AND2X2 U854 ( .A(N20), .B(n502), .Y(\data_out<1> ) );
  AND2X2 U855 ( .A(N19), .B(n502), .Y(\data_out<2> ) );
  AND2X2 U856 ( .A(N18), .B(n508), .Y(\data_out<3> ) );
  AND2X2 U857 ( .A(N17), .B(n503), .Y(\data_out<4> ) );
endmodule


module memc_Size1_0 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , N17, n1, n2,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n216), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n217), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n218), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n219), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n220), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n221), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n222), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n223), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n224), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n225), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n226), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n227), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n228), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n229), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n230), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n231), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n232), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n233), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n234), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n235), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n236), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n237), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n238), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n239), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n240), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n241), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n242), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n243), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n244), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n245), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n246), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n247), .CLK(clk), .Q(\mem<31><0> ) );
  INVX1 U2 ( .A(n172), .Y(n171) );
  INVX1 U3 ( .A(N13), .Y(n170) );
  INVX1 U4 ( .A(n158), .Y(N17) );
  INVX1 U5 ( .A(rst), .Y(n163) );
  AND2X1 U6 ( .A(n171), .B(n169), .Y(n174) );
  INVX1 U7 ( .A(n166), .Y(n159) );
  AND2X1 U8 ( .A(n165), .B(n60), .Y(n115) );
  INVX1 U9 ( .A(n164), .Y(n160) );
  NOR3X1 U10 ( .A(n170), .B(n56), .C(N14), .Y(n1) );
  INVX1 U11 ( .A(n170), .Y(n169) );
  INVX1 U12 ( .A(N14), .Y(n172) );
  OR2X2 U13 ( .A(n94), .B(write), .Y(n2) );
  INVX1 U14 ( .A(n2), .Y(\data_out<0> ) );
  AND2X2 U15 ( .A(n117), .B(n53), .Y(n4) );
  INVX1 U16 ( .A(n4), .Y(n5) );
  AND2X2 U17 ( .A(n113), .B(n53), .Y(n6) );
  INVX1 U18 ( .A(n6), .Y(n7) );
  AND2X2 U19 ( .A(n102), .B(n53), .Y(n8) );
  INVX1 U20 ( .A(n8), .Y(n9) );
  AND2X2 U21 ( .A(n104), .B(n53), .Y(n10) );
  INVX1 U22 ( .A(n10), .Y(n11) );
  AND2X2 U23 ( .A(n106), .B(n53), .Y(n12) );
  INVX1 U24 ( .A(n12), .Y(n13) );
  AND2X2 U25 ( .A(n108), .B(n53), .Y(n14) );
  INVX1 U26 ( .A(n14), .Y(n15) );
  AND2X2 U27 ( .A(n110), .B(n53), .Y(n16) );
  INVX1 U28 ( .A(n16), .Y(n17) );
  AND2X2 U29 ( .A(n115), .B(n53), .Y(n18) );
  INVX1 U30 ( .A(n18), .Y(n19) );
  AND2X2 U31 ( .A(n117), .B(n54), .Y(n20) );
  INVX1 U32 ( .A(n20), .Y(n21) );
  AND2X2 U33 ( .A(n113), .B(n54), .Y(n22) );
  INVX1 U34 ( .A(n22), .Y(n23) );
  AND2X2 U35 ( .A(n102), .B(n54), .Y(n24) );
  INVX1 U36 ( .A(n24), .Y(n25) );
  AND2X2 U37 ( .A(n104), .B(n54), .Y(n26) );
  INVX1 U38 ( .A(n26), .Y(n27) );
  AND2X2 U39 ( .A(n106), .B(n54), .Y(n28) );
  INVX1 U40 ( .A(n28), .Y(n29) );
  AND2X2 U41 ( .A(n108), .B(n54), .Y(n30) );
  INVX1 U42 ( .A(n30), .Y(n31) );
  AND2X2 U43 ( .A(n110), .B(n54), .Y(n32) );
  INVX1 U44 ( .A(n32), .Y(n33) );
  AND2X2 U45 ( .A(n115), .B(n54), .Y(n34) );
  INVX1 U46 ( .A(n34), .Y(n35) );
  AND2X2 U47 ( .A(n117), .B(n55), .Y(n36) );
  INVX1 U48 ( .A(n36), .Y(n37) );
  AND2X2 U49 ( .A(n113), .B(n55), .Y(n38) );
  INVX1 U50 ( .A(n38), .Y(n39) );
  AND2X2 U51 ( .A(n102), .B(n55), .Y(n40) );
  INVX1 U52 ( .A(n40), .Y(n41) );
  AND2X2 U53 ( .A(n104), .B(n55), .Y(n42) );
  INVX1 U54 ( .A(n42), .Y(n43) );
  AND2X2 U55 ( .A(n106), .B(n55), .Y(n44) );
  INVX1 U56 ( .A(n44), .Y(n45) );
  AND2X2 U57 ( .A(n108), .B(n55), .Y(n46) );
  INVX1 U58 ( .A(n46), .Y(n47) );
  AND2X2 U59 ( .A(n110), .B(n55), .Y(n48) );
  INVX1 U60 ( .A(n48), .Y(n49) );
  AND2X2 U61 ( .A(n115), .B(n55), .Y(n50) );
  INVX1 U62 ( .A(n50), .Y(n51) );
  BUFX2 U63 ( .A(n173), .Y(n52) );
  AND2X2 U64 ( .A(\data_in<0> ), .B(n98), .Y(n53) );
  AND2X2 U65 ( .A(\data_in<0> ), .B(n193), .Y(n54) );
  AND2X2 U66 ( .A(\data_in<0> ), .B(n123), .Y(n55) );
  OR2X2 U67 ( .A(n52), .B(\addr<5> ), .Y(n56) );
  INVX1 U68 ( .A(n56), .Y(n57) );
  INVX1 U69 ( .A(n56), .Y(n58) );
  INVX2 U70 ( .A(n123), .Y(n101) );
  INVX1 U71 ( .A(n165), .Y(n164) );
  INVX1 U72 ( .A(n168), .Y(n167) );
  OR2X1 U73 ( .A(n159), .B(n167), .Y(n59) );
  INVX1 U74 ( .A(n59), .Y(n60) );
  AND2X1 U75 ( .A(N17), .B(n163), .Y(n93) );
  INVX1 U76 ( .A(n93), .Y(n94) );
  AND2X1 U77 ( .A(n167), .B(n159), .Y(n95) );
  INVX1 U78 ( .A(n100), .Y(n193) );
  OR2X1 U79 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n96) );
  INVX1 U80 ( .A(n96), .Y(n97) );
  INVX1 U81 ( .A(n191), .Y(n98) );
  INVX1 U82 ( .A(n98), .Y(n99) );
  INVX1 U83 ( .A(n1), .Y(n100) );
  INVX1 U84 ( .A(n103), .Y(n102) );
  BUFX2 U85 ( .A(n204), .Y(n103) );
  INVX1 U86 ( .A(n105), .Y(n104) );
  BUFX2 U87 ( .A(n206), .Y(n105) );
  INVX1 U88 ( .A(n107), .Y(n106) );
  BUFX2 U89 ( .A(n208), .Y(n107) );
  INVX1 U90 ( .A(n109), .Y(n108) );
  BUFX2 U91 ( .A(n210), .Y(n109) );
  INVX1 U92 ( .A(n111), .Y(n110) );
  BUFX2 U93 ( .A(n212), .Y(n111) );
  INVX1 U94 ( .A(n113), .Y(n112) );
  AND2X1 U95 ( .A(n165), .B(n95), .Y(n113) );
  INVX1 U96 ( .A(n115), .Y(n114) );
  INVX1 U97 ( .A(n117), .Y(n116) );
  AND2X1 U98 ( .A(n164), .B(n95), .Y(n117) );
  INVX1 U99 ( .A(n122), .Y(n118) );
  INVX1 U100 ( .A(n122), .Y(n119) );
  INVX1 U101 ( .A(n122), .Y(n120) );
  INVX1 U102 ( .A(n122), .Y(n121) );
  AND2X2 U103 ( .A(\data_in<0> ), .B(n162), .Y(n122) );
  INVX1 U104 ( .A(n214), .Y(n123) );
  BUFX2 U105 ( .A(n100), .Y(n124) );
  BUFX2 U106 ( .A(n100), .Y(n125) );
  BUFX2 U107 ( .A(n99), .Y(n126) );
  BUFX2 U108 ( .A(n99), .Y(n127) );
  INVX1 U109 ( .A(N12), .Y(n168) );
  MUX2X1 U110 ( .B(n129), .A(n130), .S(n159), .Y(n128) );
  MUX2X1 U111 ( .B(n132), .A(n133), .S(n159), .Y(n131) );
  MUX2X1 U112 ( .B(n135), .A(n136), .S(n159), .Y(n134) );
  MUX2X1 U113 ( .B(n138), .A(n139), .S(n159), .Y(n137) );
  MUX2X1 U114 ( .B(n141), .A(n142), .S(n169), .Y(n140) );
  MUX2X1 U115 ( .B(n144), .A(n145), .S(n159), .Y(n143) );
  MUX2X1 U116 ( .B(n147), .A(n148), .S(n159), .Y(n146) );
  MUX2X1 U117 ( .B(n150), .A(n151), .S(n159), .Y(n149) );
  MUX2X1 U118 ( .B(n153), .A(n154), .S(n159), .Y(n152) );
  MUX2X1 U119 ( .B(n156), .A(n157), .S(n169), .Y(n155) );
  MUX2X1 U120 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n161), .Y(n130) );
  MUX2X1 U121 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n161), .Y(n129) );
  MUX2X1 U122 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n161), .Y(n133) );
  MUX2X1 U123 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n161), .Y(n132) );
  MUX2X1 U124 ( .B(n131), .A(n128), .S(n167), .Y(n142) );
  MUX2X1 U125 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n161), .Y(n136) );
  MUX2X1 U126 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n161), .Y(n135) );
  MUX2X1 U127 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n161), .Y(n139) );
  MUX2X1 U128 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n161), .Y(n138) );
  MUX2X1 U129 ( .B(n137), .A(n134), .S(n167), .Y(n141) );
  MUX2X1 U130 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n161), .Y(n145) );
  MUX2X1 U131 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n161), .Y(n144) );
  MUX2X1 U132 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n161), .Y(n148) );
  MUX2X1 U133 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n161), .Y(n147) );
  MUX2X1 U134 ( .B(n146), .A(n143), .S(n167), .Y(n157) );
  MUX2X1 U135 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n161), .Y(n151) );
  MUX2X1 U136 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n161), .Y(n150) );
  MUX2X1 U137 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n161), .Y(n154) );
  MUX2X1 U138 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n161), .Y(n153) );
  MUX2X1 U139 ( .B(n152), .A(n149), .S(n167), .Y(n156) );
  MUX2X1 U140 ( .B(n155), .A(n140), .S(n171), .Y(n158) );
  INVX8 U141 ( .A(n160), .Y(n161) );
  AND2X2 U142 ( .A(n58), .B(n174), .Y(n162) );
  INVX4 U143 ( .A(n162), .Y(n182) );
  INVX1 U144 ( .A(N11), .Y(n166) );
  INVX1 U145 ( .A(N10), .Y(n165) );
  NAND3X1 U146 ( .A(write), .B(n163), .C(n97), .Y(n173) );
  OAI21X1 U147 ( .A(n182), .B(n116), .C(\mem<31><0> ), .Y(n175) );
  OAI21X1 U148 ( .A(n118), .B(n116), .C(n175), .Y(n247) );
  OAI21X1 U149 ( .A(n112), .B(n182), .C(\mem<30><0> ), .Y(n176) );
  OAI21X1 U150 ( .A(n112), .B(n121), .C(n176), .Y(n246) );
  NAND3X1 U151 ( .A(n164), .B(n167), .C(n166), .Y(n204) );
  OAI21X1 U152 ( .A(n103), .B(n182), .C(\mem<29><0> ), .Y(n177) );
  OAI21X1 U153 ( .A(n103), .B(n119), .C(n177), .Y(n245) );
  NAND3X1 U154 ( .A(n167), .B(n166), .C(n165), .Y(n206) );
  OAI21X1 U155 ( .A(n105), .B(n182), .C(\mem<28><0> ), .Y(n178) );
  OAI21X1 U156 ( .A(n105), .B(n120), .C(n178), .Y(n244) );
  NAND3X1 U157 ( .A(n164), .B(n159), .C(n168), .Y(n208) );
  OAI21X1 U158 ( .A(n107), .B(n182), .C(\mem<27><0> ), .Y(n179) );
  OAI21X1 U159 ( .A(n107), .B(n120), .C(n179), .Y(n243) );
  NAND3X1 U160 ( .A(n168), .B(n159), .C(n165), .Y(n210) );
  OAI21X1 U161 ( .A(n109), .B(n182), .C(\mem<26><0> ), .Y(n180) );
  OAI21X1 U162 ( .A(n109), .B(n121), .C(n180), .Y(n242) );
  NAND3X1 U163 ( .A(n164), .B(n168), .C(n166), .Y(n212) );
  OAI21X1 U164 ( .A(n111), .B(n182), .C(\mem<25><0> ), .Y(n181) );
  OAI21X1 U165 ( .A(n111), .B(n119), .C(n181), .Y(n241) );
  OAI21X1 U166 ( .A(n114), .B(n182), .C(\mem<24><0> ), .Y(n183) );
  OAI21X1 U167 ( .A(n114), .B(n118), .C(n183), .Y(n240) );
  NAND3X1 U168 ( .A(n171), .B(n170), .C(n58), .Y(n191) );
  OAI21X1 U169 ( .A(n127), .B(n116), .C(\mem<23><0> ), .Y(n184) );
  NAND2X1 U170 ( .A(n5), .B(n184), .Y(n239) );
  OAI21X1 U171 ( .A(n126), .B(n112), .C(\mem<22><0> ), .Y(n185) );
  NAND2X1 U172 ( .A(n7), .B(n185), .Y(n238) );
  OAI21X1 U173 ( .A(n127), .B(n103), .C(\mem<21><0> ), .Y(n186) );
  NAND2X1 U174 ( .A(n9), .B(n186), .Y(n237) );
  OAI21X1 U175 ( .A(n126), .B(n105), .C(\mem<20><0> ), .Y(n187) );
  NAND2X1 U176 ( .A(n11), .B(n187), .Y(n236) );
  OAI21X1 U177 ( .A(n127), .B(n107), .C(\mem<19><0> ), .Y(n188) );
  NAND2X1 U178 ( .A(n13), .B(n188), .Y(n235) );
  OAI21X1 U179 ( .A(n126), .B(n109), .C(\mem<18><0> ), .Y(n189) );
  NAND2X1 U180 ( .A(n15), .B(n189), .Y(n234) );
  OAI21X1 U181 ( .A(n127), .B(n111), .C(\mem<17><0> ), .Y(n190) );
  NAND2X1 U182 ( .A(n17), .B(n190), .Y(n233) );
  OAI21X1 U183 ( .A(n126), .B(n114), .C(\mem<16><0> ), .Y(n192) );
  NAND2X1 U184 ( .A(n19), .B(n192), .Y(n232) );
  OAI21X1 U185 ( .A(n125), .B(n116), .C(\mem<15><0> ), .Y(n194) );
  NAND2X1 U186 ( .A(n21), .B(n194), .Y(n231) );
  OAI21X1 U187 ( .A(n124), .B(n112), .C(\mem<14><0> ), .Y(n195) );
  NAND2X1 U188 ( .A(n23), .B(n195), .Y(n230) );
  OAI21X1 U189 ( .A(n125), .B(n103), .C(\mem<13><0> ), .Y(n196) );
  NAND2X1 U190 ( .A(n25), .B(n196), .Y(n229) );
  OAI21X1 U191 ( .A(n124), .B(n105), .C(\mem<12><0> ), .Y(n197) );
  NAND2X1 U192 ( .A(n27), .B(n197), .Y(n228) );
  OAI21X1 U193 ( .A(n125), .B(n107), .C(\mem<11><0> ), .Y(n198) );
  NAND2X1 U194 ( .A(n29), .B(n198), .Y(n227) );
  OAI21X1 U195 ( .A(n124), .B(n109), .C(\mem<10><0> ), .Y(n199) );
  NAND2X1 U196 ( .A(n31), .B(n199), .Y(n226) );
  OAI21X1 U197 ( .A(n125), .B(n111), .C(\mem<9><0> ), .Y(n200) );
  NAND2X1 U198 ( .A(n33), .B(n200), .Y(n225) );
  OAI21X1 U199 ( .A(n124), .B(n114), .C(\mem<8><0> ), .Y(n201) );
  NAND2X1 U200 ( .A(n35), .B(n201), .Y(n224) );
  NAND3X1 U201 ( .A(n57), .B(n170), .C(n172), .Y(n214) );
  OAI21X1 U202 ( .A(n101), .B(n116), .C(\mem<7><0> ), .Y(n202) );
  NAND2X1 U203 ( .A(n37), .B(n202), .Y(n223) );
  OAI21X1 U204 ( .A(n101), .B(n112), .C(\mem<6><0> ), .Y(n203) );
  NAND2X1 U205 ( .A(n39), .B(n203), .Y(n222) );
  OAI21X1 U206 ( .A(n101), .B(n103), .C(\mem<5><0> ), .Y(n205) );
  NAND2X1 U207 ( .A(n41), .B(n205), .Y(n221) );
  OAI21X1 U208 ( .A(n101), .B(n105), .C(\mem<4><0> ), .Y(n207) );
  NAND2X1 U209 ( .A(n43), .B(n207), .Y(n220) );
  OAI21X1 U210 ( .A(n101), .B(n107), .C(\mem<3><0> ), .Y(n209) );
  NAND2X1 U211 ( .A(n45), .B(n209), .Y(n219) );
  OAI21X1 U212 ( .A(n101), .B(n109), .C(\mem<2><0> ), .Y(n211) );
  NAND2X1 U213 ( .A(n47), .B(n211), .Y(n218) );
  OAI21X1 U214 ( .A(n101), .B(n111), .C(\mem<1><0> ), .Y(n213) );
  NAND2X1 U215 ( .A(n49), .B(n213), .Y(n217) );
  OAI21X1 U216 ( .A(n101), .B(n114), .C(\mem<0><0> ), .Y(n215) );
  NAND2X1 U217 ( .A(n51), .B(n215), .Y(n216) );
endmodule


module memv_0 ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , N28, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n41,
         n43, n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60, n62,
         n63, n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81, n83,
         n84, n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149,
         n150, n152, n169, n171, n187, n189, n205, n207, n223, n225, n241,
         n242, n244, n260, n262, n278, n280, n296, n298, n314, n315, n317,
         n333, n335, n351, n353, n354, n360, n362, n369, n374, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n1019), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n1020), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n1021), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n1022), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n1023), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n1024), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n1025), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n1026), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n1027), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n1028), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n1029), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n1030), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n1031), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n1032), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n1033), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n1034), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n1035), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n1036), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n1037), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n1038), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n1039), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n1040), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n1041), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n1042), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n1043), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n1044), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n1045), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n1046), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n1047), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n1048), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n1049), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n1050), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n1051), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n1052), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n1053), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n1054), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n1055), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n1056), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n1057), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n1058), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n1059), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n1060), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n1061), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n1062), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n1063), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n1064), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n1065), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n1066), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n1067), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n1068), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n1069), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n1070), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n1071), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n1072), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n1073), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n1074), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n1075), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n1076), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n1077), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n1078), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n1079), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n1080), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n1081), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n1082), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n1083), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n1084), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n1085), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n1086), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n1087), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n1088), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n1089), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n1090), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n1091), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n1092), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n1093), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n1094), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n1095), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n1096), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n1097), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n1098), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n1099), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n1100), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n1101), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n1102), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n1103), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n1104), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n1105), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n1106), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n1107), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n1108), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n1109), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n1110), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n1111), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n1112), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n1113), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n1114), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n1115), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n1116), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n1117), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n1118), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n1119), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n1120), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n1121), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n1122), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n1123), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n1124), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n1125), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n1126), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n1127), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n1128), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n1129), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n1130), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n1131), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n1132), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n1133), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n1134), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n1135), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n1136), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n1137), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n1138), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n1139), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n1140), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n1141), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n1142), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n1143), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n1144), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n1145), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n1146), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n1147), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n1148), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n1149), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n1150), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n1151), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n1152), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n1153), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n1154), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n1155), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n1156), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n1157), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n1158), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n1159), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n1160), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n1161), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n1162), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n1163), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n1164), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n1165), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n1166), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n1167), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n1168), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n1169), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n1170), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n1171), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n1172), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n1173), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n1174), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n1175), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n1176), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n1177), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n1178), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n1179), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n1180), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n1181), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n1182), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n1183), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n1184), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n1185), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n1186), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n1187), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n1188), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n1189), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n1190), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n1191), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n1192), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n1193), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n1194), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n1195), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n1196), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n1197), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n1198), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n1199), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n1200), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n1201), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n1202), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n1203), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n1204), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n1205), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n1206), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n1207), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n1208), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n1209), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n1210), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n1211), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n1212), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n1213), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n1214), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n1215), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n1216), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n1217), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n1218), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n1219), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n1220), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n1221), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n1222), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n1223), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n1224), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n1225), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n1226), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n1227), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n1228), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n1229), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n1230), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n1231), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n1232), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n1233), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n1234), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n1235), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n1236), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n1237), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n1238), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n1239), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n1240), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n1241), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n1242), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n1243), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n1244), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n1245), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n1246), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n1247), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n1248), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n1249), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n1250), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n1251), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n1252), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n1253), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n1254), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n1255), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n1256), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n1257), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n1258), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n1259), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n1260), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n1261), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n1262), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n1263), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n1264), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n1265), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n1266), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n1267), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n1268), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n1269), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n1270), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n1271), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n1272), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n1273), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n1274), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U4 ( .A(N23), .B(n1016), .Y(n1521) );
  AND2X2 U5 ( .A(N23), .B(n1017), .Y(n1504) );
  AND2X2 U6 ( .A(N21), .B(n1014), .Y(n1293) );
  AND2X2 U7 ( .A(N21), .B(n1015), .Y(n1286) );
  AND2X2 U8 ( .A(n1012), .B(n954), .Y(n1292) );
  AND2X2 U9 ( .A(n1012), .B(n673), .Y(n1290) );
  OAI21X1 U49 ( .A(n982), .B(n653), .C(n1539), .Y(n1274) );
  OAI21X1 U50 ( .A(n60), .B(n1009), .C(\mem<255> ), .Y(n1539) );
  OAI21X1 U51 ( .A(n653), .B(n979), .C(n1538), .Y(n1273) );
  OAI21X1 U52 ( .A(n1010), .B(n57), .C(\mem<254> ), .Y(n1538) );
  OAI21X1 U53 ( .A(n653), .B(n978), .C(n1537), .Y(n1272) );
  OAI21X1 U54 ( .A(n1010), .B(n54), .C(\mem<253> ), .Y(n1537) );
  OAI21X1 U55 ( .A(n653), .B(n977), .C(n1536), .Y(n1271) );
  OAI21X1 U56 ( .A(n1010), .B(n51), .C(\mem<252> ), .Y(n1536) );
  OAI21X1 U57 ( .A(n653), .B(n975), .C(n1535), .Y(n1270) );
  OAI21X1 U58 ( .A(n1010), .B(n48), .C(\mem<251> ), .Y(n1535) );
  OAI21X1 U59 ( .A(n653), .B(n973), .C(n1534), .Y(n1269) );
  OAI21X1 U60 ( .A(n1010), .B(n45), .C(\mem<250> ), .Y(n1534) );
  OAI21X1 U61 ( .A(n653), .B(n971), .C(n1533), .Y(n1268) );
  OAI21X1 U62 ( .A(n1010), .B(n43), .C(\mem<249> ), .Y(n1533) );
  OAI21X1 U63 ( .A(n653), .B(n969), .C(n1532), .Y(n1267) );
  OAI21X1 U64 ( .A(n1010), .B(n40), .C(\mem<248> ), .Y(n1532) );
  OAI21X1 U65 ( .A(n653), .B(n968), .C(n1531), .Y(n1266) );
  OAI21X1 U66 ( .A(n1010), .B(n37), .C(\mem<247> ), .Y(n1531) );
  OAI21X1 U67 ( .A(n653), .B(n967), .C(n1530), .Y(n1265) );
  OAI21X1 U68 ( .A(n1009), .B(n35), .C(\mem<246> ), .Y(n1530) );
  OAI21X1 U69 ( .A(n653), .B(n966), .C(n1529), .Y(n1264) );
  OAI21X1 U70 ( .A(n1009), .B(n33), .C(\mem<245> ), .Y(n1529) );
  OAI21X1 U71 ( .A(n653), .B(n965), .C(n1528), .Y(n1263) );
  OAI21X1 U72 ( .A(n1009), .B(n31), .C(\mem<244> ), .Y(n1528) );
  OAI21X1 U73 ( .A(n653), .B(n964), .C(n1527), .Y(n1262) );
  OAI21X1 U74 ( .A(n1009), .B(n29), .C(\mem<243> ), .Y(n1527) );
  OAI21X1 U75 ( .A(n653), .B(n963), .C(n1526), .Y(n1261) );
  OAI21X1 U76 ( .A(n1009), .B(n27), .C(\mem<242> ), .Y(n1526) );
  OAI21X1 U77 ( .A(n653), .B(n962), .C(n1525), .Y(n1260) );
  OAI21X1 U78 ( .A(n1009), .B(n25), .C(\mem<241> ), .Y(n1525) );
  OAI21X1 U79 ( .A(n653), .B(n959), .C(n1524), .Y(n1259) );
  OAI21X1 U80 ( .A(n1009), .B(n23), .C(\mem<240> ), .Y(n1524) );
  OAI21X1 U83 ( .A(n982), .B(n649), .C(n1520), .Y(n1258) );
  OAI21X1 U84 ( .A(n60), .B(n1008), .C(\mem<239> ), .Y(n1520) );
  OAI21X1 U85 ( .A(n980), .B(n649), .C(n1519), .Y(n1257) );
  OAI21X1 U86 ( .A(n57), .B(n1008), .C(\mem<238> ), .Y(n1519) );
  OAI21X1 U87 ( .A(n978), .B(n649), .C(n1518), .Y(n1256) );
  OAI21X1 U88 ( .A(n54), .B(n1008), .C(\mem<237> ), .Y(n1518) );
  OAI21X1 U89 ( .A(n977), .B(n649), .C(n1517), .Y(n1255) );
  OAI21X1 U90 ( .A(n51), .B(n1008), .C(\mem<236> ), .Y(n1517) );
  OAI21X1 U91 ( .A(n976), .B(n649), .C(n1516), .Y(n1254) );
  OAI21X1 U92 ( .A(n48), .B(n1008), .C(\mem<235> ), .Y(n1516) );
  OAI21X1 U93 ( .A(n974), .B(n649), .C(n1515), .Y(n1253) );
  OAI21X1 U94 ( .A(n45), .B(n1008), .C(\mem<234> ), .Y(n1515) );
  OAI21X1 U95 ( .A(n972), .B(n649), .C(n1514), .Y(n1252) );
  OAI21X1 U96 ( .A(n43), .B(n1008), .C(\mem<233> ), .Y(n1514) );
  OAI21X1 U97 ( .A(n970), .B(n649), .C(n1513), .Y(n1251) );
  OAI21X1 U98 ( .A(n40), .B(n1008), .C(\mem<232> ), .Y(n1513) );
  OAI21X1 U99 ( .A(n968), .B(n649), .C(n1512), .Y(n1250) );
  OAI21X1 U100 ( .A(n37), .B(n1007), .C(\mem<231> ), .Y(n1512) );
  OAI21X1 U101 ( .A(n967), .B(n649), .C(n1511), .Y(n1249) );
  OAI21X1 U102 ( .A(n35), .B(n1007), .C(\mem<230> ), .Y(n1511) );
  OAI21X1 U103 ( .A(n966), .B(n649), .C(n1510), .Y(n1248) );
  OAI21X1 U104 ( .A(n33), .B(n1007), .C(\mem<229> ), .Y(n1510) );
  OAI21X1 U105 ( .A(n965), .B(n649), .C(n1509), .Y(n1247) );
  OAI21X1 U106 ( .A(n31), .B(n1007), .C(\mem<228> ), .Y(n1509) );
  OAI21X1 U107 ( .A(n964), .B(n649), .C(n1508), .Y(n1246) );
  OAI21X1 U108 ( .A(n29), .B(n1007), .C(\mem<227> ), .Y(n1508) );
  OAI21X1 U109 ( .A(n963), .B(n649), .C(n1507), .Y(n1245) );
  OAI21X1 U110 ( .A(n27), .B(n1007), .C(\mem<226> ), .Y(n1507) );
  OAI21X1 U111 ( .A(n962), .B(n649), .C(n1506), .Y(n1244) );
  OAI21X1 U112 ( .A(n25), .B(n1007), .C(\mem<225> ), .Y(n1506) );
  OAI21X1 U113 ( .A(n959), .B(n649), .C(n1505), .Y(n1243) );
  OAI21X1 U114 ( .A(n23), .B(n1007), .C(\mem<224> ), .Y(n1505) );
  OAI21X1 U117 ( .A(n982), .B(n645), .C(n1503), .Y(n1242) );
  OAI21X1 U118 ( .A(n60), .B(n1006), .C(\mem<223> ), .Y(n1503) );
  OAI21X1 U119 ( .A(n980), .B(n645), .C(n1502), .Y(n1241) );
  OAI21X1 U120 ( .A(n57), .B(n1006), .C(\mem<222> ), .Y(n1502) );
  OAI21X1 U121 ( .A(n978), .B(n645), .C(n1501), .Y(n1240) );
  OAI21X1 U122 ( .A(n54), .B(n1006), .C(\mem<221> ), .Y(n1501) );
  OAI21X1 U123 ( .A(n977), .B(n645), .C(n1500), .Y(n1239) );
  OAI21X1 U124 ( .A(n51), .B(n1006), .C(\mem<220> ), .Y(n1500) );
  OAI21X1 U125 ( .A(n976), .B(n645), .C(n1499), .Y(n1238) );
  OAI21X1 U126 ( .A(n48), .B(n1006), .C(\mem<219> ), .Y(n1499) );
  OAI21X1 U127 ( .A(n974), .B(n645), .C(n1498), .Y(n1237) );
  OAI21X1 U128 ( .A(n45), .B(n1006), .C(\mem<218> ), .Y(n1498) );
  OAI21X1 U129 ( .A(n972), .B(n645), .C(n1497), .Y(n1236) );
  OAI21X1 U130 ( .A(n43), .B(n1006), .C(\mem<217> ), .Y(n1497) );
  OAI21X1 U131 ( .A(n970), .B(n645), .C(n1496), .Y(n1235) );
  OAI21X1 U132 ( .A(n40), .B(n1006), .C(\mem<216> ), .Y(n1496) );
  OAI21X1 U133 ( .A(n968), .B(n645), .C(n1495), .Y(n1234) );
  OAI21X1 U134 ( .A(n37), .B(n1006), .C(\mem<215> ), .Y(n1495) );
  OAI21X1 U135 ( .A(n967), .B(n645), .C(n1494), .Y(n1233) );
  OAI21X1 U136 ( .A(n35), .B(n1006), .C(\mem<214> ), .Y(n1494) );
  OAI21X1 U137 ( .A(n966), .B(n645), .C(n1493), .Y(n1232) );
  OAI21X1 U138 ( .A(n33), .B(n1006), .C(\mem<213> ), .Y(n1493) );
  OAI21X1 U139 ( .A(n965), .B(n645), .C(n1492), .Y(n1231) );
  OAI21X1 U140 ( .A(n31), .B(n1006), .C(\mem<212> ), .Y(n1492) );
  OAI21X1 U141 ( .A(n964), .B(n645), .C(n1491), .Y(n1230) );
  OAI21X1 U142 ( .A(n29), .B(n1006), .C(\mem<211> ), .Y(n1491) );
  OAI21X1 U143 ( .A(n963), .B(n645), .C(n1490), .Y(n1229) );
  OAI21X1 U144 ( .A(n27), .B(n1006), .C(\mem<210> ), .Y(n1490) );
  OAI21X1 U145 ( .A(n962), .B(n645), .C(n1489), .Y(n1228) );
  OAI21X1 U146 ( .A(n25), .B(n1006), .C(\mem<209> ), .Y(n1489) );
  OAI21X1 U147 ( .A(n959), .B(n645), .C(n1488), .Y(n1227) );
  OAI21X1 U148 ( .A(n23), .B(n1006), .C(\mem<208> ), .Y(n1488) );
  OAI21X1 U151 ( .A(n982), .B(n643), .C(n1487), .Y(n1226) );
  OAI21X1 U152 ( .A(n60), .B(n1005), .C(\mem<207> ), .Y(n1487) );
  OAI21X1 U153 ( .A(n980), .B(n643), .C(n1486), .Y(n1225) );
  OAI21X1 U154 ( .A(n57), .B(n1005), .C(\mem<206> ), .Y(n1486) );
  OAI21X1 U155 ( .A(n978), .B(n643), .C(n1485), .Y(n1224) );
  OAI21X1 U156 ( .A(n54), .B(n1005), .C(\mem<205> ), .Y(n1485) );
  OAI21X1 U157 ( .A(n977), .B(n643), .C(n1484), .Y(n1223) );
  OAI21X1 U158 ( .A(n51), .B(n1005), .C(\mem<204> ), .Y(n1484) );
  OAI21X1 U159 ( .A(n976), .B(n643), .C(n1483), .Y(n1222) );
  OAI21X1 U160 ( .A(n48), .B(n1005), .C(\mem<203> ), .Y(n1483) );
  OAI21X1 U161 ( .A(n974), .B(n643), .C(n1482), .Y(n1221) );
  OAI21X1 U162 ( .A(n45), .B(n1005), .C(\mem<202> ), .Y(n1482) );
  OAI21X1 U163 ( .A(n972), .B(n643), .C(n1481), .Y(n1220) );
  OAI21X1 U164 ( .A(n43), .B(n1005), .C(\mem<201> ), .Y(n1481) );
  OAI21X1 U165 ( .A(n970), .B(n643), .C(n1480), .Y(n1219) );
  OAI21X1 U166 ( .A(n40), .B(n1005), .C(\mem<200> ), .Y(n1480) );
  OAI21X1 U167 ( .A(n968), .B(n643), .C(n1479), .Y(n1218) );
  OAI21X1 U168 ( .A(n37), .B(n1005), .C(\mem<199> ), .Y(n1479) );
  OAI21X1 U169 ( .A(n967), .B(n643), .C(n1478), .Y(n1217) );
  OAI21X1 U170 ( .A(n35), .B(n1005), .C(\mem<198> ), .Y(n1478) );
  OAI21X1 U171 ( .A(n966), .B(n643), .C(n1477), .Y(n1216) );
  OAI21X1 U172 ( .A(n33), .B(n1005), .C(\mem<197> ), .Y(n1477) );
  OAI21X1 U173 ( .A(n965), .B(n643), .C(n1476), .Y(n1215) );
  OAI21X1 U174 ( .A(n31), .B(n1005), .C(\mem<196> ), .Y(n1476) );
  OAI21X1 U175 ( .A(n964), .B(n643), .C(n1475), .Y(n1214) );
  OAI21X1 U176 ( .A(n29), .B(n1005), .C(\mem<195> ), .Y(n1475) );
  OAI21X1 U177 ( .A(n963), .B(n643), .C(n1474), .Y(n1213) );
  OAI21X1 U178 ( .A(n27), .B(n1005), .C(\mem<194> ), .Y(n1474) );
  OAI21X1 U179 ( .A(n962), .B(n643), .C(n1473), .Y(n1212) );
  OAI21X1 U180 ( .A(n25), .B(n1005), .C(\mem<193> ), .Y(n1473) );
  OAI21X1 U181 ( .A(n959), .B(n643), .C(n1472), .Y(n1211) );
  OAI21X1 U182 ( .A(n23), .B(n1005), .C(\mem<192> ), .Y(n1472) );
  OAI21X1 U185 ( .A(n982), .B(n641), .C(n1471), .Y(n1210) );
  OAI21X1 U186 ( .A(n60), .B(n1004), .C(\mem<191> ), .Y(n1471) );
  OAI21X1 U187 ( .A(n980), .B(n641), .C(n1470), .Y(n1209) );
  OAI21X1 U188 ( .A(n57), .B(n1004), .C(\mem<190> ), .Y(n1470) );
  OAI21X1 U189 ( .A(n978), .B(n641), .C(n1469), .Y(n1208) );
  OAI21X1 U190 ( .A(n54), .B(n1004), .C(\mem<189> ), .Y(n1469) );
  OAI21X1 U191 ( .A(n977), .B(n641), .C(n1468), .Y(n1207) );
  OAI21X1 U192 ( .A(n51), .B(n1004), .C(\mem<188> ), .Y(n1468) );
  OAI21X1 U193 ( .A(n976), .B(n641), .C(n1467), .Y(n1206) );
  OAI21X1 U194 ( .A(n48), .B(n1004), .C(\mem<187> ), .Y(n1467) );
  OAI21X1 U195 ( .A(n974), .B(n641), .C(n1466), .Y(n1205) );
  OAI21X1 U196 ( .A(n45), .B(n1004), .C(\mem<186> ), .Y(n1466) );
  OAI21X1 U197 ( .A(n972), .B(n641), .C(n1465), .Y(n1204) );
  OAI21X1 U198 ( .A(n43), .B(n1004), .C(\mem<185> ), .Y(n1465) );
  OAI21X1 U199 ( .A(n970), .B(n641), .C(n1464), .Y(n1203) );
  OAI21X1 U200 ( .A(n40), .B(n1004), .C(\mem<184> ), .Y(n1464) );
  OAI21X1 U201 ( .A(n968), .B(n641), .C(n1463), .Y(n1202) );
  OAI21X1 U202 ( .A(n37), .B(n1003), .C(\mem<183> ), .Y(n1463) );
  OAI21X1 U203 ( .A(n967), .B(n641), .C(n1462), .Y(n1201) );
  OAI21X1 U204 ( .A(n35), .B(n1003), .C(\mem<182> ), .Y(n1462) );
  OAI21X1 U205 ( .A(n966), .B(n641), .C(n1461), .Y(n1200) );
  OAI21X1 U206 ( .A(n33), .B(n1003), .C(\mem<181> ), .Y(n1461) );
  OAI21X1 U207 ( .A(n965), .B(n641), .C(n1460), .Y(n1199) );
  OAI21X1 U208 ( .A(n31), .B(n1003), .C(\mem<180> ), .Y(n1460) );
  OAI21X1 U209 ( .A(n964), .B(n641), .C(n1459), .Y(n1198) );
  OAI21X1 U210 ( .A(n29), .B(n1003), .C(\mem<179> ), .Y(n1459) );
  OAI21X1 U211 ( .A(n963), .B(n641), .C(n1458), .Y(n1197) );
  OAI21X1 U212 ( .A(n27), .B(n1003), .C(\mem<178> ), .Y(n1458) );
  OAI21X1 U213 ( .A(n962), .B(n641), .C(n1457), .Y(n1196) );
  OAI21X1 U214 ( .A(n25), .B(n1003), .C(\mem<177> ), .Y(n1457) );
  OAI21X1 U215 ( .A(n959), .B(n641), .C(n1456), .Y(n1195) );
  OAI21X1 U216 ( .A(n23), .B(n1003), .C(\mem<176> ), .Y(n1456) );
  OAI21X1 U219 ( .A(n982), .B(n637), .C(n1454), .Y(n1194) );
  OAI21X1 U220 ( .A(n60), .B(n1002), .C(\mem<175> ), .Y(n1454) );
  OAI21X1 U221 ( .A(n980), .B(n637), .C(n1453), .Y(n1193) );
  OAI21X1 U222 ( .A(n57), .B(n1002), .C(\mem<174> ), .Y(n1453) );
  OAI21X1 U223 ( .A(n978), .B(n637), .C(n1452), .Y(n1192) );
  OAI21X1 U224 ( .A(n54), .B(n1002), .C(\mem<173> ), .Y(n1452) );
  OAI21X1 U225 ( .A(n977), .B(n637), .C(n1451), .Y(n1191) );
  OAI21X1 U226 ( .A(n51), .B(n1002), .C(\mem<172> ), .Y(n1451) );
  OAI21X1 U227 ( .A(n976), .B(n637), .C(n1450), .Y(n1190) );
  OAI21X1 U228 ( .A(n48), .B(n1002), .C(\mem<171> ), .Y(n1450) );
  OAI21X1 U229 ( .A(n974), .B(n637), .C(n1449), .Y(n1189) );
  OAI21X1 U230 ( .A(n45), .B(n1002), .C(\mem<170> ), .Y(n1449) );
  OAI21X1 U231 ( .A(n972), .B(n637), .C(n1448), .Y(n1188) );
  OAI21X1 U232 ( .A(n43), .B(n1002), .C(\mem<169> ), .Y(n1448) );
  OAI21X1 U233 ( .A(n970), .B(n637), .C(n1447), .Y(n1187) );
  OAI21X1 U234 ( .A(n40), .B(n1002), .C(\mem<168> ), .Y(n1447) );
  OAI21X1 U235 ( .A(n968), .B(n637), .C(n1446), .Y(n1186) );
  OAI21X1 U236 ( .A(n37), .B(n1001), .C(\mem<167> ), .Y(n1446) );
  OAI21X1 U237 ( .A(n967), .B(n637), .C(n1445), .Y(n1185) );
  OAI21X1 U238 ( .A(n35), .B(n1001), .C(\mem<166> ), .Y(n1445) );
  OAI21X1 U239 ( .A(n966), .B(n637), .C(n1444), .Y(n1184) );
  OAI21X1 U240 ( .A(n33), .B(n1001), .C(\mem<165> ), .Y(n1444) );
  OAI21X1 U241 ( .A(n965), .B(n637), .C(n1443), .Y(n1183) );
  OAI21X1 U242 ( .A(n31), .B(n1001), .C(\mem<164> ), .Y(n1443) );
  OAI21X1 U243 ( .A(n964), .B(n637), .C(n1442), .Y(n1182) );
  OAI21X1 U244 ( .A(n29), .B(n1001), .C(\mem<163> ), .Y(n1442) );
  OAI21X1 U245 ( .A(n963), .B(n637), .C(n1441), .Y(n1181) );
  OAI21X1 U246 ( .A(n27), .B(n1001), .C(\mem<162> ), .Y(n1441) );
  OAI21X1 U247 ( .A(n962), .B(n637), .C(n1440), .Y(n1180) );
  OAI21X1 U248 ( .A(n25), .B(n1001), .C(\mem<161> ), .Y(n1440) );
  OAI21X1 U249 ( .A(n959), .B(n637), .C(n1439), .Y(n1179) );
  OAI21X1 U250 ( .A(n23), .B(n1001), .C(\mem<160> ), .Y(n1439) );
  OAI21X1 U253 ( .A(n982), .B(n374), .C(n1438), .Y(n1178) );
  OAI21X1 U254 ( .A(n60), .B(n1000), .C(\mem<159> ), .Y(n1438) );
  OAI21X1 U255 ( .A(n980), .B(n374), .C(n1437), .Y(n1177) );
  OAI21X1 U256 ( .A(n57), .B(n1000), .C(\mem<158> ), .Y(n1437) );
  OAI21X1 U257 ( .A(n978), .B(n374), .C(n1436), .Y(n1176) );
  OAI21X1 U258 ( .A(n54), .B(n1000), .C(\mem<157> ), .Y(n1436) );
  OAI21X1 U259 ( .A(n977), .B(n374), .C(n1435), .Y(n1175) );
  OAI21X1 U260 ( .A(n51), .B(n1000), .C(\mem<156> ), .Y(n1435) );
  OAI21X1 U261 ( .A(n976), .B(n374), .C(n1434), .Y(n1174) );
  OAI21X1 U262 ( .A(n48), .B(n1000), .C(\mem<155> ), .Y(n1434) );
  OAI21X1 U263 ( .A(n974), .B(n374), .C(n1433), .Y(n1173) );
  OAI21X1 U264 ( .A(n45), .B(n1000), .C(\mem<154> ), .Y(n1433) );
  OAI21X1 U265 ( .A(n972), .B(n374), .C(n1432), .Y(n1172) );
  OAI21X1 U266 ( .A(n43), .B(n1000), .C(\mem<153> ), .Y(n1432) );
  OAI21X1 U267 ( .A(n970), .B(n374), .C(n1431), .Y(n1171) );
  OAI21X1 U268 ( .A(n40), .B(n1000), .C(\mem<152> ), .Y(n1431) );
  OAI21X1 U269 ( .A(n968), .B(n374), .C(n1430), .Y(n1170) );
  OAI21X1 U270 ( .A(n37), .B(n999), .C(\mem<151> ), .Y(n1430) );
  OAI21X1 U271 ( .A(n967), .B(n374), .C(n1429), .Y(n1169) );
  OAI21X1 U272 ( .A(n35), .B(n999), .C(\mem<150> ), .Y(n1429) );
  OAI21X1 U273 ( .A(n966), .B(n374), .C(n1428), .Y(n1168) );
  OAI21X1 U274 ( .A(n33), .B(n999), .C(\mem<149> ), .Y(n1428) );
  OAI21X1 U275 ( .A(n965), .B(n374), .C(n1427), .Y(n1167) );
  OAI21X1 U276 ( .A(n31), .B(n999), .C(\mem<148> ), .Y(n1427) );
  OAI21X1 U277 ( .A(n964), .B(n374), .C(n1426), .Y(n1166) );
  OAI21X1 U278 ( .A(n29), .B(n999), .C(\mem<147> ), .Y(n1426) );
  OAI21X1 U279 ( .A(n963), .B(n374), .C(n1425), .Y(n1165) );
  OAI21X1 U280 ( .A(n27), .B(n999), .C(\mem<146> ), .Y(n1425) );
  OAI21X1 U281 ( .A(n962), .B(n374), .C(n1424), .Y(n1164) );
  OAI21X1 U282 ( .A(n25), .B(n999), .C(\mem<145> ), .Y(n1424) );
  OAI21X1 U283 ( .A(n959), .B(n374), .C(n1423), .Y(n1163) );
  OAI21X1 U284 ( .A(n23), .B(n999), .C(\mem<144> ), .Y(n1423) );
  OAI21X1 U287 ( .A(n982), .B(n354), .C(n1422), .Y(n1162) );
  OAI21X1 U288 ( .A(n60), .B(n998), .C(\mem<143> ), .Y(n1422) );
  OAI21X1 U289 ( .A(n980), .B(n354), .C(n1421), .Y(n1161) );
  OAI21X1 U290 ( .A(n57), .B(n998), .C(\mem<142> ), .Y(n1421) );
  OAI21X1 U291 ( .A(n978), .B(n354), .C(n1420), .Y(n1160) );
  OAI21X1 U292 ( .A(n54), .B(n998), .C(\mem<141> ), .Y(n1420) );
  OAI21X1 U293 ( .A(n977), .B(n354), .C(n1419), .Y(n1159) );
  OAI21X1 U294 ( .A(n51), .B(n998), .C(\mem<140> ), .Y(n1419) );
  OAI21X1 U295 ( .A(n976), .B(n354), .C(n1418), .Y(n1158) );
  OAI21X1 U296 ( .A(n48), .B(n998), .C(\mem<139> ), .Y(n1418) );
  OAI21X1 U297 ( .A(n974), .B(n354), .C(n1417), .Y(n1157) );
  OAI21X1 U298 ( .A(n45), .B(n998), .C(\mem<138> ), .Y(n1417) );
  OAI21X1 U299 ( .A(n972), .B(n354), .C(n1416), .Y(n1156) );
  OAI21X1 U300 ( .A(n43), .B(n998), .C(\mem<137> ), .Y(n1416) );
  OAI21X1 U301 ( .A(n970), .B(n354), .C(n1415), .Y(n1155) );
  OAI21X1 U302 ( .A(n40), .B(n998), .C(\mem<136> ), .Y(n1415) );
  OAI21X1 U303 ( .A(n968), .B(n354), .C(n1414), .Y(n1154) );
  OAI21X1 U304 ( .A(n37), .B(n997), .C(\mem<135> ), .Y(n1414) );
  OAI21X1 U305 ( .A(n967), .B(n354), .C(n1413), .Y(n1153) );
  OAI21X1 U306 ( .A(n35), .B(n997), .C(\mem<134> ), .Y(n1413) );
  OAI21X1 U307 ( .A(n966), .B(n354), .C(n1412), .Y(n1152) );
  OAI21X1 U308 ( .A(n33), .B(n997), .C(\mem<133> ), .Y(n1412) );
  OAI21X1 U309 ( .A(n965), .B(n354), .C(n1411), .Y(n1151) );
  OAI21X1 U310 ( .A(n31), .B(n997), .C(\mem<132> ), .Y(n1411) );
  OAI21X1 U311 ( .A(n964), .B(n354), .C(n1410), .Y(n1150) );
  OAI21X1 U312 ( .A(n29), .B(n997), .C(\mem<131> ), .Y(n1410) );
  OAI21X1 U313 ( .A(n963), .B(n354), .C(n1409), .Y(n1149) );
  OAI21X1 U314 ( .A(n27), .B(n997), .C(\mem<130> ), .Y(n1409) );
  OAI21X1 U315 ( .A(n962), .B(n354), .C(n1408), .Y(n1148) );
  OAI21X1 U316 ( .A(n25), .B(n997), .C(\mem<129> ), .Y(n1408) );
  OAI21X1 U317 ( .A(n959), .B(n354), .C(n1407), .Y(n1147) );
  OAI21X1 U318 ( .A(n23), .B(n997), .C(\mem<128> ), .Y(n1407) );
  OAI21X1 U321 ( .A(n981), .B(n333), .C(n1406), .Y(n1146) );
  OAI21X1 U322 ( .A(n60), .B(n995), .C(\mem<127> ), .Y(n1406) );
  OAI21X1 U323 ( .A(n980), .B(n333), .C(n1405), .Y(n1145) );
  OAI21X1 U324 ( .A(n57), .B(n995), .C(\mem<126> ), .Y(n1405) );
  OAI21X1 U325 ( .A(n978), .B(n996), .C(n1404), .Y(n1144) );
  OAI21X1 U326 ( .A(n54), .B(n995), .C(\mem<125> ), .Y(n1404) );
  OAI21X1 U327 ( .A(n977), .B(n996), .C(n1403), .Y(n1143) );
  OAI21X1 U328 ( .A(n51), .B(n995), .C(\mem<124> ), .Y(n1403) );
  OAI21X1 U329 ( .A(n976), .B(n333), .C(n1402), .Y(n1142) );
  OAI21X1 U330 ( .A(n48), .B(n995), .C(\mem<123> ), .Y(n1402) );
  OAI21X1 U331 ( .A(n974), .B(n333), .C(n1401), .Y(n1141) );
  OAI21X1 U332 ( .A(n45), .B(n995), .C(\mem<122> ), .Y(n1401) );
  OAI21X1 U333 ( .A(n972), .B(n333), .C(n1400), .Y(n1140) );
  OAI21X1 U334 ( .A(n43), .B(n995), .C(\mem<121> ), .Y(n1400) );
  OAI21X1 U335 ( .A(n970), .B(n333), .C(n1399), .Y(n1139) );
  OAI21X1 U336 ( .A(n40), .B(n995), .C(\mem<120> ), .Y(n1399) );
  OAI21X1 U337 ( .A(n968), .B(n996), .C(n1398), .Y(n1138) );
  OAI21X1 U338 ( .A(n37), .B(n995), .C(\mem<119> ), .Y(n1398) );
  OAI21X1 U339 ( .A(n967), .B(n996), .C(n1397), .Y(n1137) );
  OAI21X1 U340 ( .A(n35), .B(n995), .C(\mem<118> ), .Y(n1397) );
  OAI21X1 U341 ( .A(n966), .B(n996), .C(n1396), .Y(n1136) );
  OAI21X1 U342 ( .A(n33), .B(n995), .C(\mem<117> ), .Y(n1396) );
  OAI21X1 U343 ( .A(n965), .B(n996), .C(n1395), .Y(n1135) );
  OAI21X1 U344 ( .A(n31), .B(n995), .C(\mem<116> ), .Y(n1395) );
  OAI21X1 U345 ( .A(n964), .B(n996), .C(n1394), .Y(n1134) );
  OAI21X1 U346 ( .A(n29), .B(n995), .C(\mem<115> ), .Y(n1394) );
  OAI21X1 U347 ( .A(n963), .B(n996), .C(n1393), .Y(n1133) );
  OAI21X1 U348 ( .A(n27), .B(n995), .C(\mem<114> ), .Y(n1393) );
  OAI21X1 U349 ( .A(n962), .B(n996), .C(n1392), .Y(n1132) );
  OAI21X1 U350 ( .A(n25), .B(n995), .C(\mem<113> ), .Y(n1392) );
  OAI21X1 U351 ( .A(n959), .B(n996), .C(n1391), .Y(n1131) );
  OAI21X1 U352 ( .A(n23), .B(n995), .C(\mem<112> ), .Y(n1391) );
  OAI21X1 U355 ( .A(n981), .B(n315), .C(n1390), .Y(n1130) );
  OAI21X1 U356 ( .A(n60), .B(n993), .C(\mem<111> ), .Y(n1390) );
  OAI21X1 U357 ( .A(n979), .B(n315), .C(n1389), .Y(n1129) );
  OAI21X1 U358 ( .A(n57), .B(n993), .C(\mem<110> ), .Y(n1389) );
  OAI21X1 U359 ( .A(n978), .B(n994), .C(n1388), .Y(n1128) );
  OAI21X1 U360 ( .A(n54), .B(n993), .C(\mem<109> ), .Y(n1388) );
  OAI21X1 U361 ( .A(n977), .B(n994), .C(n1387), .Y(n1127) );
  OAI21X1 U362 ( .A(n51), .B(n993), .C(\mem<108> ), .Y(n1387) );
  OAI21X1 U363 ( .A(n975), .B(n315), .C(n1386), .Y(n1126) );
  OAI21X1 U364 ( .A(n48), .B(n993), .C(\mem<107> ), .Y(n1386) );
  OAI21X1 U365 ( .A(n973), .B(n315), .C(n1385), .Y(n1125) );
  OAI21X1 U366 ( .A(n45), .B(n993), .C(\mem<106> ), .Y(n1385) );
  OAI21X1 U367 ( .A(n971), .B(n315), .C(n1384), .Y(n1124) );
  OAI21X1 U368 ( .A(n43), .B(n993), .C(\mem<105> ), .Y(n1384) );
  OAI21X1 U369 ( .A(n969), .B(n315), .C(n1383), .Y(n1123) );
  OAI21X1 U370 ( .A(n40), .B(n993), .C(\mem<104> ), .Y(n1383) );
  OAI21X1 U371 ( .A(n968), .B(n994), .C(n1382), .Y(n1122) );
  OAI21X1 U372 ( .A(n37), .B(n993), .C(\mem<103> ), .Y(n1382) );
  OAI21X1 U373 ( .A(n967), .B(n994), .C(n1381), .Y(n1121) );
  OAI21X1 U374 ( .A(n35), .B(n993), .C(\mem<102> ), .Y(n1381) );
  OAI21X1 U375 ( .A(n966), .B(n994), .C(n1380), .Y(n1120) );
  OAI21X1 U376 ( .A(n33), .B(n993), .C(\mem<101> ), .Y(n1380) );
  OAI21X1 U377 ( .A(n965), .B(n994), .C(n1379), .Y(n1119) );
  OAI21X1 U378 ( .A(n31), .B(n993), .C(\mem<100> ), .Y(n1379) );
  OAI21X1 U379 ( .A(n964), .B(n994), .C(n1378), .Y(n1118) );
  OAI21X1 U380 ( .A(n29), .B(n993), .C(\mem<99> ), .Y(n1378) );
  OAI21X1 U381 ( .A(n963), .B(n994), .C(n1377), .Y(n1117) );
  OAI21X1 U382 ( .A(n27), .B(n993), .C(\mem<98> ), .Y(n1377) );
  OAI21X1 U383 ( .A(n962), .B(n994), .C(n1376), .Y(n1116) );
  OAI21X1 U384 ( .A(n25), .B(n993), .C(\mem<97> ), .Y(n1376) );
  OAI21X1 U385 ( .A(n959), .B(n994), .C(n1375), .Y(n1115) );
  OAI21X1 U386 ( .A(n23), .B(n993), .C(\mem<96> ), .Y(n1375) );
  OAI21X1 U389 ( .A(n981), .B(n298), .C(n1374), .Y(n1114) );
  OAI21X1 U390 ( .A(n60), .B(n991), .C(\mem<95> ), .Y(n1374) );
  OAI21X1 U391 ( .A(n979), .B(n298), .C(n1373), .Y(n1113) );
  OAI21X1 U392 ( .A(n57), .B(n991), .C(\mem<94> ), .Y(n1373) );
  OAI21X1 U393 ( .A(n978), .B(n992), .C(n1372), .Y(n1112) );
  OAI21X1 U394 ( .A(n54), .B(n991), .C(\mem<93> ), .Y(n1372) );
  OAI21X1 U395 ( .A(n977), .B(n992), .C(n1371), .Y(n1111) );
  OAI21X1 U396 ( .A(n51), .B(n991), .C(\mem<92> ), .Y(n1371) );
  OAI21X1 U397 ( .A(n975), .B(n298), .C(n1370), .Y(n1110) );
  OAI21X1 U398 ( .A(n48), .B(n991), .C(\mem<91> ), .Y(n1370) );
  OAI21X1 U399 ( .A(n973), .B(n298), .C(n1369), .Y(n1109) );
  OAI21X1 U400 ( .A(n45), .B(n991), .C(\mem<90> ), .Y(n1369) );
  OAI21X1 U401 ( .A(n971), .B(n298), .C(n1368), .Y(n1108) );
  OAI21X1 U402 ( .A(n43), .B(n991), .C(\mem<89> ), .Y(n1368) );
  OAI21X1 U403 ( .A(n969), .B(n298), .C(n1367), .Y(n1107) );
  OAI21X1 U404 ( .A(n40), .B(n991), .C(\mem<88> ), .Y(n1367) );
  OAI21X1 U405 ( .A(n968), .B(n992), .C(n1366), .Y(n1106) );
  OAI21X1 U406 ( .A(n37), .B(n991), .C(\mem<87> ), .Y(n1366) );
  OAI21X1 U407 ( .A(n967), .B(n992), .C(n1365), .Y(n1105) );
  OAI21X1 U408 ( .A(n35), .B(n991), .C(\mem<86> ), .Y(n1365) );
  OAI21X1 U409 ( .A(n966), .B(n992), .C(n1364), .Y(n1104) );
  OAI21X1 U410 ( .A(n33), .B(n991), .C(\mem<85> ), .Y(n1364) );
  OAI21X1 U411 ( .A(n965), .B(n992), .C(n1363), .Y(n1103) );
  OAI21X1 U412 ( .A(n31), .B(n991), .C(\mem<84> ), .Y(n1363) );
  OAI21X1 U413 ( .A(n964), .B(n992), .C(n1362), .Y(n1102) );
  OAI21X1 U414 ( .A(n29), .B(n991), .C(\mem<83> ), .Y(n1362) );
  OAI21X1 U415 ( .A(n963), .B(n992), .C(n1361), .Y(n1101) );
  OAI21X1 U416 ( .A(n27), .B(n991), .C(\mem<82> ), .Y(n1361) );
  OAI21X1 U417 ( .A(n962), .B(n992), .C(n1360), .Y(n1100) );
  OAI21X1 U418 ( .A(n25), .B(n991), .C(\mem<81> ), .Y(n1360) );
  OAI21X1 U419 ( .A(n959), .B(n992), .C(n1359), .Y(n1099) );
  OAI21X1 U420 ( .A(n23), .B(n991), .C(\mem<80> ), .Y(n1359) );
  OAI21X1 U423 ( .A(n981), .B(n280), .C(n1358), .Y(n1098) );
  OAI21X1 U424 ( .A(n60), .B(n989), .C(\mem<79> ), .Y(n1358) );
  OAI21X1 U425 ( .A(n979), .B(n280), .C(n1357), .Y(n1097) );
  OAI21X1 U426 ( .A(n57), .B(n989), .C(\mem<78> ), .Y(n1357) );
  OAI21X1 U427 ( .A(n978), .B(n990), .C(n1356), .Y(n1096) );
  OAI21X1 U428 ( .A(n54), .B(n989), .C(\mem<77> ), .Y(n1356) );
  OAI21X1 U429 ( .A(n977), .B(n990), .C(n1355), .Y(n1095) );
  OAI21X1 U430 ( .A(n51), .B(n989), .C(\mem<76> ), .Y(n1355) );
  OAI21X1 U431 ( .A(n975), .B(n280), .C(n1354), .Y(n1094) );
  OAI21X1 U432 ( .A(n48), .B(n989), .C(\mem<75> ), .Y(n1354) );
  OAI21X1 U433 ( .A(n973), .B(n280), .C(n1353), .Y(n1093) );
  OAI21X1 U434 ( .A(n45), .B(n989), .C(\mem<74> ), .Y(n1353) );
  OAI21X1 U435 ( .A(n971), .B(n280), .C(n1352), .Y(n1092) );
  OAI21X1 U436 ( .A(n43), .B(n989), .C(\mem<73> ), .Y(n1352) );
  OAI21X1 U437 ( .A(n969), .B(n280), .C(n1351), .Y(n1091) );
  OAI21X1 U438 ( .A(n40), .B(n989), .C(\mem<72> ), .Y(n1351) );
  OAI21X1 U439 ( .A(n968), .B(n990), .C(n1350), .Y(n1090) );
  OAI21X1 U440 ( .A(n37), .B(n989), .C(\mem<71> ), .Y(n1350) );
  OAI21X1 U441 ( .A(n967), .B(n990), .C(n1349), .Y(n1089) );
  OAI21X1 U442 ( .A(n35), .B(n989), .C(\mem<70> ), .Y(n1349) );
  OAI21X1 U443 ( .A(n966), .B(n990), .C(n1348), .Y(n1088) );
  OAI21X1 U444 ( .A(n33), .B(n989), .C(\mem<69> ), .Y(n1348) );
  OAI21X1 U445 ( .A(n965), .B(n990), .C(n1347), .Y(n1087) );
  OAI21X1 U446 ( .A(n31), .B(n989), .C(\mem<68> ), .Y(n1347) );
  OAI21X1 U447 ( .A(n964), .B(n990), .C(n1346), .Y(n1086) );
  OAI21X1 U448 ( .A(n29), .B(n989), .C(\mem<67> ), .Y(n1346) );
  OAI21X1 U449 ( .A(n963), .B(n990), .C(n1345), .Y(n1085) );
  OAI21X1 U450 ( .A(n27), .B(n989), .C(\mem<66> ), .Y(n1345) );
  OAI21X1 U451 ( .A(n962), .B(n990), .C(n1344), .Y(n1084) );
  OAI21X1 U452 ( .A(n25), .B(n989), .C(\mem<65> ), .Y(n1344) );
  OAI21X1 U453 ( .A(n959), .B(n990), .C(n1343), .Y(n1083) );
  OAI21X1 U454 ( .A(n23), .B(n989), .C(\mem<64> ), .Y(n1343) );
  OAI21X1 U458 ( .A(n981), .B(n262), .C(n1342), .Y(n1082) );
  OAI21X1 U459 ( .A(n60), .B(n987), .C(\mem<63> ), .Y(n1342) );
  OAI21X1 U460 ( .A(n979), .B(n262), .C(n1341), .Y(n1081) );
  OAI21X1 U461 ( .A(n57), .B(n987), .C(\mem<62> ), .Y(n1341) );
  OAI21X1 U462 ( .A(n978), .B(n988), .C(n1340), .Y(n1080) );
  OAI21X1 U463 ( .A(n54), .B(n987), .C(\mem<61> ), .Y(n1340) );
  OAI21X1 U464 ( .A(n977), .B(n988), .C(n1339), .Y(n1079) );
  OAI21X1 U465 ( .A(n51), .B(n987), .C(\mem<60> ), .Y(n1339) );
  OAI21X1 U466 ( .A(n975), .B(n262), .C(n1338), .Y(n1078) );
  OAI21X1 U467 ( .A(n48), .B(n987), .C(\mem<59> ), .Y(n1338) );
  OAI21X1 U468 ( .A(n973), .B(n262), .C(n1337), .Y(n1077) );
  OAI21X1 U469 ( .A(n45), .B(n987), .C(\mem<58> ), .Y(n1337) );
  OAI21X1 U470 ( .A(n971), .B(n262), .C(n1336), .Y(n1076) );
  OAI21X1 U471 ( .A(n43), .B(n987), .C(\mem<57> ), .Y(n1336) );
  OAI21X1 U472 ( .A(n969), .B(n262), .C(n1335), .Y(n1075) );
  OAI21X1 U473 ( .A(n40), .B(n987), .C(\mem<56> ), .Y(n1335) );
  OAI21X1 U474 ( .A(n968), .B(n988), .C(n1334), .Y(n1074) );
  OAI21X1 U475 ( .A(n37), .B(n987), .C(\mem<55> ), .Y(n1334) );
  OAI21X1 U476 ( .A(n967), .B(n988), .C(n1333), .Y(n1073) );
  OAI21X1 U477 ( .A(n35), .B(n987), .C(\mem<54> ), .Y(n1333) );
  OAI21X1 U478 ( .A(n966), .B(n988), .C(n1332), .Y(n1072) );
  OAI21X1 U479 ( .A(n33), .B(n987), .C(\mem<53> ), .Y(n1332) );
  OAI21X1 U480 ( .A(n965), .B(n988), .C(n1331), .Y(n1071) );
  OAI21X1 U481 ( .A(n31), .B(n987), .C(\mem<52> ), .Y(n1331) );
  OAI21X1 U482 ( .A(n964), .B(n988), .C(n1330), .Y(n1070) );
  OAI21X1 U483 ( .A(n29), .B(n987), .C(\mem<51> ), .Y(n1330) );
  OAI21X1 U484 ( .A(n963), .B(n988), .C(n1329), .Y(n1069) );
  OAI21X1 U485 ( .A(n27), .B(n987), .C(\mem<50> ), .Y(n1329) );
  OAI21X1 U486 ( .A(n962), .B(n988), .C(n1328), .Y(n1068) );
  OAI21X1 U487 ( .A(n25), .B(n987), .C(\mem<49> ), .Y(n1328) );
  OAI21X1 U488 ( .A(n959), .B(n988), .C(n1327), .Y(n1067) );
  OAI21X1 U489 ( .A(n23), .B(n987), .C(\mem<48> ), .Y(n1327) );
  OAI21X1 U492 ( .A(n981), .B(n244), .C(n1326), .Y(n1066) );
  OAI21X1 U493 ( .A(n60), .B(n985), .C(\mem<47> ), .Y(n1326) );
  OAI21X1 U494 ( .A(n979), .B(n244), .C(n1325), .Y(n1065) );
  OAI21X1 U495 ( .A(n57), .B(n985), .C(\mem<46> ), .Y(n1325) );
  OAI21X1 U496 ( .A(n978), .B(n986), .C(n1324), .Y(n1064) );
  OAI21X1 U497 ( .A(n54), .B(n985), .C(\mem<45> ), .Y(n1324) );
  OAI21X1 U498 ( .A(n977), .B(n986), .C(n1323), .Y(n1063) );
  OAI21X1 U499 ( .A(n51), .B(n985), .C(\mem<44> ), .Y(n1323) );
  OAI21X1 U500 ( .A(n975), .B(n244), .C(n1322), .Y(n1062) );
  OAI21X1 U501 ( .A(n48), .B(n985), .C(\mem<43> ), .Y(n1322) );
  OAI21X1 U502 ( .A(n973), .B(n244), .C(n1321), .Y(n1061) );
  OAI21X1 U503 ( .A(n45), .B(n985), .C(\mem<42> ), .Y(n1321) );
  OAI21X1 U504 ( .A(n971), .B(n244), .C(n1320), .Y(n1060) );
  OAI21X1 U505 ( .A(n43), .B(n985), .C(\mem<41> ), .Y(n1320) );
  OAI21X1 U506 ( .A(n969), .B(n244), .C(n1319), .Y(n1059) );
  OAI21X1 U507 ( .A(n40), .B(n985), .C(\mem<40> ), .Y(n1319) );
  OAI21X1 U508 ( .A(n968), .B(n986), .C(n1318), .Y(n1058) );
  OAI21X1 U509 ( .A(n37), .B(n985), .C(\mem<39> ), .Y(n1318) );
  OAI21X1 U510 ( .A(n967), .B(n986), .C(n1317), .Y(n1057) );
  OAI21X1 U511 ( .A(n35), .B(n985), .C(\mem<38> ), .Y(n1317) );
  OAI21X1 U512 ( .A(n966), .B(n986), .C(n1316), .Y(n1056) );
  OAI21X1 U513 ( .A(n33), .B(n985), .C(\mem<37> ), .Y(n1316) );
  OAI21X1 U514 ( .A(n965), .B(n986), .C(n1315), .Y(n1055) );
  OAI21X1 U515 ( .A(n31), .B(n985), .C(\mem<36> ), .Y(n1315) );
  OAI21X1 U516 ( .A(n964), .B(n986), .C(n1314), .Y(n1054) );
  OAI21X1 U517 ( .A(n29), .B(n985), .C(\mem<35> ), .Y(n1314) );
  OAI21X1 U518 ( .A(n963), .B(n986), .C(n1313), .Y(n1053) );
  OAI21X1 U519 ( .A(n27), .B(n985), .C(\mem<34> ), .Y(n1313) );
  OAI21X1 U520 ( .A(n962), .B(n986), .C(n1312), .Y(n1052) );
  OAI21X1 U521 ( .A(n25), .B(n985), .C(\mem<33> ), .Y(n1312) );
  OAI21X1 U522 ( .A(n959), .B(n986), .C(n1311), .Y(n1051) );
  OAI21X1 U523 ( .A(n23), .B(n985), .C(\mem<32> ), .Y(n1311) );
  OAI21X1 U526 ( .A(n981), .B(n241), .C(n1310), .Y(n1050) );
  OAI21X1 U527 ( .A(n60), .B(n983), .C(\mem<31> ), .Y(n1310) );
  OAI21X1 U528 ( .A(n979), .B(n241), .C(n1309), .Y(n1049) );
  OAI21X1 U529 ( .A(n57), .B(n983), .C(\mem<30> ), .Y(n1309) );
  OAI21X1 U530 ( .A(n978), .B(n984), .C(n1308), .Y(n1048) );
  OAI21X1 U531 ( .A(n54), .B(n983), .C(\mem<29> ), .Y(n1308) );
  OAI21X1 U532 ( .A(n977), .B(n984), .C(n1307), .Y(n1047) );
  OAI21X1 U533 ( .A(n51), .B(n983), .C(\mem<28> ), .Y(n1307) );
  OAI21X1 U534 ( .A(n975), .B(n241), .C(n1306), .Y(n1046) );
  OAI21X1 U535 ( .A(n48), .B(n983), .C(\mem<27> ), .Y(n1306) );
  OAI21X1 U536 ( .A(n973), .B(n241), .C(n1305), .Y(n1045) );
  OAI21X1 U537 ( .A(n45), .B(n983), .C(\mem<26> ), .Y(n1305) );
  OAI21X1 U538 ( .A(n971), .B(n241), .C(n1304), .Y(n1044) );
  OAI21X1 U539 ( .A(n43), .B(n983), .C(\mem<25> ), .Y(n1304) );
  OAI21X1 U540 ( .A(n969), .B(n241), .C(n1303), .Y(n1043) );
  OAI21X1 U541 ( .A(n40), .B(n983), .C(\mem<24> ), .Y(n1303) );
  OAI21X1 U542 ( .A(n968), .B(n984), .C(n1302), .Y(n1042) );
  OAI21X1 U543 ( .A(n37), .B(n983), .C(\mem<23> ), .Y(n1302) );
  OAI21X1 U544 ( .A(n967), .B(n984), .C(n1301), .Y(n1041) );
  OAI21X1 U545 ( .A(n35), .B(n983), .C(\mem<22> ), .Y(n1301) );
  OAI21X1 U546 ( .A(n966), .B(n984), .C(n1300), .Y(n1040) );
  OAI21X1 U547 ( .A(n33), .B(n983), .C(\mem<21> ), .Y(n1300) );
  OAI21X1 U548 ( .A(n965), .B(n984), .C(n1299), .Y(n1039) );
  OAI21X1 U549 ( .A(n31), .B(n983), .C(\mem<20> ), .Y(n1299) );
  OAI21X1 U550 ( .A(n964), .B(n984), .C(n1298), .Y(n1038) );
  OAI21X1 U551 ( .A(n29), .B(n983), .C(\mem<19> ), .Y(n1298) );
  OAI21X1 U552 ( .A(n963), .B(n984), .C(n1297), .Y(n1037) );
  OAI21X1 U553 ( .A(n27), .B(n983), .C(\mem<18> ), .Y(n1297) );
  OAI21X1 U554 ( .A(n962), .B(n984), .C(n1296), .Y(n1036) );
  OAI21X1 U555 ( .A(n25), .B(n983), .C(\mem<17> ), .Y(n1296) );
  OAI21X1 U556 ( .A(n959), .B(n984), .C(n1295), .Y(n1035) );
  OAI21X1 U557 ( .A(n23), .B(n983), .C(\mem<16> ), .Y(n1295) );
  OAI21X1 U561 ( .A(n981), .B(n130), .C(n1294), .Y(n1034) );
  OAI21X1 U562 ( .A(n60), .B(n960), .C(\mem<15> ), .Y(n1294) );
  OAI21X1 U565 ( .A(n979), .B(n130), .C(n1291), .Y(n1033) );
  OAI21X1 U566 ( .A(n57), .B(n960), .C(\mem<14> ), .Y(n1291) );
  OAI21X1 U569 ( .A(n978), .B(n961), .C(n1289), .Y(n1032) );
  OAI21X1 U570 ( .A(n54), .B(n960), .C(\mem<13> ), .Y(n1289) );
  OAI21X1 U573 ( .A(n977), .B(n961), .C(n1288), .Y(n1031) );
  OAI21X1 U574 ( .A(n51), .B(n960), .C(\mem<12> ), .Y(n1288) );
  OAI21X1 U577 ( .A(n975), .B(n130), .C(n1287), .Y(n1030) );
  OAI21X1 U578 ( .A(n48), .B(n960), .C(\mem<11> ), .Y(n1287) );
  OAI21X1 U581 ( .A(n973), .B(n130), .C(n1285), .Y(n1029) );
  OAI21X1 U582 ( .A(n45), .B(n960), .C(\mem<10> ), .Y(n1285) );
  OAI21X1 U585 ( .A(n971), .B(n130), .C(n1284), .Y(n1028) );
  OAI21X1 U586 ( .A(n43), .B(n960), .C(\mem<9> ), .Y(n1284) );
  OAI21X1 U589 ( .A(n969), .B(n130), .C(n1283), .Y(n1027) );
  OAI21X1 U590 ( .A(n40), .B(n960), .C(\mem<8> ), .Y(n1283) );
  OAI21X1 U593 ( .A(n968), .B(n961), .C(n1282), .Y(n1026) );
  OAI21X1 U594 ( .A(n37), .B(n960), .C(\mem<7> ), .Y(n1282) );
  OAI21X1 U597 ( .A(n967), .B(n961), .C(n1281), .Y(n1025) );
  OAI21X1 U598 ( .A(n35), .B(n960), .C(\mem<6> ), .Y(n1281) );
  OAI21X1 U601 ( .A(n966), .B(n961), .C(n1280), .Y(n1024) );
  OAI21X1 U602 ( .A(n33), .B(n960), .C(\mem<5> ), .Y(n1280) );
  OAI21X1 U605 ( .A(n965), .B(n961), .C(n1279), .Y(n1023) );
  OAI21X1 U606 ( .A(n31), .B(n960), .C(\mem<4> ), .Y(n1279) );
  OAI21X1 U610 ( .A(n964), .B(n961), .C(n1278), .Y(n1022) );
  OAI21X1 U611 ( .A(n29), .B(n960), .C(\mem<3> ), .Y(n1278) );
  OAI21X1 U614 ( .A(n963), .B(n961), .C(n1277), .Y(n1021) );
  OAI21X1 U615 ( .A(n27), .B(n960), .C(\mem<2> ), .Y(n1277) );
  OAI21X1 U618 ( .A(n962), .B(n961), .C(n1276), .Y(n1020) );
  OAI21X1 U619 ( .A(n25), .B(n960), .C(\mem<1> ), .Y(n1276) );
  OAI21X1 U623 ( .A(n959), .B(n961), .C(n1275), .Y(n1019) );
  OAI21X1 U624 ( .A(n23), .B(n960), .C(\mem<0> ), .Y(n1275) );
  INVX2 U2 ( .A(n652), .Y(n653) );
  BUFX4 U3 ( .A(n315), .Y(n994) );
  BUFX4 U10 ( .A(n298), .Y(n992) );
  BUFX4 U11 ( .A(n280), .Y(n990) );
  BUFX4 U12 ( .A(n262), .Y(n988) );
  BUFX4 U13 ( .A(n244), .Y(n986) );
  BUFX4 U14 ( .A(n241), .Y(n984) );
  BUFX4 U15 ( .A(n130), .Y(n961) );
  BUFX4 U16 ( .A(n333), .Y(n996) );
  AND2X1 U17 ( .A(N25), .B(n1018), .Y(n1455) );
  INVX2 U18 ( .A(N22), .Y(n1017) );
  AND2X1 U19 ( .A(data_in), .B(n112), .Y(n1523) );
  INVX1 U20 ( .A(N19), .Y(n1013) );
  AND2X1 U21 ( .A(N25), .B(N24), .Y(n1522) );
  BUFX2 U22 ( .A(n1523), .Y(n1011) );
  BUFX2 U23 ( .A(n651), .Y(n1009) );
  BUFX2 U24 ( .A(n647), .Y(n1007) );
  BUFX2 U25 ( .A(n639), .Y(n1003) );
  BUFX2 U26 ( .A(n635), .Y(n1001) );
  BUFX2 U27 ( .A(n362), .Y(n999) );
  BUFX2 U28 ( .A(n351), .Y(n997) );
  BUFX2 U29 ( .A(n223), .Y(n981) );
  BUFX2 U30 ( .A(n205), .Y(n979) );
  BUFX2 U31 ( .A(n187), .Y(n975) );
  BUFX2 U32 ( .A(n169), .Y(n973) );
  BUFX2 U33 ( .A(n150), .Y(n971) );
  BUFX2 U34 ( .A(n133), .Y(n969) );
  INVX1 U35 ( .A(n63), .Y(n960) );
  INVX1 U36 ( .A(n78), .Y(n983) );
  INVX1 U37 ( .A(n83), .Y(n989) );
  INVX1 U38 ( .A(n84), .Y(n991) );
  INVX1 U39 ( .A(n89), .Y(n1005) );
  INVX1 U40 ( .A(n93), .Y(n1006) );
  INVX1 U41 ( .A(n80), .Y(n985) );
  INVX1 U42 ( .A(n86), .Y(n993) );
  INVX1 U43 ( .A(n81), .Y(n987) );
  INVX1 U44 ( .A(n87), .Y(n995) );
  BUFX2 U45 ( .A(n187), .Y(n976) );
  BUFX2 U46 ( .A(n205), .Y(n980) );
  BUFX2 U47 ( .A(n223), .Y(n982) );
  BUFX2 U48 ( .A(n133), .Y(n970) );
  INVX1 U81 ( .A(n62), .Y(n959) );
  INVX1 U82 ( .A(n65), .Y(n962) );
  INVX1 U115 ( .A(n66), .Y(n963) );
  INVX1 U116 ( .A(n68), .Y(n964) );
  INVX1 U149 ( .A(n69), .Y(n965) );
  INVX1 U150 ( .A(n71), .Y(n966) );
  INVX1 U183 ( .A(n72), .Y(n967) );
  INVX1 U184 ( .A(n74), .Y(n968) );
  INVX1 U217 ( .A(n1015), .Y(n1014) );
  BUFX2 U218 ( .A(n351), .Y(n998) );
  BUFX2 U251 ( .A(n362), .Y(n1000) );
  BUFX2 U252 ( .A(n635), .Y(n1002) );
  BUFX2 U285 ( .A(n639), .Y(n1004) );
  BUFX2 U286 ( .A(n647), .Y(n1008) );
  BUFX2 U319 ( .A(n651), .Y(n1010) );
  BUFX2 U320 ( .A(n150), .Y(n972) );
  BUFX2 U353 ( .A(n169), .Y(n974) );
  INVX1 U354 ( .A(n75), .Y(n977) );
  INVX1 U387 ( .A(n77), .Y(n978) );
  INVX1 U388 ( .A(N24), .Y(n1018) );
  OR2X2 U421 ( .A(n1014), .B(N21), .Y(n1) );
  INVX1 U422 ( .A(n1), .Y(n2) );
  OR2X2 U455 ( .A(n1015), .B(N21), .Y(n3) );
  INVX1 U456 ( .A(n3), .Y(n4) );
  AND2X2 U457 ( .A(n7), .B(n21), .Y(n5) );
  AND2X2 U490 ( .A(n837), .B(n937), .Y(n6) );
  INVX1 U491 ( .A(n6), .Y(n7) );
  MUX2X1 U524 ( .B(\mem<81> ), .A(\mem<80> ), .S(n671), .Y(n839) );
  INVX1 U525 ( .A(n944), .Y(n8) );
  INVX1 U558 ( .A(n8), .Y(n9) );
  MUX2X1 U559 ( .B(n785), .A(n782), .S(n931), .Y(n796) );
  AND2X1 U560 ( .A(N28), .B(n19), .Y(data_out) );
  INVX1 U563 ( .A(n662), .Y(n10) );
  MUX2X1 U564 ( .B(n900), .A(n899), .S(n934), .Y(n898) );
  MUX2X1 U567 ( .B(\mem<87> ), .A(\mem<86> ), .S(n9), .Y(n837) );
  INVX1 U568 ( .A(n958), .Y(n11) );
  INVX1 U571 ( .A(n11), .Y(n12) );
  INVX1 U572 ( .A(n667), .Y(n13) );
  MUX2X1 U575 ( .B(n918), .A(n917), .S(n934), .Y(n916) );
  INVX2 U576 ( .A(n958), .Y(n667) );
  OR2X1 U579 ( .A(n1016), .B(N23), .Y(n14) );
  INVX1 U580 ( .A(n14), .Y(n15) );
  OR2X1 U583 ( .A(n1017), .B(N23), .Y(n16) );
  INVX1 U584 ( .A(n16), .Y(n17) );
  OR2X2 U587 ( .A(rst), .B(write), .Y(n18) );
  INVX1 U588 ( .A(n18), .Y(n19) );
  AND2X2 U591 ( .A(n836), .B(n933), .Y(n20) );
  INVX1 U592 ( .A(n20), .Y(n21) );
  AND2X1 U595 ( .A(n62), .B(n112), .Y(n22) );
  INVX1 U596 ( .A(n22), .Y(n23) );
  AND2X1 U599 ( .A(n65), .B(n112), .Y(n24) );
  INVX1 U600 ( .A(n24), .Y(n25) );
  AND2X1 U603 ( .A(n66), .B(n112), .Y(n26) );
  INVX1 U604 ( .A(n26), .Y(n27) );
  AND2X1 U607 ( .A(n68), .B(n112), .Y(n28) );
  INVX1 U608 ( .A(n28), .Y(n29) );
  AND2X1 U609 ( .A(n69), .B(n112), .Y(n30) );
  INVX1 U612 ( .A(n30), .Y(n31) );
  AND2X1 U613 ( .A(n71), .B(n112), .Y(n32) );
  INVX1 U616 ( .A(n32), .Y(n33) );
  AND2X1 U617 ( .A(n72), .B(n112), .Y(n34) );
  INVX1 U620 ( .A(n34), .Y(n35) );
  AND2X1 U621 ( .A(n74), .B(n112), .Y(n36) );
  INVX1 U622 ( .A(n36), .Y(n37) );
  AND2X1 U625 ( .A(n131), .B(n112), .Y(n38) );
  INVX1 U626 ( .A(n38), .Y(n40) );
  AND2X1 U627 ( .A(n149), .B(n112), .Y(n41) );
  INVX1 U628 ( .A(n41), .Y(n43) );
  AND2X1 U629 ( .A(n152), .B(n112), .Y(n44) );
  INVX1 U630 ( .A(n44), .Y(n45) );
  AND2X1 U631 ( .A(n171), .B(n112), .Y(n47) );
  INVX1 U632 ( .A(n47), .Y(n48) );
  AND2X1 U633 ( .A(n75), .B(n112), .Y(n50) );
  INVX1 U634 ( .A(n50), .Y(n51) );
  AND2X1 U635 ( .A(n77), .B(n112), .Y(n53) );
  INVX1 U636 ( .A(n53), .Y(n54) );
  AND2X1 U637 ( .A(n189), .B(n112), .Y(n56) );
  INVX1 U638 ( .A(n56), .Y(n57) );
  AND2X1 U639 ( .A(n207), .B(n112), .Y(n59) );
  INVX1 U640 ( .A(n59), .Y(n60) );
  AND2X1 U641 ( .A(n2), .B(n655), .Y(n62) );
  AND2X1 U642 ( .A(n659), .B(n15), .Y(n63) );
  AND2X1 U643 ( .A(n2), .B(n657), .Y(n65) );
  AND2X1 U644 ( .A(n2), .B(n1290), .Y(n66) );
  AND2X1 U645 ( .A(n2), .B(n1292), .Y(n68) );
  AND2X1 U646 ( .A(n4), .B(n655), .Y(n69) );
  AND2X1 U647 ( .A(n4), .B(n657), .Y(n71) );
  AND2X1 U648 ( .A(n4), .B(n1290), .Y(n72) );
  AND2X1 U649 ( .A(n4), .B(n1292), .Y(n74) );
  AND2X1 U650 ( .A(n655), .B(n1293), .Y(n75) );
  AND2X1 U651 ( .A(n657), .B(n1293), .Y(n77) );
  AND2X1 U652 ( .A(n659), .B(n17), .Y(n78) );
  AND2X1 U653 ( .A(n659), .B(n1504), .Y(n80) );
  AND2X1 U654 ( .A(n659), .B(n1521), .Y(n81) );
  AND2X1 U655 ( .A(n661), .B(n15), .Y(n83) );
  AND2X1 U656 ( .A(n661), .B(n17), .Y(n84) );
  AND2X1 U657 ( .A(n661), .B(n1504), .Y(n86) );
  AND2X1 U658 ( .A(n661), .B(n1521), .Y(n87) );
  AND2X1 U659 ( .A(n15), .B(n1522), .Y(n89) );
  AND2X1 U660 ( .A(n17), .B(n1522), .Y(n93) );
  OR2X1 U661 ( .A(n1540), .B(rst), .Y(n95) );
  INVX1 U662 ( .A(n95), .Y(n112) );
  AND2X1 U663 ( .A(n63), .B(n1011), .Y(n114) );
  INVX1 U664 ( .A(n114), .Y(n130) );
  AND2X1 U665 ( .A(n1286), .B(n655), .Y(n131) );
  INVX1 U666 ( .A(n131), .Y(n133) );
  AND2X1 U667 ( .A(n1286), .B(n657), .Y(n149) );
  INVX1 U668 ( .A(n149), .Y(n150) );
  AND2X1 U669 ( .A(n1286), .B(n1290), .Y(n152) );
  INVX1 U670 ( .A(n152), .Y(n169) );
  AND2X1 U671 ( .A(n1286), .B(n1292), .Y(n171) );
  INVX1 U672 ( .A(n171), .Y(n187) );
  AND2X1 U673 ( .A(n1290), .B(n1293), .Y(n189) );
  INVX1 U674 ( .A(n189), .Y(n205) );
  AND2X1 U675 ( .A(n1293), .B(n1292), .Y(n207) );
  INVX1 U676 ( .A(n207), .Y(n223) );
  AND2X1 U677 ( .A(n78), .B(n1011), .Y(n225) );
  INVX1 U678 ( .A(n225), .Y(n241) );
  AND2X1 U679 ( .A(n80), .B(n1011), .Y(n242) );
  INVX1 U680 ( .A(n242), .Y(n244) );
  AND2X1 U681 ( .A(n81), .B(n1011), .Y(n260) );
  INVX1 U682 ( .A(n260), .Y(n262) );
  AND2X1 U683 ( .A(n83), .B(n1011), .Y(n278) );
  INVX1 U684 ( .A(n278), .Y(n280) );
  AND2X1 U685 ( .A(n84), .B(n1011), .Y(n296) );
  INVX1 U686 ( .A(n296), .Y(n298) );
  AND2X1 U687 ( .A(n86), .B(n1011), .Y(n314) );
  INVX1 U688 ( .A(n314), .Y(n315) );
  AND2X1 U689 ( .A(n87), .B(n1011), .Y(n317) );
  INVX1 U690 ( .A(n317), .Y(n333) );
  AND2X1 U691 ( .A(n1455), .B(n15), .Y(n335) );
  INVX1 U692 ( .A(n335), .Y(n351) );
  AND2X1 U693 ( .A(n335), .B(n1523), .Y(n353) );
  INVX1 U694 ( .A(n353), .Y(n354) );
  AND2X1 U695 ( .A(n1455), .B(n17), .Y(n360) );
  INVX1 U696 ( .A(n360), .Y(n362) );
  AND2X1 U697 ( .A(n360), .B(n1523), .Y(n369) );
  INVX1 U698 ( .A(n369), .Y(n374) );
  AND2X1 U699 ( .A(n1455), .B(n1504), .Y(n634) );
  INVX1 U700 ( .A(n634), .Y(n635) );
  AND2X1 U701 ( .A(n634), .B(n1523), .Y(n636) );
  INVX1 U702 ( .A(n636), .Y(n637) );
  AND2X1 U703 ( .A(n1455), .B(n1521), .Y(n638) );
  INVX1 U704 ( .A(n638), .Y(n639) );
  AND2X1 U705 ( .A(n638), .B(n1523), .Y(n640) );
  INVX1 U706 ( .A(n640), .Y(n641) );
  AND2X1 U707 ( .A(n89), .B(n1523), .Y(n642) );
  INVX1 U708 ( .A(n642), .Y(n643) );
  AND2X1 U709 ( .A(n93), .B(n1523), .Y(n644) );
  INVX1 U710 ( .A(n644), .Y(n645) );
  AND2X1 U711 ( .A(n1504), .B(n1522), .Y(n646) );
  INVX1 U712 ( .A(n646), .Y(n647) );
  AND2X1 U713 ( .A(n646), .B(n1523), .Y(n648) );
  INVX1 U714 ( .A(n648), .Y(n649) );
  AND2X1 U715 ( .A(n1522), .B(n1521), .Y(n650) );
  INVX1 U716 ( .A(n650), .Y(n651) );
  AND2X1 U717 ( .A(n1011), .B(n650), .Y(n652) );
  OR2X2 U718 ( .A(n946), .B(n1012), .Y(n654) );
  INVX1 U719 ( .A(n654), .Y(n655) );
  OR2X2 U720 ( .A(n673), .B(n937), .Y(n656) );
  INVX1 U721 ( .A(n656), .Y(n657) );
  OR2X1 U722 ( .A(N24), .B(N25), .Y(n658) );
  INVX1 U723 ( .A(n658), .Y(n659) );
  OR2X1 U724 ( .A(n1018), .B(N25), .Y(n660) );
  INVX1 U725 ( .A(n660), .Y(n661) );
  INVX1 U726 ( .A(n11), .Y(n670) );
  INVX8 U727 ( .A(n944), .Y(n947) );
  INVX1 U728 ( .A(n11), .Y(n663) );
  INVX1 U729 ( .A(n942), .Y(n662) );
  INVX1 U730 ( .A(n942), .Y(n664) );
  INVX1 U731 ( .A(n664), .Y(n665) );
  INVX4 U732 ( .A(n943), .Y(n948) );
  INVX1 U733 ( .A(n664), .Y(n666) );
  MUX2X1 U734 ( .B(\mem<9> ), .A(\mem<8> ), .S(n671), .Y(n911) );
  MUX2X1 U735 ( .B(\mem<175> ), .A(\mem<174> ), .S(n10), .Y(n754) );
  INVX2 U736 ( .A(n958), .Y(n671) );
  MUX2X1 U737 ( .B(\mem<3> ), .A(\mem<2> ), .S(n667), .Y(n918) );
  INVX1 U738 ( .A(n944), .Y(n668) );
  INVX4 U739 ( .A(n944), .Y(n669) );
  MUX2X1 U740 ( .B(n688), .A(n687), .S(n672), .Y(n686) );
  INVX1 U741 ( .A(n928), .Y(n672) );
  MUX2X1 U742 ( .B(\mem<23> ), .A(\mem<22> ), .S(n671), .Y(n900) );
  MUX2X1 U743 ( .B(n796), .A(n795), .S(n927), .Y(n794) );
  MUX2X1 U744 ( .B(n876), .A(n875), .S(n672), .Y(n874) );
  MUX2X1 U745 ( .B(n821), .A(n824), .S(n1015), .Y(n828) );
  INVX1 U746 ( .A(n946), .Y(n673) );
  INVX4 U747 ( .A(n944), .Y(n945) );
  INVX8 U748 ( .A(n943), .Y(n955) );
  MUX2X1 U749 ( .B(\mem<85> ), .A(\mem<84> ), .S(n667), .Y(n836) );
  MUX2X1 U750 ( .B(\mem<17> ), .A(\mem<16> ), .S(n667), .Y(n902) );
  MUX2X1 U751 ( .B(\mem<43> ), .A(\mem<42> ), .S(n666), .Y(n882) );
  INVX1 U752 ( .A(n956), .Y(n957) );
  INVX4 U753 ( .A(n957), .Y(n941) );
  MUX2X1 U754 ( .B(\mem<21> ), .A(\mem<20> ), .S(n665), .Y(n899) );
  INVX2 U755 ( .A(N18), .Y(n956) );
  MUX2X1 U756 ( .B(\mem<89> ), .A(\mem<88> ), .S(n671), .Y(n834) );
  MUX2X1 U757 ( .B(\mem<129> ), .A(\mem<128> ), .S(n671), .Y(n792) );
  MUX2X1 U758 ( .B(n675), .A(n676), .S(n940), .Y(n674) );
  MUX2X1 U759 ( .B(n678), .A(n679), .S(n940), .Y(n677) );
  MUX2X1 U760 ( .B(n681), .A(n682), .S(n940), .Y(n680) );
  MUX2X1 U761 ( .B(n684), .A(n685), .S(n940), .Y(n683) );
  MUX2X1 U762 ( .B(n690), .A(n691), .S(n940), .Y(n689) );
  MUX2X1 U763 ( .B(n693), .A(n694), .S(n940), .Y(n692) );
  MUX2X1 U764 ( .B(n696), .A(n697), .S(n940), .Y(n695) );
  MUX2X1 U765 ( .B(n699), .A(n700), .S(n940), .Y(n698) );
  MUX2X1 U766 ( .B(n702), .A(n703), .S(n929), .Y(n701) );
  MUX2X1 U767 ( .B(n705), .A(n706), .S(n940), .Y(n704) );
  MUX2X1 U768 ( .B(n708), .A(n709), .S(n940), .Y(n707) );
  MUX2X1 U769 ( .B(n711), .A(n712), .S(n940), .Y(n710) );
  MUX2X1 U770 ( .B(n714), .A(n715), .S(n940), .Y(n713) );
  MUX2X1 U771 ( .B(n717), .A(n718), .S(n929), .Y(n716) );
  MUX2X1 U772 ( .B(n720), .A(n721), .S(n939), .Y(n719) );
  MUX2X1 U773 ( .B(n723), .A(n724), .S(n939), .Y(n722) );
  MUX2X1 U774 ( .B(n726), .A(n727), .S(n939), .Y(n725) );
  MUX2X1 U775 ( .B(n729), .A(n730), .S(n939), .Y(n728) );
  MUX2X1 U776 ( .B(n732), .A(n733), .S(n929), .Y(n731) );
  MUX2X1 U777 ( .B(n735), .A(n736), .S(N23), .Y(n734) );
  MUX2X1 U778 ( .B(n738), .A(n739), .S(n939), .Y(n737) );
  MUX2X1 U779 ( .B(n741), .A(n742), .S(n939), .Y(n740) );
  MUX2X1 U780 ( .B(n744), .A(n745), .S(n939), .Y(n743) );
  MUX2X1 U781 ( .B(n747), .A(n748), .S(n939), .Y(n746) );
  MUX2X1 U782 ( .B(n750), .A(n751), .S(n929), .Y(n749) );
  MUX2X1 U783 ( .B(n753), .A(n754), .S(n939), .Y(n752) );
  MUX2X1 U784 ( .B(n756), .A(n757), .S(n939), .Y(n755) );
  MUX2X1 U785 ( .B(n759), .A(n760), .S(n939), .Y(n758) );
  MUX2X1 U786 ( .B(n762), .A(n763), .S(n939), .Y(n761) );
  MUX2X1 U787 ( .B(n765), .A(n766), .S(n929), .Y(n764) );
  MUX2X1 U788 ( .B(n768), .A(n769), .S(n938), .Y(n767) );
  MUX2X1 U789 ( .B(n771), .A(n772), .S(n938), .Y(n770) );
  MUX2X1 U790 ( .B(n774), .A(n775), .S(n938), .Y(n773) );
  MUX2X1 U791 ( .B(n777), .A(n778), .S(n938), .Y(n776) );
  MUX2X1 U792 ( .B(n780), .A(n781), .S(n929), .Y(n779) );
  MUX2X1 U793 ( .B(n783), .A(n784), .S(n938), .Y(n782) );
  MUX2X1 U794 ( .B(n786), .A(n787), .S(n938), .Y(n785) );
  MUX2X1 U795 ( .B(n789), .A(n790), .S(n938), .Y(n788) );
  MUX2X1 U796 ( .B(n792), .A(n793), .S(n938), .Y(n791) );
  MUX2X1 U797 ( .B(n798), .A(n799), .S(N23), .Y(n797) );
  MUX2X1 U798 ( .B(n801), .A(n802), .S(n938), .Y(n800) );
  MUX2X1 U799 ( .B(n804), .A(n805), .S(n938), .Y(n803) );
  MUX2X1 U800 ( .B(n807), .A(n808), .S(n938), .Y(n806) );
  MUX2X1 U801 ( .B(n810), .A(n811), .S(n938), .Y(n809) );
  MUX2X1 U802 ( .B(n813), .A(n814), .S(n929), .Y(n812) );
  MUX2X1 U803 ( .B(n816), .A(n817), .S(n935), .Y(n815) );
  MUX2X1 U804 ( .B(n819), .A(n820), .S(n937), .Y(n818) );
  MUX2X1 U805 ( .B(n822), .A(n823), .S(n936), .Y(n821) );
  MUX2X1 U806 ( .B(n825), .A(n826), .S(n936), .Y(n824) );
  MUX2X1 U807 ( .B(n828), .A(n829), .S(n929), .Y(n827) );
  MUX2X1 U808 ( .B(n831), .A(n832), .S(n935), .Y(n830) );
  MUX2X1 U809 ( .B(n834), .A(n835), .S(n935), .Y(n833) );
  MUX2X1 U810 ( .B(n839), .A(n840), .S(n936), .Y(n838) );
  MUX2X1 U811 ( .B(n842), .A(n843), .S(n929), .Y(n841) );
  MUX2X1 U812 ( .B(n845), .A(n846), .S(n935), .Y(n844) );
  MUX2X1 U813 ( .B(n848), .A(n849), .S(n935), .Y(n847) );
  MUX2X1 U814 ( .B(n851), .A(n852), .S(n935), .Y(n850) );
  MUX2X1 U815 ( .B(n854), .A(n855), .S(n936), .Y(n853) );
  MUX2X1 U816 ( .B(n857), .A(n858), .S(n929), .Y(n856) );
  MUX2X1 U817 ( .B(n860), .A(n861), .S(N23), .Y(n859) );
  MUX2X1 U818 ( .B(n863), .A(n864), .S(n937), .Y(n862) );
  MUX2X1 U819 ( .B(n866), .A(n867), .S(n936), .Y(n865) );
  MUX2X1 U820 ( .B(n869), .A(n870), .S(n937), .Y(n868) );
  MUX2X1 U821 ( .B(n872), .A(n873), .S(n937), .Y(n871) );
  MUX2X1 U822 ( .B(n878), .A(n879), .S(n935), .Y(n877) );
  MUX2X1 U823 ( .B(n881), .A(n882), .S(n937), .Y(n880) );
  MUX2X1 U824 ( .B(n884), .A(n885), .S(n937), .Y(n883) );
  MUX2X1 U825 ( .B(n887), .A(n888), .S(n937), .Y(n886) );
  MUX2X1 U826 ( .B(n890), .A(n891), .S(n928), .Y(n889) );
  MUX2X1 U827 ( .B(n893), .A(n894), .S(n937), .Y(n892) );
  MUX2X1 U828 ( .B(n896), .A(n897), .S(n935), .Y(n895) );
  MUX2X1 U829 ( .B(n902), .A(n903), .S(n935), .Y(n901) );
  MUX2X1 U830 ( .B(n905), .A(n906), .S(n928), .Y(n904) );
  MUX2X1 U831 ( .B(n908), .A(n909), .S(n936), .Y(n907) );
  MUX2X1 U832 ( .B(n911), .A(n912), .S(n936), .Y(n910) );
  MUX2X1 U833 ( .B(n914), .A(n915), .S(n936), .Y(n913) );
  MUX2X1 U834 ( .B(n920), .A(n921), .S(n928), .Y(n919) );
  MUX2X1 U835 ( .B(n923), .A(n924), .S(N23), .Y(n922) );
  MUX2X1 U836 ( .B(n925), .A(n926), .S(N25), .Y(N28) );
  MUX2X1 U837 ( .B(\mem<254> ), .A(\mem<255> ), .S(n670), .Y(n676) );
  MUX2X1 U838 ( .B(\mem<252> ), .A(\mem<253> ), .S(n669), .Y(n675) );
  MUX2X1 U839 ( .B(\mem<250> ), .A(\mem<251> ), .S(n669), .Y(n679) );
  MUX2X1 U840 ( .B(\mem<248> ), .A(\mem<249> ), .S(n945), .Y(n678) );
  MUX2X1 U841 ( .B(n677), .A(n674), .S(n932), .Y(n688) );
  MUX2X1 U842 ( .B(\mem<246> ), .A(\mem<247> ), .S(n946), .Y(n682) );
  MUX2X1 U843 ( .B(\mem<244> ), .A(\mem<245> ), .S(n946), .Y(n681) );
  MUX2X1 U844 ( .B(\mem<242> ), .A(\mem<243> ), .S(n945), .Y(n685) );
  MUX2X1 U845 ( .B(\mem<240> ), .A(\mem<241> ), .S(n945), .Y(n684) );
  MUX2X1 U846 ( .B(n683), .A(n680), .S(n932), .Y(n687) );
  MUX2X1 U847 ( .B(\mem<238> ), .A(\mem<239> ), .S(n946), .Y(n691) );
  MUX2X1 U848 ( .B(\mem<236> ), .A(\mem<237> ), .S(n12), .Y(n690) );
  MUX2X1 U849 ( .B(\mem<234> ), .A(\mem<235> ), .S(n947), .Y(n694) );
  MUX2X1 U850 ( .B(\mem<232> ), .A(\mem<233> ), .S(n946), .Y(n693) );
  MUX2X1 U851 ( .B(n692), .A(n689), .S(n932), .Y(n703) );
  MUX2X1 U852 ( .B(\mem<230> ), .A(\mem<231> ), .S(n946), .Y(n697) );
  MUX2X1 U853 ( .B(\mem<228> ), .A(\mem<229> ), .S(n947), .Y(n696) );
  MUX2X1 U854 ( .B(\mem<226> ), .A(\mem<227> ), .S(n947), .Y(n700) );
  MUX2X1 U855 ( .B(\mem<224> ), .A(\mem<225> ), .S(n669), .Y(n699) );
  MUX2X1 U856 ( .B(n698), .A(n695), .S(n932), .Y(n702) );
  MUX2X1 U857 ( .B(n701), .A(n686), .S(n1016), .Y(n736) );
  MUX2X1 U858 ( .B(\mem<222> ), .A(\mem<223> ), .S(n669), .Y(n706) );
  MUX2X1 U859 ( .B(\mem<220> ), .A(\mem<221> ), .S(n945), .Y(n705) );
  MUX2X1 U860 ( .B(\mem<218> ), .A(\mem<219> ), .S(n946), .Y(n709) );
  MUX2X1 U861 ( .B(\mem<216> ), .A(\mem<217> ), .S(n946), .Y(n708) );
  MUX2X1 U862 ( .B(n707), .A(n704), .S(n932), .Y(n718) );
  MUX2X1 U863 ( .B(\mem<214> ), .A(\mem<215> ), .S(n669), .Y(n712) );
  MUX2X1 U864 ( .B(\mem<212> ), .A(\mem<213> ), .S(n955), .Y(n711) );
  MUX2X1 U865 ( .B(\mem<210> ), .A(\mem<211> ), .S(n669), .Y(n715) );
  MUX2X1 U866 ( .B(\mem<208> ), .A(\mem<209> ), .S(n947), .Y(n714) );
  MUX2X1 U867 ( .B(n713), .A(n710), .S(n932), .Y(n717) );
  MUX2X1 U868 ( .B(\mem<206> ), .A(\mem<207> ), .S(n945), .Y(n721) );
  MUX2X1 U869 ( .B(\mem<204> ), .A(\mem<205> ), .S(n946), .Y(n720) );
  MUX2X1 U870 ( .B(\mem<202> ), .A(\mem<203> ), .S(n947), .Y(n724) );
  MUX2X1 U871 ( .B(\mem<200> ), .A(\mem<201> ), .S(n946), .Y(n723) );
  MUX2X1 U872 ( .B(n722), .A(n719), .S(n932), .Y(n733) );
  MUX2X1 U873 ( .B(\mem<198> ), .A(\mem<199> ), .S(n12), .Y(n727) );
  MUX2X1 U874 ( .B(\mem<196> ), .A(\mem<197> ), .S(n947), .Y(n726) );
  MUX2X1 U875 ( .B(\mem<194> ), .A(\mem<195> ), .S(n945), .Y(n730) );
  MUX2X1 U876 ( .B(\mem<192> ), .A(\mem<193> ), .S(n947), .Y(n729) );
  MUX2X1 U877 ( .B(n728), .A(n725), .S(n932), .Y(n732) );
  MUX2X1 U878 ( .B(n731), .A(n716), .S(n1016), .Y(n735) );
  MUX2X1 U879 ( .B(\mem<190> ), .A(\mem<191> ), .S(n949), .Y(n739) );
  MUX2X1 U880 ( .B(\mem<188> ), .A(\mem<189> ), .S(n950), .Y(n738) );
  MUX2X1 U881 ( .B(\mem<186> ), .A(\mem<187> ), .S(n955), .Y(n742) );
  MUX2X1 U882 ( .B(\mem<184> ), .A(\mem<185> ), .S(n949), .Y(n741) );
  MUX2X1 U883 ( .B(n740), .A(n737), .S(n932), .Y(n751) );
  MUX2X1 U884 ( .B(\mem<182> ), .A(\mem<183> ), .S(n949), .Y(n745) );
  MUX2X1 U885 ( .B(\mem<180> ), .A(\mem<181> ), .S(n949), .Y(n744) );
  MUX2X1 U886 ( .B(\mem<178> ), .A(\mem<179> ), .S(n949), .Y(n748) );
  MUX2X1 U887 ( .B(\mem<176> ), .A(\mem<177> ), .S(n949), .Y(n747) );
  MUX2X1 U888 ( .B(n746), .A(n743), .S(n932), .Y(n750) );
  MUX2X1 U889 ( .B(\mem<172> ), .A(\mem<173> ), .S(n955), .Y(n753) );
  MUX2X1 U890 ( .B(\mem<170> ), .A(\mem<171> ), .S(n952), .Y(n757) );
  MUX2X1 U891 ( .B(\mem<168> ), .A(\mem<169> ), .S(n952), .Y(n756) );
  MUX2X1 U892 ( .B(n755), .A(n752), .S(n932), .Y(n766) );
  MUX2X1 U893 ( .B(\mem<166> ), .A(\mem<167> ), .S(n950), .Y(n760) );
  MUX2X1 U894 ( .B(\mem<164> ), .A(\mem<165> ), .S(n950), .Y(n759) );
  MUX2X1 U895 ( .B(\mem<162> ), .A(\mem<163> ), .S(n952), .Y(n763) );
  MUX2X1 U896 ( .B(\mem<160> ), .A(\mem<161> ), .S(n948), .Y(n762) );
  MUX2X1 U897 ( .B(n761), .A(n758), .S(n932), .Y(n765) );
  MUX2X1 U898 ( .B(n764), .A(n749), .S(n1016), .Y(n799) );
  MUX2X1 U899 ( .B(\mem<158> ), .A(\mem<159> ), .S(n955), .Y(n769) );
  MUX2X1 U900 ( .B(\mem<156> ), .A(\mem<157> ), .S(n948), .Y(n768) );
  MUX2X1 U901 ( .B(\mem<154> ), .A(\mem<155> ), .S(n949), .Y(n772) );
  MUX2X1 U902 ( .B(\mem<152> ), .A(\mem<153> ), .S(n949), .Y(n771) );
  MUX2X1 U903 ( .B(n770), .A(n767), .S(n931), .Y(n781) );
  MUX2X1 U904 ( .B(\mem<150> ), .A(\mem<151> ), .S(n950), .Y(n775) );
  MUX2X1 U905 ( .B(\mem<148> ), .A(\mem<149> ), .S(n950), .Y(n774) );
  MUX2X1 U906 ( .B(\mem<146> ), .A(\mem<147> ), .S(n949), .Y(n778) );
  MUX2X1 U907 ( .B(\mem<144> ), .A(\mem<145> ), .S(n950), .Y(n777) );
  MUX2X1 U908 ( .B(n776), .A(n773), .S(n931), .Y(n780) );
  MUX2X1 U909 ( .B(\mem<142> ), .A(\mem<143> ), .S(n955), .Y(n784) );
  MUX2X1 U910 ( .B(\mem<140> ), .A(\mem<141> ), .S(n950), .Y(n783) );
  MUX2X1 U911 ( .B(\mem<138> ), .A(\mem<139> ), .S(n950), .Y(n787) );
  MUX2X1 U912 ( .B(\mem<136> ), .A(\mem<137> ), .S(n949), .Y(n786) );
  MUX2X1 U913 ( .B(\mem<134> ), .A(\mem<135> ), .S(n948), .Y(n790) );
  MUX2X1 U914 ( .B(\mem<132> ), .A(\mem<133> ), .S(n949), .Y(n789) );
  MUX2X1 U915 ( .B(\mem<130> ), .A(\mem<131> ), .S(n952), .Y(n793) );
  MUX2X1 U916 ( .B(n791), .A(n788), .S(n931), .Y(n795) );
  MUX2X1 U917 ( .B(n794), .A(n779), .S(n1016), .Y(n798) );
  MUX2X1 U918 ( .B(n797), .A(n734), .S(N24), .Y(n926) );
  MUX2X1 U919 ( .B(\mem<126> ), .A(\mem<127> ), .S(n670), .Y(n802) );
  MUX2X1 U920 ( .B(\mem<124> ), .A(\mem<125> ), .S(n950), .Y(n801) );
  MUX2X1 U921 ( .B(\mem<122> ), .A(\mem<123> ), .S(n949), .Y(n805) );
  MUX2X1 U922 ( .B(\mem<120> ), .A(\mem<121> ), .S(n949), .Y(n804) );
  MUX2X1 U923 ( .B(n803), .A(n800), .S(n931), .Y(n814) );
  MUX2X1 U924 ( .B(\mem<118> ), .A(\mem<119> ), .S(n951), .Y(n808) );
  MUX2X1 U925 ( .B(\mem<116> ), .A(\mem<117> ), .S(n955), .Y(n807) );
  MUX2X1 U926 ( .B(\mem<114> ), .A(\mem<115> ), .S(n953), .Y(n811) );
  MUX2X1 U927 ( .B(\mem<112> ), .A(\mem<113> ), .S(n947), .Y(n810) );
  MUX2X1 U928 ( .B(n809), .A(n806), .S(n931), .Y(n813) );
  MUX2X1 U929 ( .B(\mem<110> ), .A(\mem<111> ), .S(n954), .Y(n817) );
  MUX2X1 U930 ( .B(\mem<108> ), .A(\mem<109> ), .S(n953), .Y(n816) );
  MUX2X1 U931 ( .B(\mem<106> ), .A(\mem<107> ), .S(n953), .Y(n820) );
  MUX2X1 U932 ( .B(\mem<104> ), .A(\mem<105> ), .S(n951), .Y(n819) );
  MUX2X1 U933 ( .B(n818), .A(n815), .S(n931), .Y(n829) );
  MUX2X1 U934 ( .B(\mem<102> ), .A(\mem<103> ), .S(n951), .Y(n823) );
  MUX2X1 U935 ( .B(\mem<100> ), .A(\mem<101> ), .S(n953), .Y(n822) );
  MUX2X1 U936 ( .B(\mem<98> ), .A(\mem<99> ), .S(n668), .Y(n826) );
  MUX2X1 U937 ( .B(\mem<96> ), .A(\mem<97> ), .S(n947), .Y(n825) );
  MUX2X1 U938 ( .B(n827), .A(n812), .S(n1016), .Y(n861) );
  MUX2X1 U939 ( .B(\mem<94> ), .A(\mem<95> ), .S(n953), .Y(n832) );
  MUX2X1 U940 ( .B(\mem<92> ), .A(\mem<93> ), .S(n948), .Y(n831) );
  MUX2X1 U941 ( .B(\mem<90> ), .A(\mem<91> ), .S(n663), .Y(n835) );
  MUX2X1 U942 ( .B(n833), .A(n830), .S(n931), .Y(n843) );
  MUX2X1 U943 ( .B(\mem<82> ), .A(\mem<83> ), .S(n951), .Y(n840) );
  MUX2X1 U944 ( .B(n838), .A(n5), .S(n931), .Y(n842) );
  MUX2X1 U945 ( .B(\mem<78> ), .A(\mem<79> ), .S(n668), .Y(n846) );
  MUX2X1 U946 ( .B(\mem<76> ), .A(\mem<77> ), .S(n951), .Y(n845) );
  MUX2X1 U947 ( .B(\mem<74> ), .A(\mem<75> ), .S(n13), .Y(n849) );
  MUX2X1 U948 ( .B(\mem<72> ), .A(\mem<73> ), .S(n953), .Y(n848) );
  MUX2X1 U949 ( .B(n847), .A(n844), .S(n931), .Y(n858) );
  MUX2X1 U950 ( .B(\mem<70> ), .A(\mem<71> ), .S(n953), .Y(n852) );
  MUX2X1 U951 ( .B(\mem<68> ), .A(\mem<69> ), .S(n662), .Y(n851) );
  MUX2X1 U952 ( .B(\mem<66> ), .A(\mem<67> ), .S(n953), .Y(n855) );
  MUX2X1 U953 ( .B(\mem<64> ), .A(\mem<65> ), .S(n952), .Y(n854) );
  MUX2X1 U954 ( .B(n853), .A(n850), .S(n931), .Y(n857) );
  MUX2X1 U955 ( .B(n856), .A(n841), .S(n1016), .Y(n860) );
  MUX2X1 U956 ( .B(\mem<62> ), .A(\mem<63> ), .S(n946), .Y(n864) );
  MUX2X1 U957 ( .B(\mem<60> ), .A(\mem<61> ), .S(n951), .Y(n863) );
  MUX2X1 U958 ( .B(\mem<58> ), .A(\mem<59> ), .S(n951), .Y(n867) );
  MUX2X1 U959 ( .B(\mem<56> ), .A(\mem<57> ), .S(n953), .Y(n866) );
  MUX2X1 U960 ( .B(n865), .A(n862), .S(n930), .Y(n876) );
  MUX2X1 U961 ( .B(\mem<54> ), .A(\mem<55> ), .S(n663), .Y(n870) );
  MUX2X1 U962 ( .B(\mem<52> ), .A(\mem<53> ), .S(n953), .Y(n869) );
  MUX2X1 U963 ( .B(\mem<50> ), .A(\mem<51> ), .S(n951), .Y(n873) );
  MUX2X1 U964 ( .B(\mem<48> ), .A(\mem<49> ), .S(n951), .Y(n872) );
  MUX2X1 U965 ( .B(n871), .A(n868), .S(n930), .Y(n875) );
  MUX2X1 U966 ( .B(\mem<46> ), .A(\mem<47> ), .S(n954), .Y(n879) );
  MUX2X1 U967 ( .B(\mem<44> ), .A(\mem<45> ), .S(n954), .Y(n878) );
  MUX2X1 U968 ( .B(\mem<40> ), .A(\mem<41> ), .S(n955), .Y(n881) );
  MUX2X1 U969 ( .B(n880), .A(n877), .S(n930), .Y(n891) );
  MUX2X1 U970 ( .B(\mem<38> ), .A(\mem<39> ), .S(n954), .Y(n885) );
  MUX2X1 U971 ( .B(\mem<36> ), .A(\mem<37> ), .S(n954), .Y(n884) );
  MUX2X1 U972 ( .B(\mem<34> ), .A(\mem<35> ), .S(n955), .Y(n888) );
  MUX2X1 U973 ( .B(\mem<32> ), .A(\mem<33> ), .S(n950), .Y(n887) );
  MUX2X1 U974 ( .B(n886), .A(n883), .S(n930), .Y(n890) );
  MUX2X1 U975 ( .B(n889), .A(n874), .S(n1016), .Y(n924) );
  MUX2X1 U976 ( .B(\mem<30> ), .A(\mem<31> ), .S(n954), .Y(n894) );
  MUX2X1 U977 ( .B(\mem<28> ), .A(\mem<29> ), .S(n948), .Y(n893) );
  MUX2X1 U978 ( .B(\mem<26> ), .A(\mem<27> ), .S(n954), .Y(n897) );
  MUX2X1 U979 ( .B(\mem<24> ), .A(\mem<25> ), .S(n954), .Y(n896) );
  MUX2X1 U980 ( .B(n895), .A(n892), .S(n930), .Y(n906) );
  MUX2X1 U981 ( .B(\mem<18> ), .A(\mem<19> ), .S(n954), .Y(n903) );
  MUX2X1 U982 ( .B(n901), .A(n898), .S(n930), .Y(n905) );
  MUX2X1 U983 ( .B(\mem<14> ), .A(\mem<15> ), .S(n954), .Y(n909) );
  MUX2X1 U984 ( .B(\mem<12> ), .A(\mem<13> ), .S(n954), .Y(n908) );
  MUX2X1 U985 ( .B(\mem<10> ), .A(\mem<11> ), .S(n955), .Y(n912) );
  MUX2X1 U986 ( .B(n910), .A(n907), .S(n930), .Y(n921) );
  MUX2X1 U987 ( .B(\mem<6> ), .A(\mem<7> ), .S(n954), .Y(n915) );
  MUX2X1 U988 ( .B(\mem<4> ), .A(\mem<5> ), .S(n952), .Y(n914) );
  MUX2X1 U989 ( .B(\mem<0> ), .A(\mem<1> ), .S(n955), .Y(n917) );
  MUX2X1 U990 ( .B(n916), .A(n913), .S(n930), .Y(n920) );
  MUX2X1 U991 ( .B(n919), .A(n904), .S(n1016), .Y(n923) );
  MUX2X1 U992 ( .B(n922), .A(n859), .S(N24), .Y(n925) );
  INVX8 U993 ( .A(N21), .Y(n927) );
  INVX8 U994 ( .A(n927), .Y(n928) );
  INVX8 U995 ( .A(n927), .Y(n929) );
  INVX8 U996 ( .A(n1015), .Y(n930) );
  INVX8 U997 ( .A(n1015), .Y(n931) );
  INVX8 U998 ( .A(n1015), .Y(n932) );
  INVX8 U999 ( .A(n1012), .Y(n933) );
  INVX8 U1000 ( .A(n1012), .Y(n934) );
  INVX8 U1001 ( .A(n934), .Y(n935) );
  INVX8 U1002 ( .A(n934), .Y(n936) );
  INVX8 U1003 ( .A(n934), .Y(n937) );
  INVX8 U1004 ( .A(n933), .Y(n938) );
  INVX8 U1005 ( .A(n933), .Y(n939) );
  INVX8 U1006 ( .A(n933), .Y(n940) );
  INVX8 U1007 ( .A(n958), .Y(n942) );
  INVX8 U1008 ( .A(n958), .Y(n943) );
  INVX8 U1009 ( .A(n958), .Y(n944) );
  INVX8 U1010 ( .A(n944), .Y(n946) );
  INVX8 U1011 ( .A(n941), .Y(n949) );
  INVX8 U1012 ( .A(n942), .Y(n950) );
  INVX8 U1013 ( .A(n942), .Y(n951) );
  INVX8 U1014 ( .A(n943), .Y(n952) );
  INVX8 U1015 ( .A(n942), .Y(n953) );
  INVX8 U1016 ( .A(n941), .Y(n954) );
  INVX8 U1017 ( .A(n956), .Y(n958) );
  INVX1 U1018 ( .A(write), .Y(n1540) );
  INVX8 U1019 ( .A(n1013), .Y(n1012) );
  INVX8 U1020 ( .A(N20), .Y(n1015) );
  INVX8 U1021 ( .A(n1017), .Y(n1016) );
endmodule


module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module cache_cache_id0 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   n164, n166, n167, n165, wr_word0, wr_valid, \w0<15> , \w0<14> ,
         \w0<13> , \w0<12> , \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> ,
         \w0<6> , \w0<5> , \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> ,
         \w1<15> , \w1<14> , \w1<13> , \w1<12> , \w1<11> , \w1<10> , \w1<9> ,
         \w1<8> , \w1<7> , \w1<6> , \w1<5> , \w1<4> , \w1<3> , \w1<2> ,
         \w1<1> , \w1<0> , \w2<15> , \w2<14> , \w2<13> , \w2<12> , \w2<11> ,
         \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , \w2<4> ,
         \w2<3> , \w2<2> , \w2<1> , \w2<0> , \w3<15> , \w3<14> , \w3<13> ,
         \w3<12> , \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> ,
         \w3<5> , \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> , dirtybit,
         validbit, n16, net88848, net88890, net88902, net88913, net91151,
         net91149, net96131, net102527, net102786, net102863, net102994,
         net103295, net107953, net117177, net117176, net121106, net121120,
         net121118, net121138, net121174, net121184, net121183, net121286,
         net121292, net121501, net121509, net121522, net121521, net121520,
         net121593, net121592, net121601, net121612, net121749, net122317,
         net123092, net123091, net125432, net125435, net125434, net125701,
         net125705, net125704, net126451, net126481, net129917, net129933,
         net130107, net130164, net130163, net130177, net126480, net111573,
         net111572, net126936, net126815, net126814, net125431, net121607,
         net126853, net121202, net121201, net121200, net121199, net126450,
         net123450, net123449, net121844, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n17, n19, n20, n21, n22, n24, n25, n26, n28,
         n30, n32, n34, n36, n38, n40, n42, n44, n46, n48, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162;
  assign \tag_out<0>  = net102527;
  assign \tag_out<4>  = net103295;
  assign \tag_out<1>  = net121593;
  assign \data_out<10>  = net126451;

  NOR2X1 U20 ( .A(n91), .B(n16), .Y(wr_valid) );
  memc_Size16_7 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({n139, n137, n135, 
        n133, n131, n129, n127, n111}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word0), .clk(clk), .rst(net91149), .createdump(createdump), 
        .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_6 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({n139, n137, n135, 
        n133, n131, n129, n127, n111}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(net125705), .clk(clk), .rst(net91149), .createdump(createdump), 
        .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_5 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({n139, n137, n135, 
        n133, n131, n129, n127, n111}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(net126481), .clk(clk), .rst(net91149), .createdump(createdump), 
        .file_id({1'b0, 1'b0, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_4 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({n139, n137, n135, 
        n133, n131, n129, n127, n111}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n25), .clk(clk), .rst(net91149), .createdump(createdump), 
        .file_id({1'b0, 1'b0, 1'b0, 1'b1, 1'b1}) );
  memc_Size5_1 mem_tg ( .data_out({n164, n165, \tag_out<2> , n166, n167}), 
        .addr({n139, n137, n135, n133, n131, n129, n127, n125}), .data_in({
        \tag_in<4> , \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), 
        .write(net122317), .clk(clk), .rst(net91149), .createdump(createdump), 
        .file_id({1'b0, 1'b0, 1'b1, 1'b0, 1'b0}) );
  memc_Size1_1 mem_dr ( .data_out(dirtybit), .addr({n139, n137, n135, n133, 
        n131, n129, n127, n111}), .data_in(comp), .write(n106), .clk(clk), 
        .rst(net91149), .createdump(createdump), .file_id({1'b0, 1'b0, 1'b1, 
        1'b0, 1'b1}) );
  memv_1 mem_vl ( .data_out(validbit), .addr({n139, n137, n135, n133, n131, 
        n129, n127, n125}), .data_in(valid_in), .write(net96131), .clk(clk), 
        .rst(net91149), .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  OR2X2 U3 ( .A(n2), .B(n3), .Y(\data_out<13> ) );
  INVX1 U4 ( .A(n159), .Y(n2) );
  INVX1 U5 ( .A(n158), .Y(n3) );
  INVX1 U6 ( .A(net121286), .Y(n4) );
  BUFX2 U7 ( .A(n19), .Y(n5) );
  INVX2 U8 ( .A(net107953), .Y(net130107) );
  INVX1 U9 ( .A(net121118), .Y(n6) );
  AND2X2 U10 ( .A(\offset<2> ), .B(\offset<1> ), .Y(n109) );
  INVX1 U11 ( .A(net121286), .Y(n7) );
  AND2X2 U12 ( .A(n68), .B(n81), .Y(net125434) );
  INVX1 U13 ( .A(n136), .Y(n135) );
  INVX1 U14 ( .A(\index<5> ), .Y(n136) );
  INVX1 U15 ( .A(n138), .Y(n137) );
  INVX1 U16 ( .A(\index<6> ), .Y(n138) );
  INVX1 U17 ( .A(n140), .Y(n139) );
  INVX1 U18 ( .A(\index<7> ), .Y(n140) );
  INVX1 U19 ( .A(\tag_in<4> ), .Y(n15) );
  INVX1 U21 ( .A(\tag_in<3> ), .Y(n92) );
  BUFX2 U22 ( .A(wr_valid), .Y(net122317) );
  BUFX2 U23 ( .A(net122317), .Y(net96131) );
  INVX1 U24 ( .A(net121844), .Y(n16) );
  AND2X2 U25 ( .A(net91151), .B(enable), .Y(net121844) );
  OR2X2 U26 ( .A(n16), .B(net129917), .Y(net88890) );
  INVX8 U27 ( .A(rst), .Y(net91151) );
  AND2X2 U28 ( .A(net121844), .B(validbit), .Y(net125701) );
  AND2X2 U29 ( .A(dirtybit), .B(net121844), .Y(net123091) );
  AND2X2 U30 ( .A(net121844), .B(net121199), .Y(net126853) );
  BUFX2 U31 ( .A(n11), .Y(n10) );
  AOI22X1 U32 ( .A(net121174), .B(\w3<10> ), .C(n9), .D(\w2<10> ), .Y(n11) );
  INVX4 U33 ( .A(net121749), .Y(net121174) );
  INVX1 U34 ( .A(n8), .Y(n9) );
  INVX1 U35 ( .A(net121120), .Y(n8) );
  INVX8 U36 ( .A(net121118), .Y(net121120) );
  AND2X2 U37 ( .A(net123450), .B(n10), .Y(net126450) );
  INVX1 U38 ( .A(net126450), .Y(net126451) );
  INVX1 U39 ( .A(net123449), .Y(net123450) );
  OR2X2 U40 ( .A(n13), .B(n14), .Y(net123449) );
  AND2X2 U41 ( .A(\w0<10> ), .B(net121292), .Y(n13) );
  INVX8 U42 ( .A(net121286), .Y(net121292) );
  AND2X2 U43 ( .A(\w1<10> ), .B(n12), .Y(n14) );
  INVX1 U44 ( .A(net121522), .Y(n12) );
  INVX1 U45 ( .A(net88848), .Y(net121522) );
  NOR3X1 U46 ( .A(net121200), .B(net121201), .C(net121202), .Y(net121199) );
  XOR2X1 U47 ( .A(n166), .B(\tag_in<1> ), .Y(net121200) );
  XNOR2X1 U48 ( .A(n164), .B(n15), .Y(net121201) );
  XOR2X1 U49 ( .A(n167), .B(\tag_in<0> ), .Y(net121202) );
  BUFX2 U50 ( .A(net121199), .Y(net121106) );
  AND2X2 U51 ( .A(net121601), .B(net126853), .Y(hit) );
  AND2X2 U52 ( .A(net125435), .B(net88913), .Y(net121601) );
  INVX1 U53 ( .A(hit), .Y(net126814) );
  AND2X2 U54 ( .A(net126936), .B(net88902), .Y(net121607) );
  INVX1 U55 ( .A(net125431), .Y(net126936) );
  AND2X2 U56 ( .A(net126815), .B(write), .Y(net125431) );
  INVX1 U57 ( .A(net96131), .Y(net88902) );
  INVX1 U58 ( .A(net121607), .Y(net129933) );
  OR2X2 U59 ( .A(net121607), .B(net111573), .Y(net126480) );
  OR2X2 U60 ( .A(net121607), .B(net117177), .Y(net125704) );
  INVX1 U61 ( .A(net126814), .Y(net126815) );
  INVX1 U62 ( .A(net125431), .Y(net125432) );
  INVX8 U63 ( .A(net126480), .Y(net126481) );
  INVX1 U64 ( .A(net111572), .Y(net111573) );
  AND2X1 U65 ( .A(\offset<2> ), .B(n17), .Y(net111572) );
  INVX1 U66 ( .A(\offset<1> ), .Y(n17) );
  INVX4 U67 ( .A(n128), .Y(n127) );
  INVX1 U68 ( .A(\offset<2> ), .Y(net121184) );
  INVX1 U69 ( .A(net107953), .Y(net130177) );
  INVX2 U70 ( .A(net121183), .Y(net121118) );
  INVX1 U71 ( .A(n12), .Y(net130163) );
  INVX1 U72 ( .A(net130163), .Y(net130164) );
  INVX2 U73 ( .A(net121501), .Y(net121286) );
  INVX8 U74 ( .A(n24), .Y(n25) );
  BUFX2 U75 ( .A(net121612), .Y(net129917) );
  OR2X2 U76 ( .A(n64), .B(n86), .Y(\data_out<9> ) );
  AND2X2 U77 ( .A(net125432), .B(net88902), .Y(n19) );
  OR2X2 U78 ( .A(n21), .B(net121749), .Y(n20) );
  INVX1 U79 ( .A(\w3<8> ), .Y(n21) );
  AND2X2 U80 ( .A(n97), .B(n74), .Y(n22) );
  INVX1 U81 ( .A(n22), .Y(\data_out<8> ) );
  OR2X2 U82 ( .A(n19), .B(n110), .Y(n24) );
  AND2X2 U83 ( .A(n69), .B(n53), .Y(n26) );
  INVX1 U84 ( .A(n26), .Y(\data_out<0> ) );
  AND2X2 U85 ( .A(n66), .B(n70), .Y(n28) );
  INVX1 U86 ( .A(n28), .Y(\data_out<1> ) );
  AND2X2 U87 ( .A(n54), .B(n71), .Y(n30) );
  INVX1 U88 ( .A(n30), .Y(\data_out<2> ) );
  AND2X2 U89 ( .A(n55), .B(n72), .Y(n32) );
  INVX1 U90 ( .A(n32), .Y(\data_out<3> ) );
  AND2X2 U91 ( .A(n77), .B(n56), .Y(n34) );
  INVX1 U92 ( .A(n34), .Y(\data_out<4> ) );
  AND2X2 U93 ( .A(n73), .B(n57), .Y(n36) );
  INVX1 U94 ( .A(n36), .Y(\data_out<5> ) );
  AND2X2 U95 ( .A(n79), .B(n58), .Y(n38) );
  INVX1 U96 ( .A(n38), .Y(\data_out<6> ) );
  AND2X2 U97 ( .A(n83), .B(n59), .Y(n40) );
  INVX1 U98 ( .A(n40), .Y(\data_out<7> ) );
  AND2X2 U99 ( .A(n75), .B(n60), .Y(n42) );
  INVX1 U100 ( .A(n42), .Y(\data_out<11> ) );
  AND2X2 U101 ( .A(n85), .B(n61), .Y(n44) );
  INVX1 U102 ( .A(n44), .Y(\data_out<12> ) );
  AND2X2 U103 ( .A(n88), .B(n62), .Y(n46) );
  INVX1 U104 ( .A(n46), .Y(\data_out<14> ) );
  AND2X2 U105 ( .A(n90), .B(n63), .Y(n48) );
  INVX1 U106 ( .A(n48), .Y(\data_out<15> ) );
  AND2X2 U107 ( .A(\offset<1> ), .B(net121184), .Y(n50) );
  INVX1 U108 ( .A(net125704), .Y(net125705) );
  AND2X2 U109 ( .A(\w2<8> ), .B(n6), .Y(n51) );
  INVX1 U110 ( .A(n51), .Y(n52) );
  INVX1 U111 ( .A(net125434), .Y(net125435) );
  BUFX2 U112 ( .A(n142), .Y(n53) );
  BUFX2 U113 ( .A(n145), .Y(n54) );
  BUFX2 U114 ( .A(n147), .Y(n55) );
  BUFX2 U115 ( .A(n149), .Y(n56) );
  BUFX2 U116 ( .A(n151), .Y(n57) );
  BUFX2 U117 ( .A(n152), .Y(n58) );
  BUFX2 U118 ( .A(n153), .Y(n59) );
  BUFX2 U119 ( .A(n156), .Y(n60) );
  BUFX2 U120 ( .A(n157), .Y(n61) );
  BUFX2 U121 ( .A(n160), .Y(n62) );
  BUFX2 U122 ( .A(n161), .Y(n63) );
  OR2X2 U123 ( .A(n98), .B(n99), .Y(n64) );
  OR2X2 U124 ( .A(n100), .B(n101), .Y(n65) );
  INVX1 U125 ( .A(n65), .Y(n66) );
  AND2X2 U126 ( .A(n112), .B(n113), .Y(n67) );
  INVX1 U127 ( .A(n67), .Y(n68) );
  BUFX2 U128 ( .A(n143), .Y(n69) );
  BUFX2 U129 ( .A(n144), .Y(n70) );
  BUFX2 U130 ( .A(n146), .Y(n71) );
  BUFX2 U131 ( .A(n148), .Y(n72) );
  BUFX2 U132 ( .A(n150), .Y(n73) );
  BUFX2 U133 ( .A(n154), .Y(n74) );
  BUFX2 U134 ( .A(n155), .Y(n75) );
  OR2X2 U135 ( .A(n102), .B(n103), .Y(n76) );
  INVX1 U136 ( .A(n76), .Y(n77) );
  OR2X2 U137 ( .A(n104), .B(n105), .Y(n78) );
  INVX1 U138 ( .A(n78), .Y(n79) );
  AND2X2 U139 ( .A(\tag_out<2> ), .B(\tag_in<2> ), .Y(n80) );
  INVX1 U140 ( .A(n80), .Y(n81) );
  OR2X2 U141 ( .A(n115), .B(n116), .Y(n82) );
  INVX1 U142 ( .A(n82), .Y(n83) );
  OR2X2 U143 ( .A(n117), .B(n118), .Y(n84) );
  INVX1 U144 ( .A(n84), .Y(n85) );
  OR2X2 U145 ( .A(n119), .B(n120), .Y(n86) );
  OR2X2 U146 ( .A(n121), .B(n122), .Y(n87) );
  INVX1 U147 ( .A(n87), .Y(n88) );
  OR2X2 U148 ( .A(n124), .B(n123), .Y(n89) );
  INVX1 U149 ( .A(n89), .Y(n90) );
  INVX1 U150 ( .A(n93), .Y(n91) );
  INVX1 U151 ( .A(net123091), .Y(net123092) );
  XOR2X1 U152 ( .A(n165), .B(n92), .Y(net88913) );
  INVX1 U153 ( .A(n93), .Y(n94) );
  AND2X2 U154 ( .A(net121612), .B(n162), .Y(n93) );
  OR2X2 U155 ( .A(net88890), .B(n110), .Y(net121749) );
  INVX1 U156 ( .A(net88890), .Y(net121138) );
  INVX1 U157 ( .A(net121509), .Y(net121612) );
  INVX1 U158 ( .A(net129917), .Y(net121592) );
  BUFX2 U159 ( .A(n166), .Y(net121593) );
  AND2X2 U160 ( .A(net125701), .B(n94), .Y(valid) );
  INVX1 U161 ( .A(net121522), .Y(net121520) );
  INVX1 U162 ( .A(net121522), .Y(net121521) );
  INVX1 U163 ( .A(write), .Y(net121509) );
  NOR3X1 U164 ( .A(\offset<1> ), .B(\offset<2> ), .C(net88890), .Y(net121501)
         );
  BUFX2 U165 ( .A(n165), .Y(\tag_out<3> ) );
  AND2X2 U166 ( .A(n109), .B(net121138), .Y(n96) );
  AND2X2 U167 ( .A(n108), .B(net129933), .Y(wr_word0) );
  AND2X2 U168 ( .A(n52), .B(n20), .Y(n97) );
  AND2X2 U169 ( .A(net121138), .B(n50), .Y(net88848) );
  NOR3X1 U170 ( .A(net121184), .B(\offset<1> ), .C(net88890), .Y(net121183) );
  AND2X2 U171 ( .A(\w0<9> ), .B(n7), .Y(n98) );
  AND2X2 U172 ( .A(net130177), .B(\w1<9> ), .Y(n99) );
  AND2X2 U173 ( .A(\w0<1> ), .B(n7), .Y(n100) );
  AND2X2 U174 ( .A(\w1<1> ), .B(n12), .Y(n101) );
  AND2X2 U175 ( .A(\w2<4> ), .B(n6), .Y(n102) );
  AND2X2 U176 ( .A(\w3<4> ), .B(net121174), .Y(n103) );
  AND2X2 U177 ( .A(n6), .B(\w2<6> ), .Y(n104) );
  AND2X2 U178 ( .A(\w3<6> ), .B(n96), .Y(n105) );
  INVX1 U179 ( .A(n5), .Y(n106) );
  AND2X2 U180 ( .A(net121184), .B(\offset<1> ), .Y(net117176) );
  INVX1 U181 ( .A(net117176), .Y(net117177) );
  OR2X1 U182 ( .A(\offset<1> ), .B(\offset<2> ), .Y(n107) );
  INVX1 U183 ( .A(n107), .Y(n108) );
  INVX1 U184 ( .A(net88848), .Y(net107953) );
  INVX1 U185 ( .A(n109), .Y(n110) );
  BUFX2 U186 ( .A(n164), .Y(net103295) );
  BUFX2 U187 ( .A(n125), .Y(n111) );
  INVX1 U188 ( .A(net121106), .Y(net102994) );
  INVX1 U189 ( .A(net121592), .Y(net102863) );
  INVX1 U190 ( .A(net121601), .Y(net102786) );
  INVX4 U191 ( .A(n126), .Y(n125) );
  INVX1 U192 ( .A(\index<0> ), .Y(n126) );
  INVX1 U193 ( .A(\tag_in<2> ), .Y(n112) );
  INVX1 U194 ( .A(\tag_out<2> ), .Y(n113) );
  INVX1 U195 ( .A(\index<1> ), .Y(n128) );
  BUFX2 U196 ( .A(n167), .Y(net102527) );
  BUFX2 U197 ( .A(\offset<0> ), .Y(err) );
  AND2X2 U198 ( .A(net121120), .B(\w2<7> ), .Y(n115) );
  AND2X2 U199 ( .A(\w3<7> ), .B(net121174), .Y(n116) );
  AND2X2 U200 ( .A(\w2<12> ), .B(n6), .Y(n117) );
  AND2X2 U201 ( .A(\w3<12> ), .B(net121174), .Y(n118) );
  AND2X2 U202 ( .A(\w2<9> ), .B(net121120), .Y(n119) );
  AND2X2 U203 ( .A(\w3<9> ), .B(net121174), .Y(n120) );
  AND2X2 U204 ( .A(\w2<14> ), .B(net121120), .Y(n121) );
  AND2X2 U205 ( .A(\w3<14> ), .B(net121174), .Y(n122) );
  AND2X2 U206 ( .A(\w2<15> ), .B(net121120), .Y(n123) );
  AND2X2 U207 ( .A(\w3<15> ), .B(net121174), .Y(n124) );
  INVX1 U208 ( .A(comp), .Y(n162) );
  INVX8 U209 ( .A(net91151), .Y(net91149) );
  INVX8 U210 ( .A(n130), .Y(n129) );
  INVX8 U211 ( .A(\index<2> ), .Y(n130) );
  INVX8 U212 ( .A(n132), .Y(n131) );
  INVX8 U213 ( .A(\index<3> ), .Y(n132) );
  INVX8 U214 ( .A(n134), .Y(n133) );
  INVX8 U215 ( .A(\index<4> ), .Y(n134) );
  OAI21X1 U216 ( .A(net102994), .B(net102786), .C(comp), .Y(n141) );
  AOI21X1 U217 ( .A(net102863), .B(n141), .C(net123092), .Y(dirty) );
  AOI22X1 U218 ( .A(net121120), .B(\w2<0> ), .C(\w3<0> ), .D(net121174), .Y(
        n143) );
  AOI22X1 U219 ( .A(net121292), .B(\w0<0> ), .C(\w1<0> ), .D(net130107), .Y(
        n142) );
  AOI22X1 U220 ( .A(net121120), .B(\w2<1> ), .C(\w3<1> ), .D(n96), .Y(n144) );
  AOI22X1 U221 ( .A(net121120), .B(\w2<2> ), .C(net121174), .D(\w3<2> ), .Y(
        n146) );
  AOI22X1 U222 ( .A(net121292), .B(\w0<2> ), .C(net121521), .D(\w1<2> ), .Y(
        n145) );
  AOI22X1 U223 ( .A(net121120), .B(\w2<3> ), .C(\w3<3> ), .D(n96), .Y(n148) );
  AOI22X1 U224 ( .A(net121292), .B(\w0<3> ), .C(\w1<3> ), .D(net130107), .Y(
        n147) );
  AOI22X1 U225 ( .A(net121292), .B(\w0<4> ), .C(net121520), .D(\w1<4> ), .Y(
        n149) );
  AOI22X1 U226 ( .A(net121120), .B(\w2<5> ), .C(\w3<5> ), .D(n96), .Y(n151) );
  AOI22X1 U227 ( .A(net121292), .B(\w0<5> ), .C(net130107), .D(\w1<5> ), .Y(
        n150) );
  AOI22X1 U228 ( .A(net121292), .B(\w0<6> ), .C(\w1<6> ), .D(net130107), .Y(
        n152) );
  AOI22X1 U229 ( .A(n7), .B(\w0<7> ), .C(net130164), .D(\w1<7> ), .Y(n153) );
  AOI22X1 U230 ( .A(\w0<8> ), .B(n4), .C(\w1<8> ), .D(net121521), .Y(n154) );
  AOI22X1 U231 ( .A(net121120), .B(\w2<11> ), .C(\w3<11> ), .D(n96), .Y(n156)
         );
  AOI22X1 U232 ( .A(net121292), .B(\w0<11> ), .C(\w1<11> ), .D(net121520), .Y(
        n155) );
  AOI22X1 U233 ( .A(n4), .B(\w0<12> ), .C(net121520), .D(\w1<12> ), .Y(n157)
         );
  AOI22X1 U234 ( .A(net121120), .B(\w2<13> ), .C(net121174), .D(\w3<13> ), .Y(
        n159) );
  AOI22X1 U235 ( .A(\w0<13> ), .B(net121292), .C(net130177), .D(\w1<13> ), .Y(
        n158) );
  AOI22X1 U236 ( .A(net121292), .B(\w0<14> ), .C(net130107), .D(\w1<14> ), .Y(
        n160) );
  AOI22X1 U237 ( .A(\w0<15> ), .B(n4), .C(net121521), .D(\w1<15> ), .Y(n161)
         );
endmodule


module cache_cache_id2 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   n240, n241, n242, wr_word0, wr_word1, wr_word2, wr_word3, \w0<15> ,
         \w0<14> , \w0<13> , \w0<12> , \w0<11> , \w0<10> , \w0<9> , \w0<8> ,
         \w0<7> , \w0<6> , \w0<5> , \w0<4> , \w0<3> , \w0<2> , \w0<1> ,
         \w0<0> , \w1<15> , \w1<14> , \w1<13> , \w1<12> , \w1<11> , \w1<10> ,
         \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , \w1<4> , \w1<3> ,
         \w1<2> , \w1<1> , \w1<0> , \w2<15> , \w2<14> , \w2<13> , \w2<12> ,
         \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> ,
         \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> , \w3<15> , \w3<14> ,
         \w3<13> , \w3<12> , \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> ,
         \w3<6> , \w3<5> , \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> ,
         dirtybit, validbit, n15, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n16, n17, n18, n19, n20, n22, n24, n26, n28, n30, n32,
         n34, n36, n38, n40, n42, n44, n46, n48, n50, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n129, n130, n131, n132, n133, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239;

  NAND2X1 U22 ( .A(n135), .B(n239), .Y(n15) );
  memc_Size16_3 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({n192, n190, n188, 
        n186, n184, n182, n154, n179}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word0), .clk(clk), .rst(n177), .createdump(createdump), 
        .file_id({1'b1, 1'b0, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_2 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({n192, n190, n188, 
        n186, n184, n182, n154, n179}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word1), .clk(clk), .rst(n177), .createdump(createdump), 
        .file_id({1'b1, 1'b0, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_1 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({n192, n190, n188, 
        n186, n184, n182, n157, n179}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word2), .clk(clk), .rst(n177), .createdump(createdump), 
        .file_id({1'b1, 1'b0, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_0 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({n192, n190, n188, 
        n186, n184, n182, n154, n179}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word3), .clk(clk), .rst(n177), .createdump(createdump), 
        .file_id({1'b1, 1'b0, 1'b0, 1'b1, 1'b1}) );
  memc_Size5_0 mem_tg ( .data_out({\tag_out<4> , n240, n241, \tag_out<1> , 
        n242}), .addr({n192, n190, n188, n186, n184, n182, n157, n162}), 
        .data_in({\tag_in<4> , \tag_in<3> , \tag_in<2> , \tag_in<1> , 
        \tag_in<0> }), .write(n160), .clk(clk), .rst(n177), .createdump(
        createdump), .file_id({1'b1, 1'b0, 1'b1, 1'b0, 1'b0}) );
  memc_Size1_0 mem_dr ( .data_out(dirtybit), .addr({n192, n190, n188, n186, 
        n184, n182, n154, n179}), .data_in(comp), .write(n19), .clk(clk), 
        .rst(n177), .createdump(createdump), .file_id({1'b1, 1'b0, 1'b1, 1'b0, 
        1'b1}) );
  memv_0 mem_vl ( .data_out(validbit), .addr({n192, n190, n188, n186, n184, 
        n182, n180, n156}), .data_in(valid_in), .write(n11), .clk(clk), .rst(
        n177), .createdump(createdump), .file_id({1'b1, 1'b0, 1'b0, 1'b0, 1'b0}) );
  AND2X2 U3 ( .A(n205), .B(n55), .Y(n236) );
  INVX2 U4 ( .A(n189), .Y(n188) );
  INVX1 U5 ( .A(\index<5> ), .Y(n189) );
  INVX2 U6 ( .A(n191), .Y(n190) );
  INVX1 U7 ( .A(\index<6> ), .Y(n191) );
  INVX1 U8 ( .A(n193), .Y(n192) );
  INVX1 U9 ( .A(\index<7> ), .Y(n193) );
  INVX1 U10 ( .A(\tag_in<4> ), .Y(n159) );
  BUFX2 U11 ( .A(enable), .Y(n1) );
  BUFX2 U12 ( .A(n168), .Y(n2) );
  AND2X2 U13 ( .A(n124), .B(n3), .Y(n173) );
  AND2X2 U14 ( .A(\offset<2> ), .B(n203), .Y(n3) );
  AND2X2 U15 ( .A(n108), .B(n158), .Y(n58) );
  INVX4 U16 ( .A(n130), .Y(n131) );
  INVX1 U17 ( .A(n241), .Y(n4) );
  AND2X2 U18 ( .A(n124), .B(n5), .Y(n163) );
  OR2X2 U19 ( .A(n204), .B(n203), .Y(n6) );
  INVX8 U20 ( .A(n6), .Y(n5) );
  INVX8 U21 ( .A(n142), .Y(n143) );
  BUFX2 U23 ( .A(n198), .Y(n7) );
  INVX4 U24 ( .A(n201), .Y(n8) );
  INVX1 U25 ( .A(n201), .Y(n235) );
  AND2X2 U26 ( .A(n10), .B(n147), .Y(n20) );
  OR2X2 U27 ( .A(n13), .B(n14), .Y(n9) );
  INVX1 U28 ( .A(n9), .Y(n10) );
  BUFX2 U29 ( .A(n160), .Y(n11) );
  XNOR2X1 U30 ( .A(n159), .B(\tag_out<4> ), .Y(n12) );
  AND2X2 U31 ( .A(n235), .B(\w2<0> ), .Y(n13) );
  AND2X2 U32 ( .A(\w3<0> ), .B(n143), .Y(n14) );
  INVX1 U33 ( .A(n52), .Y(n16) );
  INVX1 U34 ( .A(n242), .Y(n17) );
  AND2X2 U35 ( .A(n195), .B(n141), .Y(n18) );
  INVX1 U36 ( .A(n18), .Y(n19) );
  INVX1 U37 ( .A(n20), .Y(\data_out<0> ) );
  AND2X2 U38 ( .A(n88), .B(n70), .Y(n22) );
  INVX1 U39 ( .A(n22), .Y(\data_out<1> ) );
  AND2X2 U40 ( .A(n89), .B(n71), .Y(n24) );
  INVX1 U41 ( .A(n24), .Y(\data_out<2> ) );
  AND2X2 U42 ( .A(n90), .B(n72), .Y(n26) );
  INVX1 U43 ( .A(n26), .Y(\data_out<3> ) );
  AND2X2 U44 ( .A(n91), .B(n149), .Y(n28) );
  INVX1 U45 ( .A(n28), .Y(\data_out<4> ) );
  AND2X2 U46 ( .A(n92), .B(n73), .Y(n30) );
  INVX1 U47 ( .A(n30), .Y(\data_out<5> ) );
  AND2X2 U48 ( .A(n93), .B(n74), .Y(n32) );
  INVX1 U49 ( .A(n32), .Y(\data_out<6> ) );
  AND2X2 U50 ( .A(n94), .B(n75), .Y(n34) );
  INVX1 U51 ( .A(n34), .Y(\data_out<7> ) );
  AND2X2 U52 ( .A(n95), .B(n76), .Y(n36) );
  INVX1 U53 ( .A(n36), .Y(\data_out<8> ) );
  AND2X2 U54 ( .A(n96), .B(n77), .Y(n38) );
  INVX1 U55 ( .A(n38), .Y(\data_out<9> ) );
  AND2X2 U56 ( .A(n97), .B(n78), .Y(n40) );
  INVX1 U57 ( .A(n40), .Y(\data_out<10> ) );
  AND2X2 U58 ( .A(n98), .B(n79), .Y(n42) );
  INVX1 U59 ( .A(n42), .Y(\data_out<11> ) );
  AND2X2 U60 ( .A(n99), .B(n80), .Y(n44) );
  INVX1 U61 ( .A(n44), .Y(\data_out<12> ) );
  AND2X2 U62 ( .A(n100), .B(n81), .Y(n46) );
  INVX1 U63 ( .A(n46), .Y(\data_out<13> ) );
  AND2X2 U64 ( .A(n101), .B(n82), .Y(n48) );
  INVX1 U65 ( .A(n48), .Y(\data_out<14> ) );
  AND2X2 U66 ( .A(n102), .B(n83), .Y(n50) );
  INVX1 U67 ( .A(n50), .Y(\data_out<15> ) );
  OR2X2 U68 ( .A(n56), .B(n54), .Y(n52) );
  INVX1 U69 ( .A(n52), .Y(n53) );
  OR2X2 U70 ( .A(n57), .B(n12), .Y(n54) );
  AND2X2 U71 ( .A(\offset<1> ), .B(n204), .Y(n55) );
  AND2X2 U72 ( .A(n104), .B(n85), .Y(n56) );
  AND2X2 U73 ( .A(n87), .B(n106), .Y(n57) );
  AND2X2 U74 ( .A(n240), .B(n167), .Y(n59) );
  INVX1 U75 ( .A(n59), .Y(n60) );
  AND2X2 U76 ( .A(n241), .B(n172), .Y(n61) );
  INVX1 U77 ( .A(n61), .Y(n62) );
  OR2X2 U78 ( .A(n200), .B(n7), .Y(n63) );
  INVX1 U79 ( .A(n63), .Y(n64) );
  BUFX2 U80 ( .A(n194), .Y(n65) );
  AND2X2 U81 ( .A(\tag_in<3> ), .B(n168), .Y(n66) );
  INVX1 U82 ( .A(n66), .Y(n67) );
  AND2X2 U83 ( .A(\tag_in<2> ), .B(n4), .Y(n68) );
  INVX1 U84 ( .A(n68), .Y(n69) );
  BUFX2 U85 ( .A(n207), .Y(n70) );
  BUFX2 U86 ( .A(n209), .Y(n71) );
  BUFX2 U87 ( .A(n211), .Y(n72) );
  BUFX2 U88 ( .A(n215), .Y(n73) );
  BUFX2 U89 ( .A(n217), .Y(n74) );
  BUFX2 U90 ( .A(n219), .Y(n75) );
  BUFX2 U91 ( .A(n221), .Y(n76) );
  BUFX2 U92 ( .A(n223), .Y(n77) );
  BUFX2 U93 ( .A(n226), .Y(n78) );
  BUFX2 U94 ( .A(n227), .Y(n79) );
  BUFX2 U95 ( .A(n229), .Y(n80) );
  BUFX2 U96 ( .A(n231), .Y(n81) );
  BUFX2 U97 ( .A(n233), .Y(n82) );
  BUFX2 U98 ( .A(n237), .Y(n83) );
  AND2X2 U99 ( .A(n165), .B(n166), .Y(n84) );
  INVX1 U100 ( .A(n84), .Y(n85) );
  AND2X2 U101 ( .A(n170), .B(n17), .Y(n86) );
  INVX1 U102 ( .A(n86), .Y(n87) );
  BUFX2 U103 ( .A(n208), .Y(n88) );
  BUFX2 U104 ( .A(n210), .Y(n89) );
  BUFX2 U105 ( .A(n212), .Y(n90) );
  BUFX2 U106 ( .A(n214), .Y(n91) );
  BUFX2 U107 ( .A(n216), .Y(n92) );
  BUFX2 U108 ( .A(n218), .Y(n93) );
  BUFX2 U109 ( .A(n220), .Y(n94) );
  BUFX2 U110 ( .A(n222), .Y(n95) );
  BUFX2 U111 ( .A(n224), .Y(n96) );
  BUFX2 U112 ( .A(n225), .Y(n97) );
  BUFX2 U113 ( .A(n228), .Y(n98) );
  BUFX2 U114 ( .A(n230), .Y(n99) );
  BUFX2 U115 ( .A(n232), .Y(n100) );
  BUFX2 U116 ( .A(n234), .Y(n101) );
  BUFX2 U117 ( .A(n238), .Y(n102) );
  AND2X2 U118 ( .A(\tag_in<1> ), .B(\tag_out<1> ), .Y(n103) );
  INVX1 U119 ( .A(n103), .Y(n104) );
  AND2X2 U120 ( .A(\tag_in<0> ), .B(n242), .Y(n105) );
  INVX1 U121 ( .A(n105), .Y(n106) );
  OR2X2 U122 ( .A(n113), .B(n116), .Y(n107) );
  INVX1 U123 ( .A(n107), .Y(n108) );
  AND2X2 U124 ( .A(dirtybit), .B(n158), .Y(n109) );
  INVX1 U125 ( .A(n109), .Y(n110) );
  INVX1 U126 ( .A(n129), .Y(n111) );
  AND2X2 U127 ( .A(n69), .B(n62), .Y(n112) );
  INVX1 U128 ( .A(n112), .Y(n113) );
  INVX1 U129 ( .A(n112), .Y(n114) );
  AND2X2 U130 ( .A(n67), .B(n60), .Y(n115) );
  INVX1 U131 ( .A(n115), .Y(n116) );
  INVX1 U132 ( .A(n115), .Y(n117) );
  AND2X2 U133 ( .A(n153), .B(n174), .Y(n118) );
  INVX1 U134 ( .A(n118), .Y(n119) );
  INVX1 U135 ( .A(n118), .Y(n120) );
  INVX1 U136 ( .A(n118), .Y(n121) );
  AND2X2 U137 ( .A(n195), .B(n65), .Y(n122) );
  INVX1 U138 ( .A(n122), .Y(n123) );
  INVX1 U139 ( .A(n122), .Y(n124) );
  INVX1 U140 ( .A(n122), .Y(n125) );
  AND2X2 U141 ( .A(enable), .B(n126), .Y(n160) );
  AND2X2 U142 ( .A(n198), .B(n178), .Y(n126) );
  INVX1 U143 ( .A(n2), .Y(\tag_out<3> ) );
  INVX1 U144 ( .A(n4), .Y(\tag_out<2> ) );
  OR2X2 U145 ( .A(n114), .B(n117), .Y(n129) );
  OR2X2 U146 ( .A(n139), .B(n202), .Y(n201) );
  INVX8 U147 ( .A(n131), .Y(n132) );
  NOR3X1 U148 ( .A(\offset<1> ), .B(n202), .C(\offset<2> ), .Y(n130) );
  INVX2 U149 ( .A(\offset<1> ), .Y(n203) );
  INVX2 U150 ( .A(\offset<2> ), .Y(n204) );
  INVX2 U151 ( .A(n150), .Y(n133) );
  INVX1 U152 ( .A(n202), .Y(n205) );
  AND2X2 U153 ( .A(n16), .B(n58), .Y(hit) );
  INVX1 U154 ( .A(n153), .Y(n135) );
  INVX2 U155 ( .A(n150), .Y(n136) );
  INVX1 U156 ( .A(\index<0> ), .Y(n137) );
  AND2X2 U157 ( .A(\offset<2> ), .B(n203), .Y(n138) );
  INVX1 U158 ( .A(n138), .Y(n139) );
  AND2X2 U159 ( .A(n169), .B(n135), .Y(n140) );
  INVX1 U160 ( .A(n140), .Y(n141) );
  OR2X2 U161 ( .A(n202), .B(n152), .Y(n142) );
  INVX1 U162 ( .A(n171), .Y(\tag_out<0> ) );
  BUFX2 U163 ( .A(n162), .Y(n145) );
  INVX1 U164 ( .A(n206), .Y(n146) );
  INVX1 U165 ( .A(n146), .Y(n147) );
  INVX1 U166 ( .A(n213), .Y(n148) );
  INVX1 U167 ( .A(n148), .Y(n149) );
  INVX1 U168 ( .A(n236), .Y(n150) );
  AND2X1 U169 ( .A(\offset<1> ), .B(\offset<2> ), .Y(n151) );
  INVX1 U170 ( .A(n151), .Y(n152) );
  INVX1 U171 ( .A(write), .Y(n153) );
  INVX1 U172 ( .A(n196), .Y(n164) );
  BUFX2 U173 ( .A(n180), .Y(n154) );
  INVX1 U174 ( .A(n145), .Y(n155) );
  INVX1 U175 ( .A(n137), .Y(n156) );
  INVX1 U176 ( .A(n181), .Y(n157) );
  INVX1 U177 ( .A(n181), .Y(n180) );
  INVX1 U178 ( .A(n197), .Y(n175) );
  INVX1 U179 ( .A(\index<1> ), .Y(n181) );
  BUFX2 U180 ( .A(n176), .Y(n158) );
  INVX1 U181 ( .A(n11), .Y(n195) );
  BUFX2 U182 ( .A(\offset<0> ), .Y(err) );
  INVX1 U183 ( .A(n137), .Y(n162) );
  INVX1 U184 ( .A(n155), .Y(n179) );
  AND2X2 U185 ( .A(n121), .B(n163), .Y(wr_word3) );
  AND2X2 U186 ( .A(n121), .B(n164), .Y(wr_word1) );
  INVX1 U187 ( .A(\tag_in<1> ), .Y(n165) );
  INVX1 U188 ( .A(\tag_out<1> ), .Y(n166) );
  INVX1 U189 ( .A(\tag_in<3> ), .Y(n167) );
  INVX1 U190 ( .A(n240), .Y(n168) );
  BUFX2 U191 ( .A(hit), .Y(n169) );
  INVX1 U192 ( .A(\tag_in<0> ), .Y(n170) );
  INVX1 U193 ( .A(n242), .Y(n171) );
  INVX1 U194 ( .A(\tag_in<2> ), .Y(n172) );
  AND2X2 U195 ( .A(n120), .B(n173), .Y(wr_word2) );
  INVX1 U196 ( .A(n11), .Y(n174) );
  AND2X2 U197 ( .A(n175), .B(n119), .Y(wr_word0) );
  INVX1 U198 ( .A(comp), .Y(n239) );
  AND2X2 U199 ( .A(n1), .B(n178), .Y(n176) );
  INVX1 U200 ( .A(n158), .Y(n200) );
  INVX1 U201 ( .A(n15), .Y(n198) );
  INVX8 U202 ( .A(n178), .Y(n177) );
  INVX8 U203 ( .A(rst), .Y(n178) );
  INVX8 U204 ( .A(n183), .Y(n182) );
  INVX8 U205 ( .A(\index<2> ), .Y(n183) );
  INVX8 U206 ( .A(n185), .Y(n184) );
  INVX8 U207 ( .A(\index<3> ), .Y(n185) );
  INVX8 U208 ( .A(n187), .Y(n186) );
  INVX8 U209 ( .A(\index<4> ), .Y(n187) );
  NAND3X1 U210 ( .A(n158), .B(n111), .C(n53), .Y(n194) );
  NAND3X1 U211 ( .A(\offset<1> ), .B(n125), .C(n204), .Y(n196) );
  NAND3X1 U212 ( .A(n204), .B(n203), .C(n123), .Y(n197) );
  AND2X2 U213 ( .A(n64), .B(validbit), .Y(valid) );
  OAI21X1 U214 ( .A(n52), .B(n129), .C(comp), .Y(n199) );
  AOI21X1 U215 ( .A(n135), .B(n199), .C(n110), .Y(dirty) );
  OR2X2 U216 ( .A(n200), .B(n135), .Y(n202) );
  AOI22X1 U217 ( .A(\w0<0> ), .B(n132), .C(\w1<0> ), .D(n136), .Y(n206) );
  AOI22X1 U218 ( .A(n8), .B(\w2<1> ), .C(\w3<1> ), .D(n143), .Y(n208) );
  AOI22X1 U219 ( .A(\w0<1> ), .B(n132), .C(\w1<1> ), .D(n136), .Y(n207) );
  AOI22X1 U220 ( .A(n8), .B(\w2<2> ), .C(n143), .D(\w3<2> ), .Y(n210) );
  AOI22X1 U221 ( .A(\w0<2> ), .B(n132), .C(\w1<2> ), .D(n136), .Y(n209) );
  AOI22X1 U222 ( .A(n8), .B(\w2<3> ), .C(n143), .D(\w3<3> ), .Y(n212) );
  AOI22X1 U223 ( .A(\w0<3> ), .B(n132), .C(\w1<3> ), .D(n136), .Y(n211) );
  AOI22X1 U224 ( .A(n8), .B(\w2<4> ), .C(\w3<4> ), .D(n143), .Y(n214) );
  AOI22X1 U225 ( .A(\w0<4> ), .B(n132), .C(\w1<4> ), .D(n136), .Y(n213) );
  AOI22X1 U226 ( .A(n8), .B(\w2<5> ), .C(n143), .D(\w3<5> ), .Y(n216) );
  AOI22X1 U227 ( .A(\w0<5> ), .B(n132), .C(\w1<5> ), .D(n133), .Y(n215) );
  AOI22X1 U228 ( .A(n8), .B(\w2<6> ), .C(\w3<6> ), .D(n143), .Y(n218) );
  AOI22X1 U229 ( .A(\w0<6> ), .B(n132), .C(\w1<6> ), .D(n136), .Y(n217) );
  AOI22X1 U230 ( .A(n8), .B(\w2<7> ), .C(n143), .D(\w3<7> ), .Y(n220) );
  AOI22X1 U231 ( .A(\w0<7> ), .B(n132), .C(\w1<7> ), .D(n133), .Y(n219) );
  AOI22X1 U232 ( .A(n235), .B(\w2<8> ), .C(n143), .D(\w3<8> ), .Y(n222) );
  AOI22X1 U233 ( .A(\w0<8> ), .B(n132), .C(\w1<8> ), .D(n136), .Y(n221) );
  AOI22X1 U234 ( .A(n8), .B(\w2<9> ), .C(\w3<9> ), .D(n143), .Y(n224) );
  AOI22X1 U235 ( .A(\w0<9> ), .B(n132), .C(\w1<9> ), .D(n133), .Y(n223) );
  AOI22X1 U236 ( .A(\w2<10> ), .B(n8), .C(n143), .D(\w3<10> ), .Y(n226) );
  AOI22X1 U237 ( .A(\w0<10> ), .B(n132), .C(\w1<10> ), .D(n133), .Y(n225) );
  AOI22X1 U238 ( .A(n8), .B(\w2<11> ), .C(\w3<11> ), .D(n143), .Y(n228) );
  AOI22X1 U239 ( .A(\w0<11> ), .B(n132), .C(\w1<11> ), .D(n133), .Y(n227) );
  AOI22X1 U240 ( .A(n8), .B(\w2<12> ), .C(\w3<12> ), .D(n143), .Y(n230) );
  AOI22X1 U241 ( .A(\w0<12> ), .B(n132), .C(\w1<12> ), .D(n133), .Y(n229) );
  AOI22X1 U242 ( .A(n235), .B(\w2<13> ), .C(\w3<13> ), .D(n143), .Y(n232) );
  AOI22X1 U243 ( .A(\w0<13> ), .B(n132), .C(\w1<13> ), .D(n136), .Y(n231) );
  AOI22X1 U244 ( .A(n8), .B(\w2<14> ), .C(\w3<14> ), .D(n143), .Y(n234) );
  AOI22X1 U245 ( .A(\w0<14> ), .B(n132), .C(\w1<14> ), .D(n136), .Y(n233) );
  AOI22X1 U246 ( .A(n8), .B(\w2<15> ), .C(n143), .D(\w3<15> ), .Y(n238) );
  AOI22X1 U247 ( .A(n132), .B(\w0<15> ), .C(\w1<15> ), .D(n136), .Y(n237) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module final_memory_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1050, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n373, n374, n375, n376, n377, n378, n380,
         n382, n383, n384, n385, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n403, n404, n405, n406, n407,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n584, n585, n586, n587,
         n588, n589, n590, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n50, n150, n189, n289, n348, n372, n379, n381, n386, n387,
         n401, n402, n409, n421, n422, n434, n435, n447, n448, n460, n461,
         n473, n474, n486, n487, n507, n508, n522, n523, n537, n538, n552,
         n553, n567, n568, n582, n583, n591, n592, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n870), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n869), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n868), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n867), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n866), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n865), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n864), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n863), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n862), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n861), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n860), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n859), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n858), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n857), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n856), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n855), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n854), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n853), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n852), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n851), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n850), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n849), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n848), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n847), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n846), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n845), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n844), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n843), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n842), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n841), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n840), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n839), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n838), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n837), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n836), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n835), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n834), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n833), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n832), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n831), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n830), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n829), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n828), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n827), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n826), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n825), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n824), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n823), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n822), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n821), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n820), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n819), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n818), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n817), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n816), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n815), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n814), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n813), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n812), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n811), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n810), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n809), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n808), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n807), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n806), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n805), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n804), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n803), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n802), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n801), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n800), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n799), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n798), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n797), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n796), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n795), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n794), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n793), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n792), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n791), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n790), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n789), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n788), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n787), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n786), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n785), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n784), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n783), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n782), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n781), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n780), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n779), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n778), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n777), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n776), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n775), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n774), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n773), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n772), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n771), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n770), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n769), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n768), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n767), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n766), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n765), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n764), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n763), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n762), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n761), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n760), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n759), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n758), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n757), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n756), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n755), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n754), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n753), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n752), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n751), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n750), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n749), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n748), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n747), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n746), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n745), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n744), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n743), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n742), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n741), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n740), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n739), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n738), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n737), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n736), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n735), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n734), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n733), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n732), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n731), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n730), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n729), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n728), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n727), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n726), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n725), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n724), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n723), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n722), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n721), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n720), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n719), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n718), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n717), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n716), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n715), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n714), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n713), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n712), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n711), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n710), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n709), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n708), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n707), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n706), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n705), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n704), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n703), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n702), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n701), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n700), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n699), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n698), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n697), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n696), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n695), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n694), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n693), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n692), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n691), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n690), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n689), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n688), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n687), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n686), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n685), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n684), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n683), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n682), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n681), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n680), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n679), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n678), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n677), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n676), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n675), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n674), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n673), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n672), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n671), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n670), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n669), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n668), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n667), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n666), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n665), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n664), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n663), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n662), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n661), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n660), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n659), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n658), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n657), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n656), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n655), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n654), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n653), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n652), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n651), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n650), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n649), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n648), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n647), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n646), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n645), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n644), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n643), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n642), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n641), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n640), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n639), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n638), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n637), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n636), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n635), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n634), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n633), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n632), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n631), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n630), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n629), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n628), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n627), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n626), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n625), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n624), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n623), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n622), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n621), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n620), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n619), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n618), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n617), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n616), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n615), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n614), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n613), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n612), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n611), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n610), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n609), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n608), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n607), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n413), .B(n414), .Y(n412) );
  AND2X2 U10 ( .A(n418), .B(n419), .Y(n417) );
  AND2X2 U11 ( .A(n426), .B(n427), .Y(n425) );
  AND2X2 U12 ( .A(n431), .B(n432), .Y(n430) );
  AND2X2 U13 ( .A(n439), .B(n440), .Y(n438) );
  AND2X2 U14 ( .A(n444), .B(n445), .Y(n443) );
  AND2X2 U15 ( .A(n452), .B(n453), .Y(n451) );
  AND2X2 U16 ( .A(n457), .B(n458), .Y(n456) );
  AND2X2 U17 ( .A(n465), .B(n466), .Y(n464) );
  AND2X2 U18 ( .A(n470), .B(n471), .Y(n469) );
  AND2X2 U19 ( .A(n478), .B(n479), .Y(n477) );
  AND2X2 U20 ( .A(n483), .B(n484), .Y(n482) );
  AND2X2 U21 ( .A(n491), .B(n492), .Y(n490) );
  AND2X2 U22 ( .A(n496), .B(n497), .Y(n495) );
  AND2X2 U30 ( .A(n588), .B(n1030), .Y(n248) );
  AND2X2 U31 ( .A(n589), .B(n1030), .Y(n91) );
  AND2X2 U32 ( .A(n588), .B(\addr_1c<0> ), .Y(n228) );
  AND2X2 U33 ( .A(n589), .B(\addr_1c<0> ), .Y(n71) );
  AND2X2 U34 ( .A(n596), .B(n597), .Y(n595) );
  AND2X2 U45 ( .A(n603), .B(n604), .Y(n602) );
  NOR3X1 U94 ( .A(n1019), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1018), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1042), .C(n40), .Y(n607) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n40) );
  OAI21X1 U98 ( .A(n1011), .B(n1043), .C(n41), .Y(n608) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n41) );
  OAI21X1 U100 ( .A(n1011), .B(n1044), .C(n42), .Y(n609) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n42) );
  OAI21X1 U102 ( .A(n1011), .B(n1045), .C(n43), .Y(n610) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n43) );
  OAI21X1 U104 ( .A(n1011), .B(n1046), .C(n44), .Y(n611) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n44) );
  OAI21X1 U106 ( .A(n1011), .B(n1047), .C(n45), .Y(n612) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n45) );
  OAI21X1 U108 ( .A(n1011), .B(n1048), .C(n46), .Y(n613) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n46) );
  OAI21X1 U110 ( .A(n1011), .B(n1049), .C(n47), .Y(n614) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n47) );
  NAND3X1 U112 ( .A(n48), .B(n49), .C(n964), .Y(n39) );
  OAI21X1 U113 ( .A(n6), .B(n1034), .C(n51), .Y(n615) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n51) );
  OAI21X1 U115 ( .A(n6), .B(n1035), .C(n52), .Y(n616) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n52) );
  OAI21X1 U117 ( .A(n6), .B(n1036), .C(n53), .Y(n617) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n53) );
  OAI21X1 U119 ( .A(n6), .B(n1037), .C(n54), .Y(n618) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n54) );
  OAI21X1 U121 ( .A(n6), .B(n1038), .C(n55), .Y(n619) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n55) );
  OAI21X1 U123 ( .A(n6), .B(n1039), .C(n56), .Y(n620) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n56) );
  OAI21X1 U125 ( .A(n6), .B(n1040), .C(n57), .Y(n621) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n57) );
  OAI21X1 U127 ( .A(n6), .B(n1041), .C(n58), .Y(n622) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n58) );
  OAI21X1 U130 ( .A(n1042), .B(n1010), .C(n62), .Y(n623) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n62) );
  OAI21X1 U132 ( .A(n1043), .B(n1009), .C(n63), .Y(n624) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n63) );
  OAI21X1 U134 ( .A(n1044), .B(n1009), .C(n64), .Y(n625) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n64) );
  OAI21X1 U136 ( .A(n1045), .B(n1009), .C(n65), .Y(n626) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n65) );
  OAI21X1 U138 ( .A(n1046), .B(n1009), .C(n66), .Y(n627) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n66) );
  OAI21X1 U140 ( .A(n1047), .B(n1009), .C(n67), .Y(n628) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n67) );
  OAI21X1 U142 ( .A(n1048), .B(n1009), .C(n68), .Y(n629) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n68) );
  OAI21X1 U144 ( .A(n1049), .B(n1009), .C(n69), .Y(n630) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n69) );
  NAND3X1 U146 ( .A(n70), .B(n48), .C(n71), .Y(n61) );
  OAI21X1 U147 ( .A(n1034), .B(n1008), .C(n73), .Y(n631) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n73) );
  OAI21X1 U149 ( .A(n1035), .B(n1008), .C(n74), .Y(n632) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n74) );
  OAI21X1 U151 ( .A(n1036), .B(n1008), .C(n75), .Y(n633) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n75) );
  OAI21X1 U153 ( .A(n1037), .B(n1008), .C(n76), .Y(n634) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n76) );
  OAI21X1 U155 ( .A(n1038), .B(n1008), .C(n77), .Y(n635) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n77) );
  OAI21X1 U157 ( .A(n1039), .B(n1008), .C(n78), .Y(n636) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n78) );
  OAI21X1 U159 ( .A(n1040), .B(n1008), .C(n79), .Y(n637) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n79) );
  OAI21X1 U161 ( .A(n1041), .B(n1008), .C(n80), .Y(n638) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n80) );
  NAND3X1 U163 ( .A(n973), .B(n48), .C(n81), .Y(n72) );
  OAI21X1 U164 ( .A(n1042), .B(n1007), .C(n83), .Y(n639) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n83) );
  OAI21X1 U166 ( .A(n1043), .B(n1006), .C(n84), .Y(n640) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n84) );
  OAI21X1 U168 ( .A(n1044), .B(n1006), .C(n85), .Y(n641) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n85) );
  OAI21X1 U170 ( .A(n1045), .B(n1006), .C(n86), .Y(n642) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n86) );
  OAI21X1 U172 ( .A(n1046), .B(n1006), .C(n87), .Y(n643) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n87) );
  OAI21X1 U174 ( .A(n1047), .B(n1006), .C(n88), .Y(n644) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n88) );
  OAI21X1 U176 ( .A(n1048), .B(n1006), .C(n89), .Y(n645) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n89) );
  OAI21X1 U178 ( .A(n1049), .B(n1006), .C(n90), .Y(n646) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n90) );
  NAND3X1 U180 ( .A(n70), .B(n48), .C(n91), .Y(n82) );
  OAI21X1 U181 ( .A(n1034), .B(n1005), .C(n93), .Y(n647) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n93) );
  OAI21X1 U183 ( .A(n1035), .B(n1005), .C(n94), .Y(n648) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n94) );
  OAI21X1 U185 ( .A(n1036), .B(n1005), .C(n95), .Y(n649) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n95) );
  OAI21X1 U187 ( .A(n1037), .B(n1005), .C(n96), .Y(n650) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n96) );
  OAI21X1 U189 ( .A(n1038), .B(n1005), .C(n97), .Y(n651) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n97) );
  OAI21X1 U191 ( .A(n1039), .B(n1005), .C(n98), .Y(n652) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n98) );
  OAI21X1 U193 ( .A(n1040), .B(n1005), .C(n99), .Y(n653) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n99) );
  OAI21X1 U195 ( .A(n1041), .B(n1005), .C(n100), .Y(n654) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n100) );
  NAND3X1 U197 ( .A(n973), .B(n48), .C(n101), .Y(n92) );
  OAI21X1 U198 ( .A(n1042), .B(n1004), .C(n103), .Y(n655) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n103) );
  OAI21X1 U200 ( .A(n1043), .B(n1003), .C(n104), .Y(n656) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n104) );
  OAI21X1 U202 ( .A(n1044), .B(n1003), .C(n105), .Y(n657) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n105) );
  OAI21X1 U204 ( .A(n1045), .B(n1003), .C(n106), .Y(n658) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n106) );
  OAI21X1 U206 ( .A(n1046), .B(n1003), .C(n107), .Y(n659) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n107) );
  OAI21X1 U208 ( .A(n1047), .B(n1003), .C(n108), .Y(n660) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n108) );
  OAI21X1 U210 ( .A(n1048), .B(n1003), .C(n109), .Y(n661) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n109) );
  OAI21X1 U212 ( .A(n1049), .B(n1003), .C(n110), .Y(n662) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n110) );
  NAND3X1 U214 ( .A(n71), .B(n1013), .C(n111), .Y(n102) );
  OAI21X1 U215 ( .A(n1034), .B(n1002), .C(n113), .Y(n663) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n113) );
  OAI21X1 U217 ( .A(n1035), .B(n1002), .C(n114), .Y(n664) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n114) );
  OAI21X1 U219 ( .A(n1036), .B(n1002), .C(n115), .Y(n665) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n115) );
  OAI21X1 U221 ( .A(n1037), .B(n1002), .C(n116), .Y(n666) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n116) );
  OAI21X1 U223 ( .A(n1038), .B(n1002), .C(n117), .Y(n667) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n117) );
  OAI21X1 U225 ( .A(n1039), .B(n1002), .C(n118), .Y(n668) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n118) );
  OAI21X1 U227 ( .A(n1040), .B(n1002), .C(n119), .Y(n669) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n119) );
  OAI21X1 U229 ( .A(n1041), .B(n1002), .C(n120), .Y(n670) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n120) );
  NAND3X1 U231 ( .A(n973), .B(n1013), .C(n121), .Y(n112) );
  OAI21X1 U232 ( .A(n1042), .B(n1001), .C(n123), .Y(n671) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n123) );
  OAI21X1 U234 ( .A(n1043), .B(n1000), .C(n124), .Y(n672) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n124) );
  OAI21X1 U236 ( .A(n1044), .B(n1000), .C(n125), .Y(n673) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n125) );
  OAI21X1 U238 ( .A(n1045), .B(n1000), .C(n126), .Y(n674) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n126) );
  OAI21X1 U240 ( .A(n1046), .B(n1000), .C(n127), .Y(n675) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n127) );
  OAI21X1 U242 ( .A(n1047), .B(n1000), .C(n128), .Y(n676) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n128) );
  OAI21X1 U244 ( .A(n1048), .B(n1000), .C(n129), .Y(n677) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n129) );
  OAI21X1 U246 ( .A(n1049), .B(n1000), .C(n130), .Y(n678) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n130) );
  NAND3X1 U248 ( .A(n91), .B(n1013), .C(n111), .Y(n122) );
  OAI21X1 U249 ( .A(n1034), .B(n999), .C(n132), .Y(n679) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n132) );
  OAI21X1 U251 ( .A(n1035), .B(n999), .C(n133), .Y(n680) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n133) );
  OAI21X1 U253 ( .A(n1036), .B(n999), .C(n134), .Y(n681) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n134) );
  OAI21X1 U255 ( .A(n1037), .B(n999), .C(n135), .Y(n682) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n135) );
  OAI21X1 U257 ( .A(n1038), .B(n999), .C(n136), .Y(n683) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n136) );
  OAI21X1 U259 ( .A(n1039), .B(n999), .C(n137), .Y(n684) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n137) );
  OAI21X1 U261 ( .A(n1040), .B(n999), .C(n138), .Y(n685) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n138) );
  OAI21X1 U263 ( .A(n1041), .B(n999), .C(n139), .Y(n686) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n139) );
  NAND3X1 U265 ( .A(n973), .B(n1013), .C(n140), .Y(n131) );
  OAI21X1 U266 ( .A(n1042), .B(n998), .C(n142), .Y(n687) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n142) );
  OAI21X1 U268 ( .A(n1043), .B(n998), .C(n143), .Y(n688) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n143) );
  OAI21X1 U270 ( .A(n1044), .B(n998), .C(n144), .Y(n689) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n144) );
  OAI21X1 U272 ( .A(n1045), .B(n998), .C(n145), .Y(n690) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n145) );
  OAI21X1 U274 ( .A(n1046), .B(n998), .C(n146), .Y(n691) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n146) );
  OAI21X1 U276 ( .A(n1047), .B(n998), .C(n147), .Y(n692) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n147) );
  OAI21X1 U278 ( .A(n1048), .B(n998), .C(n148), .Y(n693) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n148) );
  OAI21X1 U280 ( .A(n1049), .B(n998), .C(n149), .Y(n694) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n149) );
  NAND3X1 U282 ( .A(n71), .B(n1013), .C(n969), .Y(n141) );
  OAI21X1 U283 ( .A(n1034), .B(n997), .C(n152), .Y(n695) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n152) );
  OAI21X1 U285 ( .A(n1035), .B(n997), .C(n153), .Y(n696) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n153) );
  OAI21X1 U287 ( .A(n1036), .B(n997), .C(n154), .Y(n697) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n154) );
  OAI21X1 U289 ( .A(n1037), .B(n997), .C(n155), .Y(n698) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n155) );
  OAI21X1 U291 ( .A(n1038), .B(n997), .C(n156), .Y(n699) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n156) );
  OAI21X1 U293 ( .A(n1039), .B(n997), .C(n157), .Y(n700) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n157) );
  OAI21X1 U295 ( .A(n1040), .B(n997), .C(n158), .Y(n701) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n158) );
  OAI21X1 U297 ( .A(n1041), .B(n997), .C(n159), .Y(n702) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n159) );
  NAND3X1 U299 ( .A(n973), .B(n1013), .C(n160), .Y(n151) );
  OAI21X1 U300 ( .A(n1042), .B(n996), .C(n162), .Y(n703) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n162) );
  OAI21X1 U302 ( .A(n1043), .B(n996), .C(n163), .Y(n704) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n163) );
  OAI21X1 U304 ( .A(n1044), .B(n996), .C(n164), .Y(n705) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n164) );
  OAI21X1 U306 ( .A(n1045), .B(n996), .C(n165), .Y(n706) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n165) );
  OAI21X1 U308 ( .A(n1046), .B(n996), .C(n166), .Y(n707) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n166) );
  OAI21X1 U310 ( .A(n1047), .B(n996), .C(n167), .Y(n708) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n167) );
  OAI21X1 U312 ( .A(n1048), .B(n996), .C(n168), .Y(n709) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n168) );
  OAI21X1 U314 ( .A(n1049), .B(n996), .C(n169), .Y(n710) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n169) );
  NAND3X1 U316 ( .A(n91), .B(n1013), .C(n969), .Y(n161) );
  OAI21X1 U317 ( .A(n1034), .B(n995), .C(n171), .Y(n711) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n171) );
  OAI21X1 U319 ( .A(n1035), .B(n995), .C(n172), .Y(n712) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n172) );
  OAI21X1 U321 ( .A(n1036), .B(n995), .C(n173), .Y(n713) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n173) );
  OAI21X1 U323 ( .A(n1037), .B(n995), .C(n174), .Y(n714) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n174) );
  OAI21X1 U325 ( .A(n1038), .B(n995), .C(n175), .Y(n715) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n175) );
  OAI21X1 U327 ( .A(n1039), .B(n995), .C(n176), .Y(n716) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n176) );
  OAI21X1 U329 ( .A(n1040), .B(n995), .C(n177), .Y(n717) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n177) );
  OAI21X1 U331 ( .A(n1041), .B(n995), .C(n178), .Y(n718) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n178) );
  NAND3X1 U333 ( .A(n973), .B(n1013), .C(n179), .Y(n170) );
  OAI21X1 U334 ( .A(n1042), .B(n994), .C(n181), .Y(n719) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n181) );
  OAI21X1 U336 ( .A(n1043), .B(n994), .C(n182), .Y(n720) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n182) );
  OAI21X1 U338 ( .A(n1044), .B(n994), .C(n183), .Y(n721) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n183) );
  OAI21X1 U340 ( .A(n1045), .B(n994), .C(n184), .Y(n722) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n184) );
  OAI21X1 U342 ( .A(n1046), .B(n994), .C(n185), .Y(n723) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n185) );
  OAI21X1 U344 ( .A(n1047), .B(n994), .C(n186), .Y(n724) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n186) );
  OAI21X1 U346 ( .A(n1048), .B(n994), .C(n187), .Y(n725) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n187) );
  OAI21X1 U348 ( .A(n1049), .B(n994), .C(n188), .Y(n726) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n188) );
  NAND3X1 U350 ( .A(n71), .B(n1013), .C(n967), .Y(n180) );
  OAI21X1 U351 ( .A(n1034), .B(n993), .C(n191), .Y(n727) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n191) );
  OAI21X1 U353 ( .A(n1035), .B(n993), .C(n192), .Y(n728) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n192) );
  OAI21X1 U355 ( .A(n1036), .B(n993), .C(n193), .Y(n729) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n193) );
  OAI21X1 U357 ( .A(n1037), .B(n993), .C(n194), .Y(n730) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n194) );
  OAI21X1 U359 ( .A(n1038), .B(n993), .C(n195), .Y(n731) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n195) );
  OAI21X1 U361 ( .A(n1039), .B(n993), .C(n196), .Y(n732) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n196) );
  OAI21X1 U363 ( .A(n1040), .B(n993), .C(n197), .Y(n733) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n197) );
  OAI21X1 U365 ( .A(n1041), .B(n993), .C(n198), .Y(n734) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n198) );
  NAND3X1 U367 ( .A(n973), .B(n1013), .C(n199), .Y(n190) );
  OAI21X1 U368 ( .A(n1042), .B(n992), .C(n201), .Y(n735) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n201) );
  OAI21X1 U370 ( .A(n1043), .B(n992), .C(n202), .Y(n736) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n202) );
  OAI21X1 U372 ( .A(n1044), .B(n992), .C(n203), .Y(n737) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n203) );
  OAI21X1 U374 ( .A(n1045), .B(n992), .C(n204), .Y(n738) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n204) );
  OAI21X1 U376 ( .A(n1046), .B(n992), .C(n205), .Y(n739) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n205) );
  OAI21X1 U378 ( .A(n1047), .B(n992), .C(n206), .Y(n740) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n206) );
  OAI21X1 U380 ( .A(n1048), .B(n992), .C(n207), .Y(n741) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n207) );
  OAI21X1 U382 ( .A(n1049), .B(n992), .C(n208), .Y(n742) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n208) );
  NAND3X1 U384 ( .A(n91), .B(n1013), .C(n967), .Y(n200) );
  OAI21X1 U385 ( .A(n1034), .B(n991), .C(n210), .Y(n743) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n210) );
  OAI21X1 U387 ( .A(n1035), .B(n991), .C(n211), .Y(n744) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n211) );
  OAI21X1 U389 ( .A(n1036), .B(n991), .C(n212), .Y(n745) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n212) );
  OAI21X1 U391 ( .A(n1037), .B(n991), .C(n213), .Y(n746) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n213) );
  OAI21X1 U393 ( .A(n1038), .B(n991), .C(n214), .Y(n747) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n214) );
  OAI21X1 U395 ( .A(n1039), .B(n991), .C(n215), .Y(n748) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n215) );
  OAI21X1 U397 ( .A(n1040), .B(n991), .C(n216), .Y(n749) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n216) );
  OAI21X1 U399 ( .A(n1041), .B(n991), .C(n217), .Y(n750) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n217) );
  NAND3X1 U401 ( .A(n973), .B(n1013), .C(n218), .Y(n209) );
  OAI21X1 U402 ( .A(n1042), .B(n990), .C(n220), .Y(n751) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n220) );
  OAI21X1 U404 ( .A(n1043), .B(n989), .C(n221), .Y(n752) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n221) );
  OAI21X1 U406 ( .A(n1044), .B(n989), .C(n222), .Y(n753) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n222) );
  OAI21X1 U408 ( .A(n1045), .B(n989), .C(n223), .Y(n754) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n223) );
  OAI21X1 U410 ( .A(n1046), .B(n989), .C(n224), .Y(n755) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n224) );
  OAI21X1 U412 ( .A(n1047), .B(n989), .C(n225), .Y(n756) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n225) );
  OAI21X1 U414 ( .A(n1048), .B(n989), .C(n226), .Y(n757) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n226) );
  OAI21X1 U416 ( .A(n1049), .B(n989), .C(n227), .Y(n758) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n227) );
  NAND3X1 U418 ( .A(n70), .B(n1012), .C(n228), .Y(n219) );
  OAI21X1 U419 ( .A(n1034), .B(n988), .C(n230), .Y(n759) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n230) );
  OAI21X1 U421 ( .A(n1035), .B(n988), .C(n231), .Y(n760) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n231) );
  OAI21X1 U423 ( .A(n1036), .B(n988), .C(n232), .Y(n761) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n232) );
  OAI21X1 U425 ( .A(n1037), .B(n988), .C(n233), .Y(n762) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n233) );
  OAI21X1 U427 ( .A(n1038), .B(n988), .C(n234), .Y(n763) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n234) );
  OAI21X1 U429 ( .A(n1039), .B(n988), .C(n235), .Y(n764) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n235) );
  OAI21X1 U431 ( .A(n1040), .B(n988), .C(n236), .Y(n765) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n236) );
  OAI21X1 U433 ( .A(n1041), .B(n988), .C(n237), .Y(n766) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n237) );
  NAND3X1 U435 ( .A(n973), .B(n1012), .C(n238), .Y(n229) );
  OAI21X1 U436 ( .A(n1042), .B(n987), .C(n240), .Y(n767) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n240) );
  OAI21X1 U438 ( .A(n1043), .B(n986), .C(n241), .Y(n768) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n241) );
  OAI21X1 U440 ( .A(n1044), .B(n986), .C(n242), .Y(n769) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n242) );
  OAI21X1 U442 ( .A(n1045), .B(n986), .C(n243), .Y(n770) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n243) );
  OAI21X1 U444 ( .A(n1046), .B(n986), .C(n244), .Y(n771) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n244) );
  OAI21X1 U446 ( .A(n1047), .B(n986), .C(n245), .Y(n772) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n245) );
  OAI21X1 U448 ( .A(n1048), .B(n986), .C(n246), .Y(n773) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n246) );
  OAI21X1 U450 ( .A(n1049), .B(n986), .C(n247), .Y(n774) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n247) );
  NAND3X1 U452 ( .A(n70), .B(n1012), .C(n248), .Y(n239) );
  OAI21X1 U453 ( .A(n1034), .B(n985), .C(n251), .Y(n775) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n251) );
  OAI21X1 U455 ( .A(n1035), .B(n985), .C(n252), .Y(n776) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n252) );
  OAI21X1 U457 ( .A(n1036), .B(n985), .C(n253), .Y(n777) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n253) );
  OAI21X1 U459 ( .A(n1037), .B(n985), .C(n254), .Y(n778) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n254) );
  OAI21X1 U461 ( .A(n1038), .B(n985), .C(n255), .Y(n779) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n255) );
  OAI21X1 U463 ( .A(n1039), .B(n985), .C(n256), .Y(n780) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n256) );
  OAI21X1 U465 ( .A(n1040), .B(n985), .C(n257), .Y(n781) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n257) );
  OAI21X1 U467 ( .A(n1041), .B(n985), .C(n258), .Y(n782) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n258) );
  NAND3X1 U469 ( .A(n973), .B(n1012), .C(n259), .Y(n250) );
  OAI21X1 U470 ( .A(n1042), .B(n984), .C(n261), .Y(n783) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n261) );
  OAI21X1 U472 ( .A(n1043), .B(n983), .C(n262), .Y(n784) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n262) );
  OAI21X1 U474 ( .A(n1044), .B(n983), .C(n263), .Y(n785) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n263) );
  OAI21X1 U476 ( .A(n1045), .B(n983), .C(n264), .Y(n786) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n264) );
  OAI21X1 U478 ( .A(n1046), .B(n983), .C(n265), .Y(n787) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n265) );
  OAI21X1 U480 ( .A(n1047), .B(n983), .C(n266), .Y(n788) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n266) );
  OAI21X1 U482 ( .A(n1048), .B(n983), .C(n267), .Y(n789) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n267) );
  OAI21X1 U484 ( .A(n1049), .B(n983), .C(n268), .Y(n790) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n268) );
  NAND3X1 U486 ( .A(n111), .B(n1012), .C(n228), .Y(n260) );
  OAI21X1 U487 ( .A(n1034), .B(n982), .C(n270), .Y(n791) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n270) );
  OAI21X1 U489 ( .A(n1035), .B(n982), .C(n271), .Y(n792) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n271) );
  OAI21X1 U491 ( .A(n1036), .B(n982), .C(n272), .Y(n793) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n272) );
  OAI21X1 U493 ( .A(n1037), .B(n982), .C(n273), .Y(n794) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n273) );
  OAI21X1 U495 ( .A(n1038), .B(n982), .C(n274), .Y(n795) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n274) );
  OAI21X1 U497 ( .A(n1039), .B(n982), .C(n275), .Y(n796) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n275) );
  OAI21X1 U499 ( .A(n1040), .B(n982), .C(n276), .Y(n797) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n276) );
  OAI21X1 U501 ( .A(n1041), .B(n982), .C(n277), .Y(n798) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n277) );
  NAND3X1 U503 ( .A(n973), .B(n1012), .C(n278), .Y(n269) );
  OAI21X1 U504 ( .A(n1042), .B(n981), .C(n280), .Y(n799) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n280) );
  OAI21X1 U506 ( .A(n1043), .B(n980), .C(n281), .Y(n800) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n281) );
  OAI21X1 U508 ( .A(n1044), .B(n980), .C(n282), .Y(n801) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n282) );
  OAI21X1 U510 ( .A(n1045), .B(n980), .C(n283), .Y(n802) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n283) );
  OAI21X1 U512 ( .A(n1046), .B(n980), .C(n284), .Y(n803) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n284) );
  OAI21X1 U514 ( .A(n1047), .B(n980), .C(n285), .Y(n804) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n285) );
  OAI21X1 U516 ( .A(n1048), .B(n980), .C(n286), .Y(n805) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n286) );
  OAI21X1 U518 ( .A(n1049), .B(n980), .C(n287), .Y(n806) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n287) );
  NAND3X1 U520 ( .A(n111), .B(n1012), .C(n248), .Y(n279) );
  OAI21X1 U521 ( .A(n1034), .B(n979), .C(n291), .Y(n807) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n291) );
  OAI21X1 U523 ( .A(n1035), .B(n979), .C(n292), .Y(n808) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n292) );
  OAI21X1 U525 ( .A(n1036), .B(n979), .C(n293), .Y(n809) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n293) );
  OAI21X1 U527 ( .A(n1037), .B(n979), .C(n294), .Y(n810) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n294) );
  OAI21X1 U529 ( .A(n1038), .B(n979), .C(n295), .Y(n811) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n295) );
  OAI21X1 U531 ( .A(n1039), .B(n979), .C(n296), .Y(n812) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n296) );
  OAI21X1 U533 ( .A(n1040), .B(n979), .C(n297), .Y(n813) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n297) );
  OAI21X1 U535 ( .A(n1041), .B(n979), .C(n298), .Y(n814) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n298) );
  NAND3X1 U537 ( .A(n973), .B(n1012), .C(n299), .Y(n290) );
  OAI21X1 U538 ( .A(n1042), .B(n978), .C(n301), .Y(n815) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n301) );
  OAI21X1 U540 ( .A(n1043), .B(n978), .C(n302), .Y(n816) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n302) );
  OAI21X1 U542 ( .A(n1044), .B(n978), .C(n303), .Y(n817) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n303) );
  OAI21X1 U544 ( .A(n1045), .B(n978), .C(n304), .Y(n818) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n304) );
  OAI21X1 U546 ( .A(n1046), .B(n978), .C(n305), .Y(n819) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n305) );
  OAI21X1 U548 ( .A(n1047), .B(n978), .C(n306), .Y(n820) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n306) );
  OAI21X1 U550 ( .A(n1048), .B(n978), .C(n307), .Y(n821) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n307) );
  OAI21X1 U552 ( .A(n1049), .B(n978), .C(n308), .Y(n822) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n308) );
  NAND3X1 U554 ( .A(n969), .B(n1012), .C(n228), .Y(n300) );
  OAI21X1 U555 ( .A(n1034), .B(n977), .C(n310), .Y(n823) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n310) );
  OAI21X1 U557 ( .A(n1035), .B(n977), .C(n311), .Y(n824) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n311) );
  OAI21X1 U559 ( .A(n1036), .B(n977), .C(n312), .Y(n825) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n312) );
  OAI21X1 U561 ( .A(n1037), .B(n977), .C(n313), .Y(n826) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n313) );
  OAI21X1 U563 ( .A(n1038), .B(n977), .C(n314), .Y(n827) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n314) );
  OAI21X1 U565 ( .A(n1039), .B(n977), .C(n315), .Y(n828) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n315) );
  OAI21X1 U567 ( .A(n1040), .B(n977), .C(n316), .Y(n829) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n316) );
  OAI21X1 U569 ( .A(n1041), .B(n977), .C(n317), .Y(n830) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n317) );
  NAND3X1 U571 ( .A(n973), .B(n1012), .C(n318), .Y(n309) );
  OAI21X1 U572 ( .A(n1042), .B(n976), .C(n320), .Y(n831) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n320) );
  OAI21X1 U574 ( .A(n1043), .B(n976), .C(n321), .Y(n832) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n321) );
  OAI21X1 U576 ( .A(n1044), .B(n976), .C(n322), .Y(n833) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n322) );
  OAI21X1 U578 ( .A(n1045), .B(n976), .C(n323), .Y(n834) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n323) );
  OAI21X1 U580 ( .A(n1046), .B(n976), .C(n324), .Y(n835) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n324) );
  OAI21X1 U582 ( .A(n1047), .B(n976), .C(n325), .Y(n836) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n325) );
  OAI21X1 U584 ( .A(n1048), .B(n976), .C(n326), .Y(n837) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n326) );
  OAI21X1 U586 ( .A(n1049), .B(n976), .C(n327), .Y(n838) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n327) );
  NAND3X1 U588 ( .A(n969), .B(n1012), .C(n248), .Y(n319) );
  OAI21X1 U590 ( .A(n1034), .B(n975), .C(n330), .Y(n839) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n330) );
  OAI21X1 U592 ( .A(n1035), .B(n975), .C(n331), .Y(n840) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n331) );
  OAI21X1 U594 ( .A(n1036), .B(n975), .C(n332), .Y(n841) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n332) );
  OAI21X1 U596 ( .A(n1037), .B(n975), .C(n333), .Y(n842) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n333) );
  OAI21X1 U598 ( .A(n1038), .B(n975), .C(n334), .Y(n843) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n334) );
  OAI21X1 U600 ( .A(n1039), .B(n975), .C(n335), .Y(n844) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n335) );
  OAI21X1 U602 ( .A(n1040), .B(n975), .C(n336), .Y(n845) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n336) );
  OAI21X1 U604 ( .A(n1041), .B(n975), .C(n337), .Y(n846) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n337) );
  NAND3X1 U606 ( .A(n973), .B(n1012), .C(n338), .Y(n329) );
  OAI21X1 U607 ( .A(n1042), .B(n974), .C(n340), .Y(n847) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n340) );
  OAI21X1 U609 ( .A(n1043), .B(n974), .C(n341), .Y(n848) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n341) );
  OAI21X1 U611 ( .A(n1044), .B(n974), .C(n342), .Y(n849) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n342) );
  OAI21X1 U613 ( .A(n1045), .B(n974), .C(n343), .Y(n850) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n343) );
  OAI21X1 U615 ( .A(n1046), .B(n974), .C(n344), .Y(n851) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n344) );
  OAI21X1 U617 ( .A(n1047), .B(n974), .C(n345), .Y(n852) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n345) );
  OAI21X1 U619 ( .A(n1048), .B(n974), .C(n346), .Y(n853) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n346) );
  OAI21X1 U621 ( .A(n1049), .B(n974), .C(n347), .Y(n854) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n347) );
  NAND3X1 U623 ( .A(n967), .B(n1012), .C(n228), .Y(n339) );
  OAI21X1 U624 ( .A(n1034), .B(n8), .C(n349), .Y(n855) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n349) );
  OAI21X1 U626 ( .A(n1035), .B(n8), .C(n350), .Y(n856) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n350) );
  OAI21X1 U628 ( .A(n1036), .B(n8), .C(n351), .Y(n857) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n351) );
  OAI21X1 U630 ( .A(n1037), .B(n8), .C(n352), .Y(n858) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n352) );
  OAI21X1 U632 ( .A(n1038), .B(n8), .C(n353), .Y(n859) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n353) );
  OAI21X1 U634 ( .A(n1039), .B(n8), .C(n354), .Y(n860) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n354) );
  OAI21X1 U636 ( .A(n1040), .B(n8), .C(n355), .Y(n861) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n355) );
  OAI21X1 U638 ( .A(n1041), .B(n8), .C(n356), .Y(n862) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n356) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n59) );
  OAI21X1 U642 ( .A(n1042), .B(n972), .C(n359), .Y(n863) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n359) );
  OAI21X1 U644 ( .A(n1043), .B(n972), .C(n360), .Y(n864) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n360) );
  OAI21X1 U646 ( .A(n1044), .B(n972), .C(n361), .Y(n865) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n361) );
  OAI21X1 U648 ( .A(n1045), .B(n972), .C(n362), .Y(n866) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n362) );
  OAI21X1 U650 ( .A(n1046), .B(n972), .C(n363), .Y(n867) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n363) );
  OAI21X1 U652 ( .A(n1047), .B(n972), .C(n364), .Y(n868) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n364) );
  OAI21X1 U654 ( .A(n1048), .B(n972), .C(n365), .Y(n869) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n365) );
  OAI21X1 U656 ( .A(n1049), .B(n972), .C(n366), .Y(n870) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n366) );
  NAND3X1 U658 ( .A(n967), .B(n1013), .C(n248), .Y(n358) );
  NOR3X1 U661 ( .A(n370), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n369) );
  NOR3X1 U662 ( .A(n371), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n368) );
  AOI21X1 U663 ( .A(n473), .B(n373), .C(n963), .Y(n1050) );
  OAI21X1 U665 ( .A(rd), .B(n374), .C(wr), .Y(n373) );
  NAND3X1 U667 ( .A(n375), .B(n1029), .C(n376), .Y(n374) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n376) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n375) );
  AOI21X1 U670 ( .A(n460), .B(n378), .C(n1020), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n380), .C(n4), .Y(n378) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n91), .C(\mem<0><1> ), .D(n248), .Y(n383) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n71), .C(\mem<2><1> ), .D(n228), .Y(n382) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n91), .C(\mem<4><1> ), .D(n248), .Y(n385) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n71), .C(\mem<6><1> ), .D(n228), .Y(n384) );
  AOI22X1 U678 ( .A(n288), .B(n893), .C(n249), .D(n933), .Y(n377) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n91), .C(\mem<12><1> ), .D(n248), .Y(
        n389) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n71), .C(\mem<14><1> ), .D(n228), .Y(
        n388) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n91), .C(\mem<8><1> ), .D(n248), .Y(n391) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n71), .C(\mem<10><1> ), .D(n228), .Y(
        n390) );
  AOI21X1 U685 ( .A(n448), .B(n393), .C(n1020), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n940), .B(n395), .C(n950), .Y(n393) );
  AOI21X1 U687 ( .A(n397), .B(n398), .C(n971), .Y(n396) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n91), .C(\mem<0><0> ), .D(n248), .Y(n398) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n71), .C(\mem<2><0> ), .D(n228), .Y(n397) );
  AOI21X1 U690 ( .A(n399), .B(n400), .C(n970), .Y(n394) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n91), .C(\mem<4><0> ), .D(n248), .Y(n400) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n71), .C(\mem<6><0> ), .D(n228), .Y(n399) );
  AOI22X1 U693 ( .A(n288), .B(n891), .C(n249), .D(n931), .Y(n392) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n91), .C(\mem<12><0> ), .D(n248), .Y(
        n404) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n71), .C(\mem<14><0> ), .D(n228), .Y(
        n403) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n91), .C(\mem<8><0> ), .D(n248), .Y(n406) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n71), .C(\mem<10><0> ), .D(n228), .Y(
        n405) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n407) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n199), .C(\mem<19><7> ), .D(n179), .Y(
        n414) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n160), .C(\mem<23><7> ), .D(n140), .Y(
        n413) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n121), .C(\mem<27><7> ), .D(n101), .Y(
        n411) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n81), .C(\mem<31><7> ), .D(n60), .Y(n410) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n357), .C(\mem<3><7> ), .D(n338), .Y(n419) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n318), .C(\mem<7><7> ), .D(n299), .Y(n418) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n278), .C(\mem<11><7> ), .D(n259), .Y(
        n416) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n238), .C(\mem<15><7> ), .D(n218), .Y(
        n415) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n420) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n199), .C(\mem<19><6> ), .D(n179), .Y(
        n427) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n160), .C(\mem<23><6> ), .D(n140), .Y(
        n426) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n121), .C(\mem<27><6> ), .D(n101), .Y(
        n424) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n81), .C(\mem<31><6> ), .D(n60), .Y(n423) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n357), .C(\mem<3><6> ), .D(n338), .Y(n432) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n318), .C(\mem<7><6> ), .D(n299), .Y(n431) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n278), .C(\mem<11><6> ), .D(n259), .Y(
        n429) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n238), .C(\mem<15><6> ), .D(n218), .Y(
        n428) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n433) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n199), .C(\mem<19><5> ), .D(n179), .Y(
        n440) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n160), .C(\mem<23><5> ), .D(n140), .Y(
        n439) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n121), .C(\mem<27><5> ), .D(n101), .Y(
        n437) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n81), .C(\mem<31><5> ), .D(n60), .Y(n436) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n357), .C(\mem<3><5> ), .D(n338), .Y(n445) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n318), .C(\mem<7><5> ), .D(n299), .Y(n444) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n278), .C(\mem<11><5> ), .D(n259), .Y(
        n442) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n238), .C(\mem<15><5> ), .D(n218), .Y(
        n441) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n446) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n199), .C(\mem<19><4> ), .D(n179), .Y(
        n453) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n160), .C(\mem<23><4> ), .D(n140), .Y(
        n452) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n121), .C(\mem<27><4> ), .D(n101), .Y(
        n450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n81), .C(\mem<31><4> ), .D(n60), .Y(n449) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n357), .C(\mem<3><4> ), .D(n338), .Y(n458) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n318), .C(\mem<7><4> ), .D(n299), .Y(n457) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n278), .C(\mem<11><4> ), .D(n259), .Y(
        n455) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n238), .C(\mem<15><4> ), .D(n218), .Y(
        n454) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n459) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n199), .C(\mem<19><3> ), .D(n179), .Y(
        n466) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n160), .C(\mem<23><3> ), .D(n140), .Y(
        n465) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n121), .C(\mem<27><3> ), .D(n101), .Y(
        n463) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n81), .C(\mem<31><3> ), .D(n60), .Y(n462) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n357), .C(\mem<3><3> ), .D(n338), .Y(n471) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n318), .C(\mem<7><3> ), .D(n299), .Y(n470) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n278), .C(\mem<11><3> ), .D(n259), .Y(
        n468) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n238), .C(\mem<15><3> ), .D(n218), .Y(
        n467) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n472) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n199), .C(\mem<19><2> ), .D(n179), .Y(
        n479) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n160), .C(\mem<23><2> ), .D(n140), .Y(
        n478) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n121), .C(\mem<27><2> ), .D(n101), .Y(
        n476) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n81), .C(\mem<31><2> ), .D(n60), .Y(n475) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n357), .C(\mem<3><2> ), .D(n338), .Y(n484) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n318), .C(\mem<7><2> ), .D(n299), .Y(n483) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n278), .C(\mem<11><2> ), .D(n259), .Y(
        n481) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n238), .C(\mem<15><2> ), .D(n218), .Y(
        n480) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n485) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n199), .C(\mem<19><1> ), .D(n179), .Y(
        n492) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n160), .C(\mem<23><1> ), .D(n140), .Y(
        n491) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n121), .C(\mem<27><1> ), .D(n101), .Y(
        n489) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n81), .C(\mem<31><1> ), .D(n60), .Y(n488) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n357), .C(\mem<3><1> ), .D(n338), .Y(n497) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n318), .C(\mem<7><1> ), .D(n299), .Y(n496) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n278), .C(\mem<11><1> ), .D(n259), .Y(
        n494) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n238), .C(\mem<15><1> ), .D(n218), .Y(
        n493) );
  AOI21X1 U777 ( .A(n447), .B(n499), .C(n1020), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n939), .B(n501), .C(n949), .Y(n499) );
  AOI21X1 U779 ( .A(n503), .B(n504), .C(n971), .Y(n502) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n91), .C(\mem<0><7> ), .D(n248), .Y(n504) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n71), .C(\mem<2><7> ), .D(n228), .Y(n503) );
  AOI21X1 U782 ( .A(n505), .B(n506), .C(n970), .Y(n500) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n91), .C(\mem<4><7> ), .D(n248), .Y(n506) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n71), .C(\mem<6><7> ), .D(n228), .Y(n505) );
  AOI22X1 U785 ( .A(n288), .B(n889), .C(n249), .D(n929), .Y(n498) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n91), .C(\mem<12><7> ), .D(n248), .Y(
        n510) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n71), .C(\mem<14><7> ), .D(n228), .Y(
        n509) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n91), .C(\mem<8><7> ), .D(n248), .Y(n512) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n71), .C(\mem<10><7> ), .D(n228), .Y(
        n511) );
  AOI21X1 U792 ( .A(n435), .B(n514), .C(n1020), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n938), .B(n516), .C(n948), .Y(n514) );
  AOI21X1 U794 ( .A(n518), .B(n519), .C(n971), .Y(n517) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n91), .C(\mem<0><6> ), .D(n248), .Y(n519) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n71), .C(\mem<2><6> ), .D(n228), .Y(n518) );
  AOI21X1 U797 ( .A(n520), .B(n521), .C(n970), .Y(n515) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n91), .C(\mem<4><6> ), .D(n248), .Y(n521) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n71), .C(\mem<6><6> ), .D(n228), .Y(n520) );
  AOI22X1 U800 ( .A(n288), .B(n887), .C(n249), .D(n927), .Y(n513) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n91), .C(\mem<12><6> ), .D(n248), .Y(
        n525) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n71), .C(\mem<14><6> ), .D(n228), .Y(
        n524) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n91), .C(\mem<8><6> ), .D(n248), .Y(n527) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n71), .C(\mem<10><6> ), .D(n228), .Y(
        n526) );
  AOI21X1 U807 ( .A(n434), .B(n529), .C(n1020), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n937), .B(n531), .C(n947), .Y(n529) );
  AOI21X1 U809 ( .A(n533), .B(n534), .C(n971), .Y(n532) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n91), .C(\mem<0><5> ), .D(n248), .Y(n534) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n71), .C(\mem<2><5> ), .D(n228), .Y(n533) );
  AOI21X1 U812 ( .A(n535), .B(n536), .C(n970), .Y(n530) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n91), .C(\mem<4><5> ), .D(n248), .Y(n536) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n71), .C(\mem<6><5> ), .D(n228), .Y(n535) );
  AOI22X1 U815 ( .A(n288), .B(n885), .C(n249), .D(n925), .Y(n528) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n91), .C(\mem<12><5> ), .D(n248), .Y(
        n540) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n71), .C(\mem<14><5> ), .D(n228), .Y(
        n539) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n91), .C(\mem<8><5> ), .D(n248), .Y(n542) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n71), .C(\mem<10><5> ), .D(n228), .Y(
        n541) );
  AOI21X1 U822 ( .A(n422), .B(n544), .C(n1020), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n936), .B(n546), .C(n946), .Y(n544) );
  AOI21X1 U824 ( .A(n548), .B(n549), .C(n971), .Y(n547) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n91), .C(\mem<0><4> ), .D(n248), .Y(n549) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n71), .C(\mem<2><4> ), .D(n228), .Y(n548) );
  AOI21X1 U827 ( .A(n550), .B(n551), .C(n970), .Y(n545) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n91), .C(\mem<4><4> ), .D(n248), .Y(n551) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n71), .C(\mem<6><4> ), .D(n228), .Y(n550) );
  AOI22X1 U830 ( .A(n288), .B(n883), .C(n249), .D(n923), .Y(n543) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n91), .C(\mem<12><4> ), .D(n248), .Y(
        n555) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n71), .C(\mem<14><4> ), .D(n228), .Y(
        n554) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n91), .C(\mem<8><4> ), .D(n248), .Y(n557) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n71), .C(\mem<10><4> ), .D(n228), .Y(
        n556) );
  AOI21X1 U837 ( .A(n421), .B(n559), .C(n1020), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n935), .B(n561), .C(n945), .Y(n559) );
  AOI21X1 U839 ( .A(n563), .B(n564), .C(n971), .Y(n562) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n91), .C(\mem<0><3> ), .D(n248), .Y(n564) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n71), .C(\mem<2><3> ), .D(n228), .Y(n563) );
  AOI21X1 U842 ( .A(n565), .B(n566), .C(n970), .Y(n560) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n91), .C(\mem<4><3> ), .D(n248), .Y(n566) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n71), .C(\mem<6><3> ), .D(n228), .Y(n565) );
  AOI22X1 U845 ( .A(n288), .B(n881), .C(n249), .D(n921), .Y(n558) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n91), .C(\mem<12><3> ), .D(n248), .Y(
        n570) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n71), .C(\mem<14><3> ), .D(n228), .Y(
        n569) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n91), .C(\mem<8><3> ), .D(n248), .Y(n572) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n71), .C(\mem<10><3> ), .D(n228), .Y(
        n571) );
  AOI21X1 U852 ( .A(n409), .B(n574), .C(n1020), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n934), .B(n576), .C(n944), .Y(n574) );
  AOI21X1 U854 ( .A(n578), .B(n579), .C(n971), .Y(n577) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n91), .C(\mem<0><2> ), .D(n248), .Y(n579) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n71), .C(\mem<2><2> ), .D(n228), .Y(n578) );
  AOI21X1 U857 ( .A(n580), .B(n581), .C(n970), .Y(n575) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n91), .C(\mem<4><2> ), .D(n248), .Y(n581) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n71), .C(\mem<6><2> ), .D(n228), .Y(n580) );
  AOI22X1 U860 ( .A(n288), .B(n879), .C(n249), .D(n919), .Y(n573) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n91), .C(\mem<12><2> ), .D(n248), .Y(
        n585) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n71), .C(\mem<14><2> ), .D(n228), .Y(
        n584) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n91), .C(\mem<8><2> ), .D(n248), .Y(n587) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n71), .C(\mem<10><2> ), .D(n228), .Y(
        n586) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n588) );
  NOR2X1 U868 ( .A(n1033), .B(\addr_1c<4> ), .Y(n589) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n590) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n199), .C(\mem<19><0> ), .D(n179), .Y(
        n597) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n160), .C(\mem<23><0> ), .D(n140), .Y(
        n596) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n121), .C(\mem<27><0> ), .D(n101), .Y(
        n594) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n81), .C(\mem<31><0> ), .D(n60), .Y(n593) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n357), .C(\mem<3><0> ), .D(n338), .Y(n604) );
  NAND2X1 U877 ( .A(n1031), .B(n1032), .Y(n367) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n318), .C(\mem<7><0> ), .D(n299), .Y(n603) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1032), .Y(n328) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n278), .C(\mem<11><0> ), .D(n259), .Y(
        n601) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n238), .C(\mem<15><0> ), .D(n218), .Y(
        n600) );
  dff_203 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1015) );
  dff_202 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1016) );
  dff_185 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1016)
         );
  dff_186 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1016)
         );
  dff_187 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1016)
         );
  dff_188 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1016)
         );
  dff_189 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1016)
         );
  dff_190 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1016)
         );
  dff_191 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1016)
         );
  dff_192 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1016)
         );
  dff_193 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1015)
         );
  dff_194 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1015)
         );
  dff_195 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1015) );
  dff_196 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1015) );
  dff_197 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1015) );
  dff_169 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1015) );
  dff_170 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1015) );
  dff_171 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1015) );
  dff_172 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1015) );
  dff_173 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1015) );
  dff_174 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1015) );
  dff_175 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1015) );
  dff_176 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1015) );
  dff_177 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1015) );
  dff_178 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1015) );
  dff_179 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1015) );
  dff_180 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1015) );
  dff_181 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1015) );
  dff_182 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1015) );
  dff_183 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1015) );
  dff_184 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1015) );
  dff_153 \reg2[0]  ( .q(\data_out<0> ), .d(n1028), .clk(clk), .rst(n1016) );
  dff_154 \reg2[1]  ( .q(\data_out<1> ), .d(n1027), .clk(clk), .rst(n1016) );
  dff_155 \reg2[2]  ( .q(\data_out<2> ), .d(n1026), .clk(clk), .rst(n1016) );
  dff_156 \reg2[3]  ( .q(\data_out<3> ), .d(n1025), .clk(clk), .rst(n1016) );
  dff_157 \reg2[4]  ( .q(\data_out<4> ), .d(n1024), .clk(clk), .rst(n1016) );
  dff_158 \reg2[5]  ( .q(\data_out<5> ), .d(n1023), .clk(clk), .rst(n1016) );
  dff_159 \reg2[6]  ( .q(\data_out<6> ), .d(n1022), .clk(clk), .rst(n1015) );
  dff_160 \reg2[7]  ( .q(\data_out<7> ), .d(n1021), .clk(clk), .rst(n1015) );
  dff_161 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1015) );
  dff_162 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1015) );
  dff_163 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1015) );
  dff_164 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1015) );
  dff_165 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1015) );
  dff_166 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1015) );
  dff_167 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1015) );
  dff_168 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1015) );
  dff_201 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1015) );
  dff_200 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1015) );
  dff_199 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1015) );
  dff_198 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1016) );
  INVX1 U2 ( .A(wr1), .Y(n1029) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n371) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n357), .Y(n49) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1033) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1032) );
  INVX1 U7 ( .A(\addr_1c<1> ), .Y(n1031) );
  OR2X1 U8 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n370) );
  AND2X1 U23 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n598) );
  AND2X1 U24 ( .A(\addr_1c<3> ), .B(n1030), .Y(n599) );
  AND2X1 U25 ( .A(\addr_1c<0> ), .B(n1033), .Y(n605) );
  AND2X1 U26 ( .A(n1030), .B(n1033), .Y(n606) );
  INVX1 U27 ( .A(\addr_1c<0> ), .Y(n1030) );
  AND2X1 U28 ( .A(\addr_1c<2> ), .B(n1031), .Y(n288) );
  AND2X1 U29 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n249) );
  AND2X1 U35 ( .A(n599), .B(n249), .Y(n81) );
  AND2X1 U36 ( .A(n288), .B(n598), .Y(n101) );
  AND2X1 U37 ( .A(n288), .B(n599), .Y(n121) );
  AND2X1 U38 ( .A(n941), .B(n598), .Y(n140) );
  AND2X1 U39 ( .A(n941), .B(n599), .Y(n160) );
  AND2X1 U40 ( .A(n598), .B(n951), .Y(n179) );
  AND2X1 U41 ( .A(n599), .B(n951), .Y(n199) );
  AND2X1 U42 ( .A(n605), .B(n249), .Y(n218) );
  AND2X1 U43 ( .A(n249), .B(n606), .Y(n238) );
  AND2X1 U44 ( .A(n605), .B(n288), .Y(n259) );
  AND2X1 U46 ( .A(n288), .B(n606), .Y(n278) );
  AND2X1 U47 ( .A(n605), .B(n941), .Y(n299) );
  AND2X1 U48 ( .A(n941), .B(n606), .Y(n318) );
  OR2X1 U49 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U50 ( .A(n605), .B(n951), .Y(n338) );
  OR2X1 U51 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U52 ( .A(n49), .B(\mem<32><0> ), .Y(n395) );
  AND2X1 U53 ( .A(n49), .B(\mem<32><1> ), .Y(n380) );
  AND2X1 U54 ( .A(n49), .B(\mem<32><2> ), .Y(n576) );
  AND2X1 U55 ( .A(n49), .B(\mem<32><3> ), .Y(n561) );
  AND2X1 U56 ( .A(n49), .B(\mem<32><4> ), .Y(n546) );
  AND2X1 U57 ( .A(n49), .B(\mem<32><5> ), .Y(n531) );
  AND2X1 U58 ( .A(n49), .B(\mem<32><6> ), .Y(n516) );
  AND2X1 U59 ( .A(n49), .B(\mem<32><7> ), .Y(n501) );
  INVX1 U60 ( .A(rd1), .Y(n1020) );
  BUFX2 U61 ( .A(n961), .Y(n1010) );
  BUFX2 U62 ( .A(n961), .Y(n1009) );
  BUFX2 U63 ( .A(n960), .Y(n1007) );
  BUFX2 U64 ( .A(n960), .Y(n1006) );
  BUFX2 U65 ( .A(n959), .Y(n1004) );
  BUFX2 U66 ( .A(n959), .Y(n1003) );
  BUFX2 U67 ( .A(n958), .Y(n1001) );
  BUFX2 U68 ( .A(n958), .Y(n1000) );
  BUFX2 U69 ( .A(n957), .Y(n990) );
  BUFX2 U70 ( .A(n957), .Y(n989) );
  BUFX2 U71 ( .A(n956), .Y(n987) );
  BUFX2 U72 ( .A(n956), .Y(n986) );
  BUFX2 U73 ( .A(n955), .Y(n984) );
  BUFX2 U74 ( .A(n955), .Y(n983) );
  BUFX2 U75 ( .A(n954), .Y(n981) );
  BUFX2 U76 ( .A(n954), .Y(n980) );
  INVX1 U77 ( .A(\data_in_1c<0> ), .Y(n1034) );
  INVX1 U78 ( .A(\data_in_1c<1> ), .Y(n1035) );
  INVX1 U79 ( .A(\data_in_1c<2> ), .Y(n1036) );
  INVX1 U80 ( .A(\data_in_1c<3> ), .Y(n1037) );
  INVX1 U81 ( .A(\data_in_1c<4> ), .Y(n1038) );
  INVX1 U82 ( .A(\data_in_1c<5> ), .Y(n1039) );
  INVX1 U83 ( .A(\data_in_1c<6> ), .Y(n1040) );
  INVX1 U84 ( .A(\data_in_1c<7> ), .Y(n1041) );
  INVX1 U85 ( .A(\data_in_1c<8> ), .Y(n1042) );
  INVX1 U86 ( .A(\data_in_1c<9> ), .Y(n1043) );
  INVX1 U87 ( .A(\data_in_1c<10> ), .Y(n1044) );
  INVX1 U88 ( .A(\data_in_1c<11> ), .Y(n1045) );
  INVX1 U89 ( .A(\data_in_1c<12> ), .Y(n1046) );
  INVX1 U90 ( .A(\data_in_1c<13> ), .Y(n1047) );
  INVX1 U91 ( .A(\data_in_1c<14> ), .Y(n1048) );
  INVX1 U92 ( .A(\data_in_1c<15> ), .Y(n1049) );
  INVX1 U93 ( .A(n590), .Y(n1028) );
  INVX1 U129 ( .A(n485), .Y(n1027) );
  INVX1 U589 ( .A(n472), .Y(n1026) );
  INVX1 U640 ( .A(n459), .Y(n1025) );
  INVX1 U659 ( .A(n446), .Y(n1024) );
  INVX1 U660 ( .A(n433), .Y(n1023) );
  INVX1 U664 ( .A(n420), .Y(n1022) );
  INVX1 U666 ( .A(n407), .Y(n1021) );
  INVX2 U672 ( .A(n1017), .Y(n1015) );
  INVX1 U675 ( .A(n48), .Y(n1014) );
  AND2X1 U679 ( .A(wr1), .B(n1017), .Y(n48) );
  INVX1 U682 ( .A(rst), .Y(n1017) );
  AND2X1 U694 ( .A(n249), .B(n964), .Y(n70) );
  INVX1 U697 ( .A(n1014), .Y(n1012) );
  AND2X1 U701 ( .A(n288), .B(n964), .Y(n111) );
  INVX1 U706 ( .A(n1014), .Y(n1013) );
  AND2X1 U712 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U717 ( .A(n1), .Y(n2) );
  AND2X1 U723 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U728 ( .A(n3), .Y(n4) );
  AND2X1 U734 ( .A(n60), .B(n189), .Y(n5) );
  INVX1 U739 ( .A(n5), .Y(n6) );
  AND2X1 U745 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U750 ( .A(n7), .Y(n8) );
  OR2X1 U756 ( .A(n487), .B(n10), .Y(n9) );
  OR2X1 U761 ( .A(n474), .B(n486), .Y(n10) );
  OR2X1 U767 ( .A(n522), .B(n12), .Y(n11) );
  OR2X1 U772 ( .A(n507), .B(n508), .Y(n12) );
  OR2X1 U786 ( .A(n538), .B(n14), .Y(n13) );
  OR2X1 U789 ( .A(n523), .B(n537), .Y(n14) );
  OR2X1 U801 ( .A(n567), .B(n16), .Y(n15) );
  OR2X1 U804 ( .A(n552), .B(n553), .Y(n16) );
  OR2X1 U816 ( .A(n583), .B(n18), .Y(n17) );
  OR2X1 U819 ( .A(n568), .B(n582), .Y(n18) );
  OR2X1 U831 ( .A(n871), .B(n20), .Y(n19) );
  OR2X1 U834 ( .A(n591), .B(n592), .Y(n20) );
  OR2X1 U846 ( .A(n874), .B(n22), .Y(n21) );
  OR2X1 U849 ( .A(n872), .B(n873), .Y(n22) );
  OR2X1 U861 ( .A(n877), .B(n24), .Y(n23) );
  OR2X1 U864 ( .A(n875), .B(n876), .Y(n24) );
  OR2X1 U870 ( .A(n896), .B(n26), .Y(n25) );
  OR2X1 U875 ( .A(n894), .B(n895), .Y(n26) );
  OR2X1 U882 ( .A(n899), .B(n28), .Y(n27) );
  OR2X1 U883 ( .A(n897), .B(n898), .Y(n28) );
  OR2X1 U884 ( .A(n902), .B(n30), .Y(n29) );
  OR2X1 U885 ( .A(n900), .B(n901), .Y(n30) );
  OR2X1 U886 ( .A(n905), .B(n32), .Y(n31) );
  OR2X1 U887 ( .A(n903), .B(n904), .Y(n32) );
  OR2X1 U888 ( .A(n908), .B(n34), .Y(n33) );
  OR2X1 U889 ( .A(n906), .B(n907), .Y(n34) );
  OR2X1 U890 ( .A(n911), .B(n36), .Y(n35) );
  OR2X1 U891 ( .A(n909), .B(n910), .Y(n36) );
  OR2X1 U892 ( .A(n914), .B(n38), .Y(n37) );
  OR2X1 U893 ( .A(n912), .B(n913), .Y(n38) );
  OR2X1 U894 ( .A(n917), .B(n150), .Y(n50) );
  OR2X1 U895 ( .A(n915), .B(n916), .Y(n150) );
  AND2X1 U896 ( .A(n973), .B(n48), .Y(n189) );
  AND2X1 U897 ( .A(n48), .B(n357), .Y(n289) );
  INVX1 U898 ( .A(n1017), .Y(n1016) );
  AND2X1 U899 ( .A(n941), .B(n943), .Y(n348) );
  INVX1 U900 ( .A(n348), .Y(n372) );
  AND2X1 U901 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U902 ( .A(n379), .Y(n381) );
  AND2X1 U903 ( .A(n941), .B(n942), .Y(n386) );
  INVX1 U904 ( .A(n386), .Y(n387) );
  AND2X1 U905 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U906 ( .A(n401), .Y(n402) );
  BUFX2 U907 ( .A(n1050), .Y(err) );
  BUFX2 U908 ( .A(n573), .Y(n409) );
  BUFX2 U909 ( .A(n558), .Y(n421) );
  BUFX2 U910 ( .A(n543), .Y(n422) );
  BUFX2 U911 ( .A(n528), .Y(n434) );
  BUFX2 U912 ( .A(n513), .Y(n435) );
  BUFX2 U913 ( .A(n498), .Y(n447) );
  BUFX2 U914 ( .A(n392), .Y(n448) );
  BUFX2 U915 ( .A(n377), .Y(n460) );
  AND2X2 U916 ( .A(rd), .B(n374), .Y(n461) );
  INVX1 U917 ( .A(n461), .Y(n473) );
  INVX1 U918 ( .A(n602), .Y(n474) );
  INVX1 U919 ( .A(n601), .Y(n486) );
  INVX1 U920 ( .A(n600), .Y(n487) );
  INVX1 U921 ( .A(n495), .Y(n507) );
  INVX1 U922 ( .A(n494), .Y(n508) );
  INVX1 U923 ( .A(n493), .Y(n522) );
  INVX1 U924 ( .A(n482), .Y(n523) );
  INVX1 U925 ( .A(n481), .Y(n537) );
  INVX1 U926 ( .A(n480), .Y(n538) );
  INVX1 U927 ( .A(n469), .Y(n552) );
  INVX1 U928 ( .A(n468), .Y(n553) );
  INVX1 U929 ( .A(n467), .Y(n567) );
  INVX1 U930 ( .A(n456), .Y(n568) );
  INVX1 U931 ( .A(n455), .Y(n582) );
  INVX1 U932 ( .A(n454), .Y(n583) );
  INVX1 U933 ( .A(n443), .Y(n591) );
  INVX1 U934 ( .A(n442), .Y(n592) );
  INVX1 U935 ( .A(n441), .Y(n871) );
  INVX1 U936 ( .A(n430), .Y(n872) );
  INVX1 U937 ( .A(n429), .Y(n873) );
  INVX1 U938 ( .A(n428), .Y(n874) );
  INVX1 U939 ( .A(n417), .Y(n875) );
  INVX1 U940 ( .A(n416), .Y(n876) );
  INVX1 U941 ( .A(n415), .Y(n877) );
  AND2X2 U942 ( .A(n586), .B(n587), .Y(n878) );
  INVX1 U943 ( .A(n878), .Y(n879) );
  AND2X2 U944 ( .A(n571), .B(n572), .Y(n880) );
  INVX1 U945 ( .A(n880), .Y(n881) );
  AND2X2 U946 ( .A(n556), .B(n557), .Y(n882) );
  INVX1 U947 ( .A(n882), .Y(n883) );
  AND2X2 U948 ( .A(n541), .B(n542), .Y(n884) );
  INVX1 U949 ( .A(n884), .Y(n885) );
  AND2X2 U950 ( .A(n526), .B(n527), .Y(n886) );
  INVX1 U951 ( .A(n886), .Y(n887) );
  AND2X2 U952 ( .A(n511), .B(n512), .Y(n888) );
  INVX1 U953 ( .A(n888), .Y(n889) );
  AND2X2 U954 ( .A(n405), .B(n406), .Y(n890) );
  INVX1 U955 ( .A(n890), .Y(n891) );
  AND2X2 U956 ( .A(n390), .B(n391), .Y(n892) );
  INVX1 U957 ( .A(n892), .Y(n893) );
  INVX1 U958 ( .A(n595), .Y(n894) );
  INVX1 U959 ( .A(n594), .Y(n895) );
  INVX1 U960 ( .A(n593), .Y(n896) );
  INVX1 U961 ( .A(n490), .Y(n897) );
  INVX1 U962 ( .A(n489), .Y(n898) );
  INVX1 U963 ( .A(n488), .Y(n899) );
  INVX1 U964 ( .A(n477), .Y(n900) );
  INVX1 U965 ( .A(n476), .Y(n901) );
  INVX1 U966 ( .A(n475), .Y(n902) );
  INVX1 U967 ( .A(n464), .Y(n903) );
  INVX1 U968 ( .A(n463), .Y(n904) );
  INVX1 U969 ( .A(n462), .Y(n905) );
  INVX1 U970 ( .A(n451), .Y(n906) );
  INVX1 U971 ( .A(n450), .Y(n907) );
  INVX1 U972 ( .A(n449), .Y(n908) );
  INVX1 U973 ( .A(n438), .Y(n909) );
  INVX1 U974 ( .A(n437), .Y(n910) );
  INVX1 U975 ( .A(n436), .Y(n911) );
  INVX1 U976 ( .A(n425), .Y(n912) );
  INVX1 U977 ( .A(n424), .Y(n913) );
  INVX1 U978 ( .A(n423), .Y(n914) );
  INVX1 U979 ( .A(n412), .Y(n915) );
  INVX1 U980 ( .A(n411), .Y(n916) );
  INVX1 U981 ( .A(n410), .Y(n917) );
  AND2X2 U982 ( .A(n584), .B(n585), .Y(n918) );
  INVX1 U983 ( .A(n918), .Y(n919) );
  AND2X2 U984 ( .A(n569), .B(n570), .Y(n920) );
  INVX1 U985 ( .A(n920), .Y(n921) );
  AND2X2 U986 ( .A(n554), .B(n555), .Y(n922) );
  INVX1 U987 ( .A(n922), .Y(n923) );
  AND2X2 U988 ( .A(n539), .B(n540), .Y(n924) );
  INVX1 U989 ( .A(n924), .Y(n925) );
  AND2X2 U990 ( .A(n524), .B(n525), .Y(n926) );
  INVX1 U991 ( .A(n926), .Y(n927) );
  AND2X2 U992 ( .A(n509), .B(n510), .Y(n928) );
  INVX1 U993 ( .A(n928), .Y(n929) );
  AND2X2 U994 ( .A(n403), .B(n404), .Y(n930) );
  INVX1 U995 ( .A(n930), .Y(n931) );
  AND2X2 U996 ( .A(n388), .B(n389), .Y(n932) );
  INVX1 U997 ( .A(n932), .Y(n933) );
  BUFX2 U998 ( .A(n575), .Y(n934) );
  BUFX2 U999 ( .A(n560), .Y(n935) );
  BUFX2 U1000 ( .A(n545), .Y(n936) );
  BUFX2 U1001 ( .A(n530), .Y(n937) );
  BUFX2 U1002 ( .A(n515), .Y(n938) );
  BUFX2 U1003 ( .A(n500), .Y(n939) );
  BUFX2 U1004 ( .A(n394), .Y(n940) );
  INVX1 U1005 ( .A(n970), .Y(n941) );
  INVX1 U1006 ( .A(n385), .Y(n942) );
  INVX1 U1007 ( .A(n384), .Y(n943) );
  BUFX2 U1008 ( .A(n328), .Y(n970) );
  BUFX2 U1009 ( .A(n577), .Y(n944) );
  BUFX2 U1010 ( .A(n562), .Y(n945) );
  BUFX2 U1011 ( .A(n547), .Y(n946) );
  BUFX2 U1012 ( .A(n532), .Y(n947) );
  BUFX2 U1013 ( .A(n517), .Y(n948) );
  BUFX2 U1014 ( .A(n502), .Y(n949) );
  BUFX2 U1015 ( .A(n396), .Y(n950) );
  INVX1 U1016 ( .A(n971), .Y(n951) );
  INVX1 U1017 ( .A(n383), .Y(n952) );
  INVX1 U1018 ( .A(n382), .Y(n953) );
  BUFX2 U1019 ( .A(n367), .Y(n971) );
  BUFX2 U1020 ( .A(n358), .Y(n972) );
  BUFX2 U1021 ( .A(n339), .Y(n974) );
  BUFX2 U1022 ( .A(n329), .Y(n975) );
  BUFX2 U1023 ( .A(n319), .Y(n976) );
  BUFX2 U1024 ( .A(n309), .Y(n977) );
  BUFX2 U1025 ( .A(n300), .Y(n978) );
  BUFX2 U1026 ( .A(n290), .Y(n979) );
  BUFX2 U1027 ( .A(n269), .Y(n982) );
  BUFX2 U1028 ( .A(n250), .Y(n985) );
  BUFX2 U1029 ( .A(n229), .Y(n988) );
  BUFX2 U1030 ( .A(n209), .Y(n991) );
  BUFX2 U1031 ( .A(n200), .Y(n992) );
  BUFX2 U1032 ( .A(n190), .Y(n993) );
  BUFX2 U1033 ( .A(n180), .Y(n994) );
  BUFX2 U1034 ( .A(n170), .Y(n995) );
  BUFX2 U1035 ( .A(n161), .Y(n996) );
  BUFX2 U1036 ( .A(n151), .Y(n997) );
  BUFX2 U1037 ( .A(n141), .Y(n998) );
  BUFX2 U1038 ( .A(n131), .Y(n999) );
  BUFX2 U1039 ( .A(n112), .Y(n1002) );
  BUFX2 U1040 ( .A(n92), .Y(n1005) );
  BUFX2 U1041 ( .A(n72), .Y(n1008) );
  BUFX2 U1042 ( .A(n59), .Y(n973) );
  AND2X1 U1043 ( .A(n249), .B(n598), .Y(n60) );
  BUFX2 U1044 ( .A(n39), .Y(n1011) );
  BUFX2 U1045 ( .A(n279), .Y(n954) );
  BUFX2 U1046 ( .A(n260), .Y(n955) );
  BUFX2 U1047 ( .A(n239), .Y(n956) );
  BUFX2 U1048 ( .A(n219), .Y(n957) );
  BUFX2 U1049 ( .A(n122), .Y(n958) );
  BUFX2 U1050 ( .A(n102), .Y(n959) );
  BUFX2 U1051 ( .A(n82), .Y(n960) );
  BUFX2 U1052 ( .A(n61), .Y(n961) );
  AND2X1 U1053 ( .A(enable), .B(n1017), .Y(n962) );
  INVX1 U1054 ( .A(n962), .Y(n963) );
  AND2X1 U1055 ( .A(n368), .B(n369), .Y(n964) );
  INVX1 U1056 ( .A(n964), .Y(n965) );
  INVX1 U1057 ( .A(n966), .Y(n967) );
  INVX1 U1058 ( .A(n968), .Y(n969) );
  AND2X1 U1059 ( .A(n951), .B(n606), .Y(n357) );
  INVX1 U1060 ( .A(rd), .Y(n1018) );
  INVX1 U1061 ( .A(wr), .Y(n1019) );
endmodule


module final_memory_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1839, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1047), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1048), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1049), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1050), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1051), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1052), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1053), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1054), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1055), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1056), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1057), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1058), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1059), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1060), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1061), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1062), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1063), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1064), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1065), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1066), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1067), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1068), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1069), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1070), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1071), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1072), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1073), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1074), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1075), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1076), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1077), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1078), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1079), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1080), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1081), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1082), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1083), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1084), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1085), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1086), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1087), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1088), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1089), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1090), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1091), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1092), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1093), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1094), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1095), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1096), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1097), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1098), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1099), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1100), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1101), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1102), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1103), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1104), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1105), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1106), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1107), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1108), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1109), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1110), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1111), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1112), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1113), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1114), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1115), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1116), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1117), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1118), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1119), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1120), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1121), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1122), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1123), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1124), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1125), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1126), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1127), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1128), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1129), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1130), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1131), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1132), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1133), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1134), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1135), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1136), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1137), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1138), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1139), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1140), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1141), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1142), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1143), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1144), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1145), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1146), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1147), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1148), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1149), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1150), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1151), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1152), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1153), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1154), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1155), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1156), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1157), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1158), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1159), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1160), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1161), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1162), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1163), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1164), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1165), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1166), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1167), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1168), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1169), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1170), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1171), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1172), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1173), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1174), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1175), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1176), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1177), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1178), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1179), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1180), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1181), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1182), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1183), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1184), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1185), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1186), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1187), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1188), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1189), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1190), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1191), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1192), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1193), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1194), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1195), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1196), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1197), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1198), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1199), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1200), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1201), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1202), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1203), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1204), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1205), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1206), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1207), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1208), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1209), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1210), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1211), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1212), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1213), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1214), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1215), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1216), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1217), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1218), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1219), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1220), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1221), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1222), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1223), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1224), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1225), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1226), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1227), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1228), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1229), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1230), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1231), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1232), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1233), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1234), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1235), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1236), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1237), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1238), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1239), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1240), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1241), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1242), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1243), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1244), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1245), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1246), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1247), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1248), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1249), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1250), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1251), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1252), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1253), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1254), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1255), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1256), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1257), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1258), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1259), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1260), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1261), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1262), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1263), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1264), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1265), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1266), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1267), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1268), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1269), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1270), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1271), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1272), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1273), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1274), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1275), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1276), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1277), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1278), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1279), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1280), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1281), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1282), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1283), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1284), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1285), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1286), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1287), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1288), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1289), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1290), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1291), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1292), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1293), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1294), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1295), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1296), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1297), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1298), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1299), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1300), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1301), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1302), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1303), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1304), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1305), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1306), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1307), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1308), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1309), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1310), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1478), .B(n1477), .Y(n1479) );
  AND2X2 U10 ( .A(n1473), .B(n1472), .Y(n1474) );
  AND2X2 U11 ( .A(n1467), .B(n1466), .Y(n1468) );
  AND2X2 U12 ( .A(n1462), .B(n1461), .Y(n1463) );
  AND2X2 U13 ( .A(n1456), .B(n1455), .Y(n1457) );
  AND2X2 U14 ( .A(n1451), .B(n1450), .Y(n1452) );
  AND2X2 U15 ( .A(n1445), .B(n1444), .Y(n1446) );
  AND2X2 U16 ( .A(n1440), .B(n1439), .Y(n1441) );
  AND2X2 U17 ( .A(n1434), .B(n1433), .Y(n1435) );
  AND2X2 U18 ( .A(n1429), .B(n1428), .Y(n1430) );
  AND2X2 U19 ( .A(n1423), .B(n1422), .Y(n1424) );
  AND2X2 U20 ( .A(n1418), .B(n1417), .Y(n1419) );
  AND2X2 U21 ( .A(n1412), .B(n1411), .Y(n1413) );
  AND2X2 U22 ( .A(n1407), .B(n1406), .Y(n1408) );
  AND2X2 U30 ( .A(n1327), .B(n1027), .Y(n1632) );
  AND2X2 U31 ( .A(n1326), .B(n1027), .Y(n1787) );
  AND2X2 U32 ( .A(n1327), .B(\addr_1c<0> ), .Y(n1652) );
  AND2X2 U33 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1807) );
  AND2X2 U34 ( .A(n1321), .B(n1320), .Y(n1322) );
  AND2X2 U45 ( .A(n1314), .B(n1313), .Y(n1315) );
  NOR3X1 U94 ( .A(n1024), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1023), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1039), .C(n1837), .Y(n1310) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1837) );
  OAI21X1 U98 ( .A(n1011), .B(n1040), .C(n1836), .Y(n1309) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1836) );
  OAI21X1 U100 ( .A(n1011), .B(n1041), .C(n1835), .Y(n1308) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1835) );
  OAI21X1 U102 ( .A(n1011), .B(n1042), .C(n1834), .Y(n1307) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1834) );
  OAI21X1 U104 ( .A(n1011), .B(n1043), .C(n1833), .Y(n1306) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1833) );
  OAI21X1 U106 ( .A(n1011), .B(n1044), .C(n1832), .Y(n1305) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1832) );
  OAI21X1 U108 ( .A(n1011), .B(n1045), .C(n1831), .Y(n1304) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1831) );
  OAI21X1 U110 ( .A(n1011), .B(n1046), .C(n1830), .Y(n1303) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1830) );
  NAND3X1 U112 ( .A(n1829), .B(n1828), .C(n964), .Y(n1838) );
  OAI21X1 U113 ( .A(n6), .B(n1031), .C(n1827), .Y(n1302) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1827) );
  OAI21X1 U115 ( .A(n6), .B(n1032), .C(n1826), .Y(n1301) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1826) );
  OAI21X1 U117 ( .A(n6), .B(n1033), .C(n1825), .Y(n1300) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1825) );
  OAI21X1 U119 ( .A(n6), .B(n1034), .C(n1824), .Y(n1299) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1824) );
  OAI21X1 U121 ( .A(n6), .B(n1035), .C(n1823), .Y(n1298) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1823) );
  OAI21X1 U123 ( .A(n6), .B(n1036), .C(n1822), .Y(n1297) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1822) );
  OAI21X1 U125 ( .A(n6), .B(n1037), .C(n1821), .Y(n1296) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1821) );
  OAI21X1 U127 ( .A(n6), .B(n1038), .C(n1820), .Y(n1295) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1820) );
  OAI21X1 U130 ( .A(n1039), .B(n1010), .C(n1816), .Y(n1294) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1816) );
  OAI21X1 U132 ( .A(n1040), .B(n1009), .C(n1815), .Y(n1293) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1815) );
  OAI21X1 U134 ( .A(n1041), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1814) );
  OAI21X1 U136 ( .A(n1042), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1813) );
  OAI21X1 U138 ( .A(n1043), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1812) );
  OAI21X1 U140 ( .A(n1044), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1811) );
  OAI21X1 U142 ( .A(n1045), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1810) );
  OAI21X1 U144 ( .A(n1046), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1809) );
  NAND3X1 U146 ( .A(n1808), .B(n1829), .C(n1807), .Y(n1817) );
  OAI21X1 U147 ( .A(n1031), .B(n1008), .C(n1805), .Y(n1286) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1805) );
  OAI21X1 U149 ( .A(n1032), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1804) );
  OAI21X1 U151 ( .A(n1033), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1803) );
  OAI21X1 U153 ( .A(n1034), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1802) );
  OAI21X1 U155 ( .A(n1035), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1801) );
  OAI21X1 U157 ( .A(n1036), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1800) );
  OAI21X1 U159 ( .A(n1037), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1799) );
  OAI21X1 U161 ( .A(n1038), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1798) );
  NAND3X1 U163 ( .A(n973), .B(n1829), .C(n1797), .Y(n1806) );
  OAI21X1 U164 ( .A(n1039), .B(n1007), .C(n1795), .Y(n1278) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1795) );
  OAI21X1 U166 ( .A(n1040), .B(n1006), .C(n1794), .Y(n1277) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1794) );
  OAI21X1 U168 ( .A(n1041), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1793) );
  OAI21X1 U170 ( .A(n1042), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1792) );
  OAI21X1 U172 ( .A(n1043), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1791) );
  OAI21X1 U174 ( .A(n1044), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1790) );
  OAI21X1 U176 ( .A(n1045), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1789) );
  OAI21X1 U178 ( .A(n1046), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1788) );
  NAND3X1 U180 ( .A(n1808), .B(n1829), .C(n1787), .Y(n1796) );
  OAI21X1 U181 ( .A(n1031), .B(n1005), .C(n1785), .Y(n1270) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1785) );
  OAI21X1 U183 ( .A(n1032), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1784) );
  OAI21X1 U185 ( .A(n1033), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1783) );
  OAI21X1 U187 ( .A(n1034), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1782) );
  OAI21X1 U189 ( .A(n1035), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1781) );
  OAI21X1 U191 ( .A(n1036), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1780) );
  OAI21X1 U193 ( .A(n1037), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1779) );
  OAI21X1 U195 ( .A(n1038), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1778) );
  NAND3X1 U197 ( .A(n973), .B(n1829), .C(n1777), .Y(n1786) );
  OAI21X1 U198 ( .A(n1039), .B(n1004), .C(n1775), .Y(n1262) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1775) );
  OAI21X1 U200 ( .A(n1040), .B(n1003), .C(n1774), .Y(n1261) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1774) );
  OAI21X1 U202 ( .A(n1041), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1773) );
  OAI21X1 U204 ( .A(n1042), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1772) );
  OAI21X1 U206 ( .A(n1043), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1771) );
  OAI21X1 U208 ( .A(n1044), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1770) );
  OAI21X1 U210 ( .A(n1045), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1769) );
  OAI21X1 U212 ( .A(n1046), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1768) );
  NAND3X1 U214 ( .A(n1807), .B(n1829), .C(n1767), .Y(n1776) );
  OAI21X1 U215 ( .A(n1031), .B(n1002), .C(n1765), .Y(n1254) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1765) );
  OAI21X1 U217 ( .A(n1032), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1764) );
  OAI21X1 U219 ( .A(n1033), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1763) );
  OAI21X1 U221 ( .A(n1034), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1762) );
  OAI21X1 U223 ( .A(n1035), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1761) );
  OAI21X1 U225 ( .A(n1036), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1760) );
  OAI21X1 U227 ( .A(n1037), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1759) );
  OAI21X1 U229 ( .A(n1038), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1758) );
  NAND3X1 U231 ( .A(n973), .B(n1829), .C(n1757), .Y(n1766) );
  OAI21X1 U232 ( .A(n1039), .B(n1001), .C(n1755), .Y(n1246) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1755) );
  OAI21X1 U234 ( .A(n1040), .B(n1000), .C(n1754), .Y(n1245) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1754) );
  OAI21X1 U236 ( .A(n1041), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1753) );
  OAI21X1 U238 ( .A(n1042), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1752) );
  OAI21X1 U240 ( .A(n1043), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1751) );
  OAI21X1 U242 ( .A(n1044), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1750) );
  OAI21X1 U244 ( .A(n1045), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1749) );
  OAI21X1 U246 ( .A(n1046), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1748) );
  NAND3X1 U248 ( .A(n1787), .B(n1829), .C(n1767), .Y(n1756) );
  OAI21X1 U249 ( .A(n1031), .B(n999), .C(n1746), .Y(n1238) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1746) );
  OAI21X1 U251 ( .A(n1032), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1745) );
  OAI21X1 U253 ( .A(n1033), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1744) );
  OAI21X1 U255 ( .A(n1034), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1743) );
  OAI21X1 U257 ( .A(n1035), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1742) );
  OAI21X1 U259 ( .A(n1036), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1741) );
  OAI21X1 U261 ( .A(n1037), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1740) );
  OAI21X1 U263 ( .A(n1038), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1739) );
  NAND3X1 U265 ( .A(n973), .B(n1829), .C(n1738), .Y(n1747) );
  OAI21X1 U266 ( .A(n1039), .B(n998), .C(n1736), .Y(n1230) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1736) );
  OAI21X1 U268 ( .A(n1040), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1735) );
  OAI21X1 U270 ( .A(n1041), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1734) );
  OAI21X1 U272 ( .A(n1042), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1733) );
  OAI21X1 U274 ( .A(n1043), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1732) );
  OAI21X1 U276 ( .A(n1044), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1731) );
  OAI21X1 U278 ( .A(n1045), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1730) );
  OAI21X1 U280 ( .A(n1046), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1729) );
  NAND3X1 U282 ( .A(n1807), .B(n1829), .C(n969), .Y(n1737) );
  OAI21X1 U283 ( .A(n1031), .B(n997), .C(n1727), .Y(n1222) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1727) );
  OAI21X1 U285 ( .A(n1032), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1726) );
  OAI21X1 U287 ( .A(n1033), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1725) );
  OAI21X1 U289 ( .A(n1034), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1724) );
  OAI21X1 U291 ( .A(n1035), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1723) );
  OAI21X1 U293 ( .A(n1036), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1722) );
  OAI21X1 U295 ( .A(n1037), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1721) );
  OAI21X1 U297 ( .A(n1038), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1720) );
  NAND3X1 U299 ( .A(n973), .B(n1829), .C(n1719), .Y(n1728) );
  OAI21X1 U300 ( .A(n1039), .B(n996), .C(n1717), .Y(n1214) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1717) );
  OAI21X1 U302 ( .A(n1040), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1716) );
  OAI21X1 U304 ( .A(n1041), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1715) );
  OAI21X1 U306 ( .A(n1042), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1714) );
  OAI21X1 U308 ( .A(n1043), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1713) );
  OAI21X1 U310 ( .A(n1044), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1712) );
  OAI21X1 U312 ( .A(n1045), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1711) );
  OAI21X1 U314 ( .A(n1046), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1710) );
  NAND3X1 U316 ( .A(n1787), .B(n1829), .C(n969), .Y(n1718) );
  OAI21X1 U317 ( .A(n1031), .B(n995), .C(n1708), .Y(n1206) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1708) );
  OAI21X1 U319 ( .A(n1032), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1707) );
  OAI21X1 U321 ( .A(n1033), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1706) );
  OAI21X1 U323 ( .A(n1034), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1705) );
  OAI21X1 U325 ( .A(n1035), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1704) );
  OAI21X1 U327 ( .A(n1036), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1703) );
  OAI21X1 U329 ( .A(n1037), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1702) );
  OAI21X1 U331 ( .A(n1038), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1701) );
  NAND3X1 U333 ( .A(n973), .B(n1829), .C(n1700), .Y(n1709) );
  OAI21X1 U334 ( .A(n1039), .B(n994), .C(n1698), .Y(n1198) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1698) );
  OAI21X1 U336 ( .A(n1040), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1697) );
  OAI21X1 U338 ( .A(n1041), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1696) );
  OAI21X1 U340 ( .A(n1042), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1695) );
  OAI21X1 U342 ( .A(n1043), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1694) );
  OAI21X1 U344 ( .A(n1044), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1693) );
  OAI21X1 U346 ( .A(n1045), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1692) );
  OAI21X1 U348 ( .A(n1046), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1691) );
  NAND3X1 U350 ( .A(n1807), .B(n1829), .C(n967), .Y(n1699) );
  OAI21X1 U351 ( .A(n1031), .B(n993), .C(n1689), .Y(n1190) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1689) );
  OAI21X1 U353 ( .A(n1032), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1688) );
  OAI21X1 U355 ( .A(n1033), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1687) );
  OAI21X1 U357 ( .A(n1034), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1686) );
  OAI21X1 U359 ( .A(n1035), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1685) );
  OAI21X1 U361 ( .A(n1036), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1684) );
  OAI21X1 U363 ( .A(n1037), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1683) );
  OAI21X1 U365 ( .A(n1038), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1682) );
  NAND3X1 U367 ( .A(n973), .B(n1829), .C(n1681), .Y(n1690) );
  OAI21X1 U368 ( .A(n1039), .B(n992), .C(n1679), .Y(n1182) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1679) );
  OAI21X1 U370 ( .A(n1040), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1678) );
  OAI21X1 U372 ( .A(n1041), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1677) );
  OAI21X1 U374 ( .A(n1042), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1676) );
  OAI21X1 U376 ( .A(n1043), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1675) );
  OAI21X1 U378 ( .A(n1044), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1674) );
  OAI21X1 U380 ( .A(n1045), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1673) );
  OAI21X1 U382 ( .A(n1046), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1672) );
  NAND3X1 U384 ( .A(n1787), .B(n1829), .C(n967), .Y(n1680) );
  OAI21X1 U385 ( .A(n1031), .B(n991), .C(n1670), .Y(n1174) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1670) );
  OAI21X1 U387 ( .A(n1032), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1669) );
  OAI21X1 U389 ( .A(n1033), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1668) );
  OAI21X1 U391 ( .A(n1034), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1667) );
  OAI21X1 U393 ( .A(n1035), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1666) );
  OAI21X1 U395 ( .A(n1036), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1665) );
  OAI21X1 U397 ( .A(n1037), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1664) );
  OAI21X1 U399 ( .A(n1038), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1663) );
  NAND3X1 U401 ( .A(n973), .B(n1829), .C(n1662), .Y(n1671) );
  OAI21X1 U402 ( .A(n1039), .B(n990), .C(n1660), .Y(n1166) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1660) );
  OAI21X1 U404 ( .A(n1040), .B(n989), .C(n1659), .Y(n1165) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1659) );
  OAI21X1 U406 ( .A(n1041), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1658) );
  OAI21X1 U408 ( .A(n1042), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1657) );
  OAI21X1 U410 ( .A(n1043), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1656) );
  OAI21X1 U412 ( .A(n1044), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1655) );
  OAI21X1 U414 ( .A(n1045), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1654) );
  OAI21X1 U416 ( .A(n1046), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1653) );
  NAND3X1 U418 ( .A(n1808), .B(n1829), .C(n1652), .Y(n1661) );
  OAI21X1 U419 ( .A(n1031), .B(n988), .C(n1650), .Y(n1158) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1650) );
  OAI21X1 U421 ( .A(n1032), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1649) );
  OAI21X1 U423 ( .A(n1033), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1648) );
  OAI21X1 U425 ( .A(n1034), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1647) );
  OAI21X1 U427 ( .A(n1035), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1646) );
  OAI21X1 U429 ( .A(n1036), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1645) );
  OAI21X1 U431 ( .A(n1037), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1644) );
  OAI21X1 U433 ( .A(n1038), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1643) );
  NAND3X1 U435 ( .A(n973), .B(n1829), .C(n1642), .Y(n1651) );
  OAI21X1 U436 ( .A(n1039), .B(n987), .C(n1640), .Y(n1150) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1640) );
  OAI21X1 U438 ( .A(n1040), .B(n986), .C(n1639), .Y(n1149) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1639) );
  OAI21X1 U440 ( .A(n1041), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1638) );
  OAI21X1 U442 ( .A(n1042), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1637) );
  OAI21X1 U444 ( .A(n1043), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1636) );
  OAI21X1 U446 ( .A(n1044), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1635) );
  OAI21X1 U448 ( .A(n1045), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1634) );
  OAI21X1 U450 ( .A(n1046), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1633) );
  NAND3X1 U452 ( .A(n1808), .B(n1829), .C(n1632), .Y(n1641) );
  OAI21X1 U453 ( .A(n1031), .B(n985), .C(n1629), .Y(n1142) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1629) );
  OAI21X1 U455 ( .A(n1032), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1628) );
  OAI21X1 U457 ( .A(n1033), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1627) );
  OAI21X1 U459 ( .A(n1034), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1626) );
  OAI21X1 U461 ( .A(n1035), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1625) );
  OAI21X1 U463 ( .A(n1036), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1624) );
  OAI21X1 U465 ( .A(n1037), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1623) );
  OAI21X1 U467 ( .A(n1038), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1622) );
  NAND3X1 U469 ( .A(n973), .B(n1829), .C(n1621), .Y(n1630) );
  OAI21X1 U470 ( .A(n1039), .B(n984), .C(n1619), .Y(n1134) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1619) );
  OAI21X1 U472 ( .A(n1040), .B(n983), .C(n1618), .Y(n1133) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1618) );
  OAI21X1 U474 ( .A(n1041), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1617) );
  OAI21X1 U476 ( .A(n1042), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1616) );
  OAI21X1 U478 ( .A(n1043), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1615) );
  OAI21X1 U480 ( .A(n1044), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1614) );
  OAI21X1 U482 ( .A(n1045), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1613) );
  OAI21X1 U484 ( .A(n1046), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1612) );
  NAND3X1 U486 ( .A(n1767), .B(n1829), .C(n1652), .Y(n1620) );
  OAI21X1 U487 ( .A(n1031), .B(n982), .C(n1610), .Y(n1126) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1610) );
  OAI21X1 U489 ( .A(n1032), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1609) );
  OAI21X1 U491 ( .A(n1033), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1608) );
  OAI21X1 U493 ( .A(n1034), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1607) );
  OAI21X1 U495 ( .A(n1035), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1606) );
  OAI21X1 U497 ( .A(n1036), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1605) );
  OAI21X1 U499 ( .A(n1037), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1604) );
  OAI21X1 U501 ( .A(n1038), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1603) );
  NAND3X1 U503 ( .A(n973), .B(n1829), .C(n1602), .Y(n1611) );
  OAI21X1 U504 ( .A(n1039), .B(n981), .C(n1600), .Y(n1118) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1600) );
  OAI21X1 U506 ( .A(n1040), .B(n980), .C(n1599), .Y(n1117) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1599) );
  OAI21X1 U508 ( .A(n1041), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1598) );
  OAI21X1 U510 ( .A(n1042), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1597) );
  OAI21X1 U512 ( .A(n1043), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1596) );
  OAI21X1 U514 ( .A(n1044), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1595) );
  OAI21X1 U516 ( .A(n1045), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1594) );
  OAI21X1 U518 ( .A(n1046), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1593) );
  NAND3X1 U520 ( .A(n1767), .B(n1829), .C(n1632), .Y(n1601) );
  OAI21X1 U521 ( .A(n1031), .B(n979), .C(n1590), .Y(n1110) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1590) );
  OAI21X1 U523 ( .A(n1032), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1589) );
  OAI21X1 U525 ( .A(n1033), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1588) );
  OAI21X1 U527 ( .A(n1034), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1587) );
  OAI21X1 U529 ( .A(n1035), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1586) );
  OAI21X1 U531 ( .A(n1036), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1585) );
  OAI21X1 U533 ( .A(n1037), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1584) );
  OAI21X1 U535 ( .A(n1038), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1583) );
  NAND3X1 U537 ( .A(n973), .B(n1829), .C(n1582), .Y(n1591) );
  OAI21X1 U538 ( .A(n1039), .B(n978), .C(n1580), .Y(n1102) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1580) );
  OAI21X1 U540 ( .A(n1040), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1579) );
  OAI21X1 U542 ( .A(n1041), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1578) );
  OAI21X1 U544 ( .A(n1042), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1577) );
  OAI21X1 U546 ( .A(n1043), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1576) );
  OAI21X1 U548 ( .A(n1044), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1575) );
  OAI21X1 U550 ( .A(n1045), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1574) );
  OAI21X1 U552 ( .A(n1046), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1573) );
  NAND3X1 U554 ( .A(n969), .B(n1829), .C(n1652), .Y(n1581) );
  OAI21X1 U555 ( .A(n1031), .B(n977), .C(n1571), .Y(n1094) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1571) );
  OAI21X1 U557 ( .A(n1032), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1570) );
  OAI21X1 U559 ( .A(n1033), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1569) );
  OAI21X1 U561 ( .A(n1034), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1568) );
  OAI21X1 U563 ( .A(n1035), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1567) );
  OAI21X1 U565 ( .A(n1036), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1566) );
  OAI21X1 U567 ( .A(n1037), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1565) );
  OAI21X1 U569 ( .A(n1038), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1564) );
  NAND3X1 U571 ( .A(n973), .B(n1829), .C(n1563), .Y(n1572) );
  OAI21X1 U572 ( .A(n1039), .B(n976), .C(n1561), .Y(n1086) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1561) );
  OAI21X1 U574 ( .A(n1040), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1560) );
  OAI21X1 U576 ( .A(n1041), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1559) );
  OAI21X1 U578 ( .A(n1042), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1558) );
  OAI21X1 U580 ( .A(n1043), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1557) );
  OAI21X1 U582 ( .A(n1044), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1556) );
  OAI21X1 U584 ( .A(n1045), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1555) );
  OAI21X1 U586 ( .A(n1046), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1554) );
  NAND3X1 U588 ( .A(n969), .B(n1829), .C(n1632), .Y(n1562) );
  OAI21X1 U590 ( .A(n1031), .B(n975), .C(n1551), .Y(n1078) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1551) );
  OAI21X1 U592 ( .A(n1032), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1550) );
  OAI21X1 U594 ( .A(n1033), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1549) );
  OAI21X1 U596 ( .A(n1034), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1548) );
  OAI21X1 U598 ( .A(n1035), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1547) );
  OAI21X1 U600 ( .A(n1036), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1546) );
  OAI21X1 U602 ( .A(n1037), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1545) );
  OAI21X1 U604 ( .A(n1038), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1544) );
  NAND3X1 U606 ( .A(n973), .B(n1829), .C(n1543), .Y(n1552) );
  OAI21X1 U607 ( .A(n1039), .B(n974), .C(n1541), .Y(n1070) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1541) );
  OAI21X1 U609 ( .A(n1040), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1540) );
  OAI21X1 U611 ( .A(n1041), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1539) );
  OAI21X1 U613 ( .A(n1042), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1538) );
  OAI21X1 U615 ( .A(n1043), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1537) );
  OAI21X1 U617 ( .A(n1044), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1536) );
  OAI21X1 U619 ( .A(n1045), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1535) );
  OAI21X1 U621 ( .A(n1046), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1534) );
  NAND3X1 U623 ( .A(n967), .B(n1829), .C(n1652), .Y(n1542) );
  OAI21X1 U624 ( .A(n1031), .B(n8), .C(n1533), .Y(n1062) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1533) );
  OAI21X1 U626 ( .A(n1032), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1532) );
  OAI21X1 U628 ( .A(n1033), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1531) );
  OAI21X1 U630 ( .A(n1034), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1530) );
  OAI21X1 U632 ( .A(n1035), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1529) );
  OAI21X1 U634 ( .A(n1036), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1528) );
  OAI21X1 U636 ( .A(n1037), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1527) );
  OAI21X1 U638 ( .A(n1038), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1526) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1819) );
  OAI21X1 U642 ( .A(n1039), .B(n972), .C(n1523), .Y(n1054) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1523) );
  OAI21X1 U644 ( .A(n1040), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1522) );
  OAI21X1 U646 ( .A(n1041), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1521) );
  OAI21X1 U648 ( .A(n1042), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1520) );
  OAI21X1 U650 ( .A(n1043), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1519) );
  OAI21X1 U652 ( .A(n1044), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1518) );
  OAI21X1 U654 ( .A(n1045), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1517) );
  OAI21X1 U656 ( .A(n1046), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1516) );
  NAND3X1 U658 ( .A(n967), .B(n1829), .C(n1632), .Y(n1524) );
  NOR3X1 U661 ( .A(n1512), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1513) );
  NOR3X1 U662 ( .A(n1511), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1514) );
  AOI21X1 U663 ( .A(n461), .B(n1510), .C(n963), .Y(n1839) );
  OAI21X1 U665 ( .A(rd), .B(n1509), .C(wr), .Y(n1510) );
  NAND3X1 U667 ( .A(n1508), .B(n1026), .C(n1507), .Y(n1509) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1507) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1508) );
  AOI21X1 U670 ( .A(n448), .B(n1505), .C(n1025), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1504), .C(n4), .Y(n1505) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1787), .C(\mem<0><1> ), .D(n1632), .Y(
        n1502) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1807), .C(\mem<2><1> ), .D(n1652), .Y(
        n1503) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1787), .C(\mem<4><1> ), .D(n1632), .Y(
        n1500) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1807), .C(\mem<6><1> ), .D(n1652), .Y(
        n1501) );
  AOI22X1 U678 ( .A(n1592), .B(n892), .C(n1631), .D(n932), .Y(n1506) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1787), .C(\mem<12><1> ), .D(n1632), .Y(
        n1498) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1807), .C(\mem<14><1> ), .D(n1652), .Y(
        n1499) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1787), .C(\mem<8><1> ), .D(n1632), .Y(
        n1496) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1807), .C(\mem<10><1> ), .D(n1652), .Y(
        n1497) );
  AOI21X1 U685 ( .A(n447), .B(n1494), .C(n1025), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1492), .C(n950), .Y(n1494) );
  AOI21X1 U687 ( .A(n1490), .B(n1489), .C(n971), .Y(n1491) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1787), .C(\mem<0><0> ), .D(n1632), .Y(
        n1489) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1807), .C(\mem<2><0> ), .D(n1652), .Y(
        n1490) );
  AOI21X1 U690 ( .A(n1488), .B(n1487), .C(n970), .Y(n1493) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1787), .C(\mem<4><0> ), .D(n1632), .Y(
        n1487) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1807), .C(\mem<6><0> ), .D(n1652), .Y(
        n1488) );
  AOI22X1 U693 ( .A(n1592), .B(n890), .C(n1631), .D(n930), .Y(n1495) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1787), .C(\mem<12><0> ), .D(n1632), .Y(
        n1485) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1807), .C(\mem<14><0> ), .D(n1652), .Y(
        n1486) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1787), .C(\mem<8><0> ), .D(n1632), .Y(
        n1483) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1807), .C(\mem<10><0> ), .D(n1652), .Y(
        n1484) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1482) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1681), .C(\mem<19><7> ), .D(n1700), .Y(
        n1477) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1719), .C(\mem<23><7> ), .D(n1738), .Y(
        n1478) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1757), .C(\mem<27><7> ), .D(n1777), .Y(
        n1480) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1797), .C(\mem<31><7> ), .D(n1818), .Y(
        n1481) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1525), .C(\mem<3><7> ), .D(n1543), .Y(
        n1472) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1563), .C(\mem<7><7> ), .D(n1582), .Y(
        n1473) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1602), .C(\mem<11><7> ), .D(n1621), .Y(
        n1475) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1642), .C(\mem<15><7> ), .D(n1662), .Y(
        n1476) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1471) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1681), .C(\mem<19><6> ), .D(n1700), .Y(
        n1466) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1719), .C(\mem<23><6> ), .D(n1738), .Y(
        n1467) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1757), .C(\mem<27><6> ), .D(n1777), .Y(
        n1469) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1797), .C(\mem<31><6> ), .D(n1818), .Y(
        n1470) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1525), .C(\mem<3><6> ), .D(n1543), .Y(
        n1461) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1563), .C(\mem<7><6> ), .D(n1582), .Y(
        n1462) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1602), .C(\mem<11><6> ), .D(n1621), .Y(
        n1464) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1642), .C(\mem<15><6> ), .D(n1662), .Y(
        n1465) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1460) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1681), .C(\mem<19><5> ), .D(n1700), .Y(
        n1455) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1719), .C(\mem<23><5> ), .D(n1738), .Y(
        n1456) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1757), .C(\mem<27><5> ), .D(n1777), .Y(
        n1458) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1797), .C(\mem<31><5> ), .D(n1818), .Y(
        n1459) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1525), .C(\mem<3><5> ), .D(n1543), .Y(
        n1450) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1563), .C(\mem<7><5> ), .D(n1582), .Y(
        n1451) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1602), .C(\mem<11><5> ), .D(n1621), .Y(
        n1453) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1642), .C(\mem<15><5> ), .D(n1662), .Y(
        n1454) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1449) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1681), .C(\mem<19><4> ), .D(n1700), .Y(
        n1444) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1719), .C(\mem<23><4> ), .D(n1738), .Y(
        n1445) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1757), .C(\mem<27><4> ), .D(n1777), .Y(
        n1447) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1797), .C(\mem<31><4> ), .D(n1818), .Y(
        n1448) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1525), .C(\mem<3><4> ), .D(n1543), .Y(
        n1439) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1563), .C(\mem<7><4> ), .D(n1582), .Y(
        n1440) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1602), .C(\mem<11><4> ), .D(n1621), .Y(
        n1442) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1642), .C(\mem<15><4> ), .D(n1662), .Y(
        n1443) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1438) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1681), .C(\mem<19><3> ), .D(n1700), .Y(
        n1433) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1719), .C(\mem<23><3> ), .D(n1738), .Y(
        n1434) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1757), .C(\mem<27><3> ), .D(n1777), .Y(
        n1436) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1797), .C(\mem<31><3> ), .D(n1818), .Y(
        n1437) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1525), .C(\mem<3><3> ), .D(n1543), .Y(
        n1428) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1563), .C(\mem<7><3> ), .D(n1582), .Y(
        n1429) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1602), .C(\mem<11><3> ), .D(n1621), .Y(
        n1431) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1642), .C(\mem<15><3> ), .D(n1662), .Y(
        n1432) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1427) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1681), .C(\mem<19><2> ), .D(n1700), .Y(
        n1422) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1719), .C(\mem<23><2> ), .D(n1738), .Y(
        n1423) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1757), .C(\mem<27><2> ), .D(n1777), .Y(
        n1425) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1797), .C(\mem<31><2> ), .D(n1818), .Y(
        n1426) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1525), .C(\mem<3><2> ), .D(n1543), .Y(
        n1417) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1563), .C(\mem<7><2> ), .D(n1582), .Y(
        n1418) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1602), .C(\mem<11><2> ), .D(n1621), .Y(
        n1420) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1642), .C(\mem<15><2> ), .D(n1662), .Y(
        n1421) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1416) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1681), .C(\mem<19><1> ), .D(n1700), .Y(
        n1411) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1719), .C(\mem<23><1> ), .D(n1738), .Y(
        n1412) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1757), .C(\mem<27><1> ), .D(n1777), .Y(
        n1414) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1797), .C(\mem<31><1> ), .D(n1818), .Y(
        n1415) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1525), .C(\mem<3><1> ), .D(n1543), .Y(
        n1406) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1563), .C(\mem<7><1> ), .D(n1582), .Y(
        n1407) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1602), .C(\mem<11><1> ), .D(n1621), .Y(
        n1409) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1642), .C(\mem<15><1> ), .D(n1662), .Y(
        n1410) );
  AOI21X1 U777 ( .A(n435), .B(n1404), .C(n1025), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1402), .C(n949), .Y(n1404) );
  AOI21X1 U779 ( .A(n1400), .B(n1399), .C(n971), .Y(n1401) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1787), .C(\mem<0><7> ), .D(n1632), .Y(
        n1399) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1807), .C(\mem<2><7> ), .D(n1652), .Y(
        n1400) );
  AOI21X1 U782 ( .A(n1398), .B(n1397), .C(n970), .Y(n1403) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1787), .C(\mem<4><7> ), .D(n1632), .Y(
        n1397) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1807), .C(\mem<6><7> ), .D(n1652), .Y(
        n1398) );
  AOI22X1 U785 ( .A(n1592), .B(n888), .C(n1631), .D(n928), .Y(n1405) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1787), .C(\mem<12><7> ), .D(n1632), .Y(
        n1395) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1807), .C(\mem<14><7> ), .D(n1652), .Y(
        n1396) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1787), .C(\mem<8><7> ), .D(n1632), .Y(
        n1393) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1807), .C(\mem<10><7> ), .D(n1652), .Y(
        n1394) );
  AOI21X1 U792 ( .A(n434), .B(n1391), .C(n1025), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1389), .C(n948), .Y(n1391) );
  AOI21X1 U794 ( .A(n1387), .B(n1386), .C(n971), .Y(n1388) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1787), .C(\mem<0><6> ), .D(n1632), .Y(
        n1386) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1807), .C(\mem<2><6> ), .D(n1652), .Y(
        n1387) );
  AOI21X1 U797 ( .A(n1385), .B(n1384), .C(n970), .Y(n1390) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1787), .C(\mem<4><6> ), .D(n1632), .Y(
        n1384) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1807), .C(\mem<6><6> ), .D(n1652), .Y(
        n1385) );
  AOI22X1 U800 ( .A(n1592), .B(n886), .C(n1631), .D(n926), .Y(n1392) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1787), .C(\mem<12><6> ), .D(n1632), .Y(
        n1382) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1807), .C(\mem<14><6> ), .D(n1652), .Y(
        n1383) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1787), .C(\mem<8><6> ), .D(n1632), .Y(
        n1380) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1807), .C(\mem<10><6> ), .D(n1652), .Y(
        n1381) );
  AOI21X1 U807 ( .A(n422), .B(n1378), .C(n1025), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1376), .C(n947), .Y(n1378) );
  AOI21X1 U809 ( .A(n1374), .B(n1373), .C(n971), .Y(n1375) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1787), .C(\mem<0><5> ), .D(n1632), .Y(
        n1373) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1807), .C(\mem<2><5> ), .D(n1652), .Y(
        n1374) );
  AOI21X1 U812 ( .A(n1372), .B(n1371), .C(n970), .Y(n1377) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1787), .C(\mem<4><5> ), .D(n1632), .Y(
        n1371) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1807), .C(\mem<6><5> ), .D(n1652), .Y(
        n1372) );
  AOI22X1 U815 ( .A(n1592), .B(n884), .C(n1631), .D(n924), .Y(n1379) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1787), .C(\mem<12><5> ), .D(n1632), .Y(
        n1369) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1807), .C(\mem<14><5> ), .D(n1652), .Y(
        n1370) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1787), .C(\mem<8><5> ), .D(n1632), .Y(
        n1367) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1807), .C(\mem<10><5> ), .D(n1652), .Y(
        n1368) );
  AOI21X1 U822 ( .A(n421), .B(n1365), .C(n1025), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1363), .C(n946), .Y(n1365) );
  AOI21X1 U824 ( .A(n1361), .B(n1360), .C(n971), .Y(n1362) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1787), .C(\mem<0><4> ), .D(n1632), .Y(
        n1360) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1807), .C(\mem<2><4> ), .D(n1652), .Y(
        n1361) );
  AOI21X1 U827 ( .A(n1359), .B(n1358), .C(n970), .Y(n1364) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1787), .C(\mem<4><4> ), .D(n1632), .Y(
        n1358) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1807), .C(\mem<6><4> ), .D(n1652), .Y(
        n1359) );
  AOI22X1 U830 ( .A(n1592), .B(n882), .C(n1631), .D(n922), .Y(n1366) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1787), .C(\mem<12><4> ), .D(n1632), .Y(
        n1356) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1807), .C(\mem<14><4> ), .D(n1652), .Y(
        n1357) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1787), .C(\mem<8><4> ), .D(n1632), .Y(
        n1354) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1807), .C(\mem<10><4> ), .D(n1652), .Y(
        n1355) );
  AOI21X1 U837 ( .A(n409), .B(n1352), .C(n1025), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1350), .C(n945), .Y(n1352) );
  AOI21X1 U839 ( .A(n1348), .B(n1347), .C(n971), .Y(n1349) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1787), .C(\mem<0><3> ), .D(n1632), .Y(
        n1347) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1807), .C(\mem<2><3> ), .D(n1652), .Y(
        n1348) );
  AOI21X1 U842 ( .A(n1346), .B(n1345), .C(n970), .Y(n1351) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1787), .C(\mem<4><3> ), .D(n1632), .Y(
        n1345) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1807), .C(\mem<6><3> ), .D(n1652), .Y(
        n1346) );
  AOI22X1 U845 ( .A(n1592), .B(n880), .C(n1631), .D(n920), .Y(n1353) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1787), .C(\mem<12><3> ), .D(n1632), .Y(
        n1343) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1807), .C(\mem<14><3> ), .D(n1652), .Y(
        n1344) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1787), .C(\mem<8><3> ), .D(n1632), .Y(
        n1341) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1807), .C(\mem<10><3> ), .D(n1652), .Y(
        n1342) );
  AOI21X1 U852 ( .A(n408), .B(n1339), .C(n1025), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1337), .C(n944), .Y(n1339) );
  AOI21X1 U854 ( .A(n1335), .B(n1334), .C(n971), .Y(n1336) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1787), .C(\mem<0><2> ), .D(n1632), .Y(
        n1334) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1807), .C(\mem<2><2> ), .D(n1652), .Y(
        n1335) );
  AOI21X1 U857 ( .A(n1333), .B(n1332), .C(n970), .Y(n1338) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1787), .C(\mem<4><2> ), .D(n1632), .Y(
        n1332) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1807), .C(\mem<6><2> ), .D(n1652), .Y(
        n1333) );
  AOI22X1 U860 ( .A(n1592), .B(n878), .C(n1631), .D(n918), .Y(n1340) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1787), .C(\mem<12><2> ), .D(n1632), .Y(
        n1330) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1807), .C(\mem<14><2> ), .D(n1652), .Y(
        n1331) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1787), .C(\mem<8><2> ), .D(n1632), .Y(
        n1328) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1807), .C(\mem<10><2> ), .D(n1652), .Y(
        n1329) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1327) );
  NOR2X1 U868 ( .A(n1030), .B(\addr_1c<4> ), .Y(n1326) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1325) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1681), .C(\mem<19><0> ), .D(n1700), .Y(
        n1320) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1719), .C(\mem<23><0> ), .D(n1738), .Y(
        n1321) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1757), .C(\mem<27><0> ), .D(n1777), .Y(
        n1323) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1797), .C(\mem<31><0> ), .D(n1818), .Y(
        n1324) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1525), .C(\mem<3><0> ), .D(n1543), .Y(
        n1313) );
  NAND2X1 U877 ( .A(n1028), .B(n1029), .Y(n1515) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1563), .C(\mem<7><0> ), .D(n1582), .Y(
        n1314) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1029), .Y(n1553) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1602), .C(\mem<11><0> ), .D(n1621), .Y(
        n1316) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1642), .C(\mem<15><0> ), .D(n1662), .Y(
        n1317) );
  dff_152 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_151 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1013) );
  dff_150 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1013)
         );
  dff_149 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1013)
         );
  dff_148 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1013)
         );
  dff_147 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1013)
         );
  dff_146 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1013)
         );
  dff_145 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1013)
         );
  dff_144 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1013)
         );
  dff_143 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1013)
         );
  dff_142 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_141 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_140 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1012) );
  dff_139 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1012) );
  dff_138 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1012) );
  dff_137 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_136 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_135 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_134 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_133 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_132 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_131 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_130 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_129 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_128 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_127 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_126 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_125 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_124 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_123 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_122 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_121 \reg2[0]  ( .q(\data_out<0> ), .d(n1022), .clk(clk), .rst(n1013) );
  dff_120 \reg2[1]  ( .q(\data_out<1> ), .d(n1021), .clk(clk), .rst(n1013) );
  dff_119 \reg2[2]  ( .q(\data_out<2> ), .d(n1020), .clk(clk), .rst(n1013) );
  dff_118 \reg2[3]  ( .q(\data_out<3> ), .d(n1019), .clk(clk), .rst(n1013) );
  dff_117 \reg2[4]  ( .q(\data_out<4> ), .d(n1018), .clk(clk), .rst(n1013) );
  dff_116 \reg2[5]  ( .q(\data_out<5> ), .d(n1017), .clk(clk), .rst(n1013) );
  dff_115 \reg2[6]  ( .q(\data_out<6> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_114 \reg2[7]  ( .q(\data_out<7> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_113 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1012) );
  dff_112 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1012) );
  dff_111 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_110 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_109 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_108 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1013) );
  dff_107 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_106 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_105 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_104 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_103 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_102 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1013) );
  OR2X1 U2 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1511) );
  AND2X1 U3 ( .A(\addr_1c<4> ), .B(n1525), .Y(n1828) );
  INVX1 U4 ( .A(rst), .Y(n1014) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1030) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1029) );
  INVX1 U7 ( .A(wr1), .Y(n1026) );
  OR2X1 U8 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1512) );
  INVX1 U23 ( .A(\addr_1c<0> ), .Y(n1027) );
  AND2X1 U24 ( .A(n1027), .B(n1030), .Y(n1311) );
  AND2X1 U25 ( .A(\addr_1c<0> ), .B(n1030), .Y(n1312) );
  AND2X1 U26 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1319) );
  AND2X1 U27 ( .A(\addr_1c<3> ), .B(n1027), .Y(n1318) );
  INVX1 U28 ( .A(\addr_1c<1> ), .Y(n1028) );
  AND2X1 U29 ( .A(n1592), .B(n1319), .Y(n1777) );
  AND2X1 U35 ( .A(n1592), .B(n1318), .Y(n1757) );
  AND2X1 U36 ( .A(n940), .B(n1319), .Y(n1738) );
  AND2X1 U37 ( .A(n940), .B(n1318), .Y(n1719) );
  AND2X1 U38 ( .A(n1319), .B(n951), .Y(n1700) );
  AND2X1 U39 ( .A(n1318), .B(n951), .Y(n1681) );
  AND2X1 U40 ( .A(n1312), .B(n1592), .Y(n1621) );
  AND2X1 U41 ( .A(n1592), .B(n1311), .Y(n1602) );
  AND2X1 U42 ( .A(n1312), .B(n940), .Y(n1582) );
  AND2X1 U43 ( .A(n940), .B(n1311), .Y(n1563) );
  OR2X1 U44 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U46 ( .A(n1312), .B(n951), .Y(n1543) );
  OR2X1 U47 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U48 ( .A(n1631), .B(n1311), .Y(n1642) );
  AND2X1 U49 ( .A(n1312), .B(n1631), .Y(n1662) );
  AND2X1 U50 ( .A(n1318), .B(n1631), .Y(n1797) );
  AND2X1 U51 ( .A(\addr_1c<2> ), .B(n1028), .Y(n1592) );
  AND2X1 U52 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1631) );
  BUFX2 U53 ( .A(n961), .Y(n1010) );
  BUFX2 U54 ( .A(n961), .Y(n1009) );
  BUFX2 U55 ( .A(n960), .Y(n1007) );
  BUFX2 U56 ( .A(n960), .Y(n1006) );
  BUFX2 U57 ( .A(n959), .Y(n1004) );
  BUFX2 U58 ( .A(n959), .Y(n1003) );
  BUFX2 U59 ( .A(n958), .Y(n1001) );
  BUFX2 U60 ( .A(n958), .Y(n1000) );
  BUFX2 U61 ( .A(n957), .Y(n990) );
  BUFX2 U62 ( .A(n957), .Y(n989) );
  BUFX2 U63 ( .A(n956), .Y(n987) );
  BUFX2 U64 ( .A(n956), .Y(n986) );
  BUFX2 U65 ( .A(n955), .Y(n984) );
  BUFX2 U66 ( .A(n955), .Y(n983) );
  BUFX2 U67 ( .A(n954), .Y(n981) );
  BUFX2 U68 ( .A(n954), .Y(n980) );
  INVX1 U69 ( .A(\data_in_1c<0> ), .Y(n1031) );
  INVX1 U70 ( .A(\data_in_1c<1> ), .Y(n1032) );
  INVX1 U71 ( .A(\data_in_1c<2> ), .Y(n1033) );
  INVX1 U72 ( .A(\data_in_1c<3> ), .Y(n1034) );
  INVX1 U73 ( .A(\data_in_1c<4> ), .Y(n1035) );
  INVX1 U74 ( .A(\data_in_1c<5> ), .Y(n1036) );
  INVX1 U75 ( .A(\data_in_1c<6> ), .Y(n1037) );
  INVX1 U76 ( .A(\data_in_1c<7> ), .Y(n1038) );
  INVX1 U77 ( .A(\data_in_1c<8> ), .Y(n1039) );
  INVX1 U78 ( .A(\data_in_1c<9> ), .Y(n1040) );
  INVX1 U79 ( .A(\data_in_1c<10> ), .Y(n1041) );
  INVX1 U80 ( .A(\data_in_1c<11> ), .Y(n1042) );
  INVX1 U81 ( .A(\data_in_1c<12> ), .Y(n1043) );
  INVX1 U82 ( .A(\data_in_1c<13> ), .Y(n1044) );
  INVX1 U83 ( .A(\data_in_1c<14> ), .Y(n1045) );
  INVX1 U84 ( .A(\data_in_1c<15> ), .Y(n1046) );
  AND2X1 U85 ( .A(n1828), .B(\mem<32><0> ), .Y(n1492) );
  AND2X1 U86 ( .A(n1828), .B(\mem<32><1> ), .Y(n1504) );
  AND2X1 U87 ( .A(n1828), .B(\mem<32><2> ), .Y(n1337) );
  AND2X1 U88 ( .A(n1828), .B(\mem<32><3> ), .Y(n1350) );
  AND2X1 U89 ( .A(n1828), .B(\mem<32><4> ), .Y(n1363) );
  AND2X1 U90 ( .A(n1828), .B(\mem<32><5> ), .Y(n1376) );
  AND2X1 U91 ( .A(n1828), .B(\mem<32><6> ), .Y(n1389) );
  AND2X1 U92 ( .A(n1828), .B(\mem<32><7> ), .Y(n1402) );
  INVX1 U93 ( .A(rd1), .Y(n1025) );
  INVX1 U129 ( .A(n1325), .Y(n1022) );
  INVX1 U589 ( .A(n1416), .Y(n1021) );
  INVX1 U640 ( .A(n1427), .Y(n1020) );
  INVX1 U659 ( .A(n1438), .Y(n1019) );
  INVX1 U660 ( .A(n1449), .Y(n1018) );
  INVX1 U664 ( .A(n1460), .Y(n1017) );
  INVX1 U666 ( .A(n1471), .Y(n1016) );
  INVX1 U672 ( .A(n1482), .Y(n1015) );
  INVX2 U675 ( .A(n1014), .Y(n1012) );
  AND2X1 U679 ( .A(wr1), .B(n1014), .Y(n1829) );
  AND2X1 U682 ( .A(n1631), .B(n964), .Y(n1808) );
  AND2X1 U694 ( .A(n1592), .B(n964), .Y(n1767) );
  AND2X1 U697 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U701 ( .A(n1), .Y(n2) );
  AND2X1 U706 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U712 ( .A(n3), .Y(n4) );
  AND2X1 U717 ( .A(n1818), .B(n189), .Y(n5) );
  INVX1 U723 ( .A(n5), .Y(n6) );
  AND2X1 U728 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U734 ( .A(n7), .Y(n8) );
  OR2X1 U739 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U745 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U750 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U756 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U761 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U767 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U772 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U786 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U789 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U801 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U804 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U816 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U819 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U831 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U834 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U846 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U849 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U861 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U864 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U870 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U875 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U882 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U883 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U884 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U885 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U886 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U887 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U888 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U889 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U890 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U891 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U892 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U893 ( .A(n973), .B(n1829), .Y(n189) );
  AND2X1 U894 ( .A(n1829), .B(n1525), .Y(n289) );
  INVX1 U895 ( .A(n1014), .Y(n1013) );
  AND2X1 U896 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U897 ( .A(n348), .Y(n372) );
  AND2X1 U898 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U899 ( .A(n379), .Y(n381) );
  AND2X1 U900 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U901 ( .A(n386), .Y(n387) );
  AND2X1 U902 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U903 ( .A(n401), .Y(n402) );
  BUFX2 U904 ( .A(n1340), .Y(n408) );
  BUFX2 U905 ( .A(n1353), .Y(n409) );
  BUFX2 U906 ( .A(n1366), .Y(n421) );
  BUFX2 U907 ( .A(n1379), .Y(n422) );
  BUFX2 U908 ( .A(n1392), .Y(n434) );
  BUFX2 U909 ( .A(n1405), .Y(n435) );
  BUFX2 U910 ( .A(n1495), .Y(n447) );
  BUFX2 U911 ( .A(n1506), .Y(n448) );
  AND2X2 U912 ( .A(rd), .B(n1509), .Y(n460) );
  INVX1 U913 ( .A(n460), .Y(n461) );
  INVX1 U914 ( .A(n1315), .Y(n473) );
  INVX1 U915 ( .A(n1316), .Y(n474) );
  INVX1 U916 ( .A(n1317), .Y(n486) );
  INVX1 U917 ( .A(n1408), .Y(n487) );
  INVX1 U918 ( .A(n1409), .Y(n507) );
  INVX1 U919 ( .A(n1410), .Y(n508) );
  INVX1 U920 ( .A(n1419), .Y(n522) );
  INVX1 U921 ( .A(n1420), .Y(n523) );
  INVX1 U922 ( .A(n1421), .Y(n537) );
  INVX1 U923 ( .A(n1430), .Y(n538) );
  INVX1 U924 ( .A(n1431), .Y(n552) );
  INVX1 U925 ( .A(n1432), .Y(n553) );
  INVX1 U926 ( .A(n1441), .Y(n567) );
  INVX1 U927 ( .A(n1442), .Y(n568) );
  INVX1 U928 ( .A(n1443), .Y(n582) );
  INVX1 U929 ( .A(n1452), .Y(n583) );
  INVX1 U930 ( .A(n1453), .Y(n591) );
  INVX1 U931 ( .A(n1454), .Y(n592) );
  INVX1 U932 ( .A(n1463), .Y(n871) );
  INVX1 U933 ( .A(n1464), .Y(n872) );
  INVX1 U934 ( .A(n1465), .Y(n873) );
  INVX1 U935 ( .A(n1474), .Y(n874) );
  INVX1 U936 ( .A(n1475), .Y(n875) );
  INVX1 U937 ( .A(n1476), .Y(n876) );
  AND2X2 U938 ( .A(n1329), .B(n1328), .Y(n877) );
  INVX1 U939 ( .A(n877), .Y(n878) );
  AND2X2 U940 ( .A(n1342), .B(n1341), .Y(n879) );
  INVX1 U941 ( .A(n879), .Y(n880) );
  AND2X2 U942 ( .A(n1355), .B(n1354), .Y(n881) );
  INVX1 U943 ( .A(n881), .Y(n882) );
  AND2X2 U944 ( .A(n1368), .B(n1367), .Y(n883) );
  INVX1 U945 ( .A(n883), .Y(n884) );
  AND2X2 U946 ( .A(n1381), .B(n1380), .Y(n885) );
  INVX1 U947 ( .A(n885), .Y(n886) );
  AND2X2 U948 ( .A(n1394), .B(n1393), .Y(n887) );
  INVX1 U949 ( .A(n887), .Y(n888) );
  AND2X2 U950 ( .A(n1484), .B(n1483), .Y(n889) );
  INVX1 U951 ( .A(n889), .Y(n890) );
  AND2X2 U952 ( .A(n1497), .B(n1496), .Y(n891) );
  INVX1 U953 ( .A(n891), .Y(n892) );
  INVX1 U954 ( .A(n1322), .Y(n893) );
  INVX1 U955 ( .A(n1323), .Y(n894) );
  INVX1 U956 ( .A(n1324), .Y(n895) );
  INVX1 U957 ( .A(n1413), .Y(n896) );
  INVX1 U958 ( .A(n1414), .Y(n897) );
  INVX1 U959 ( .A(n1415), .Y(n898) );
  INVX1 U960 ( .A(n1424), .Y(n899) );
  INVX1 U961 ( .A(n1425), .Y(n900) );
  INVX1 U962 ( .A(n1426), .Y(n901) );
  INVX1 U963 ( .A(n1435), .Y(n902) );
  INVX1 U964 ( .A(n1436), .Y(n903) );
  INVX1 U965 ( .A(n1437), .Y(n904) );
  INVX1 U966 ( .A(n1446), .Y(n905) );
  INVX1 U967 ( .A(n1447), .Y(n906) );
  INVX1 U968 ( .A(n1448), .Y(n907) );
  INVX1 U969 ( .A(n1457), .Y(n908) );
  INVX1 U970 ( .A(n1458), .Y(n909) );
  INVX1 U971 ( .A(n1459), .Y(n910) );
  INVX1 U972 ( .A(n1468), .Y(n911) );
  INVX1 U973 ( .A(n1469), .Y(n912) );
  INVX1 U974 ( .A(n1470), .Y(n913) );
  INVX1 U975 ( .A(n1479), .Y(n914) );
  INVX1 U976 ( .A(n1480), .Y(n915) );
  INVX1 U977 ( .A(n1481), .Y(n916) );
  AND2X2 U978 ( .A(n1331), .B(n1330), .Y(n917) );
  INVX1 U979 ( .A(n917), .Y(n918) );
  AND2X2 U980 ( .A(n1344), .B(n1343), .Y(n919) );
  INVX1 U981 ( .A(n919), .Y(n920) );
  AND2X2 U982 ( .A(n1357), .B(n1356), .Y(n921) );
  INVX1 U983 ( .A(n921), .Y(n922) );
  AND2X2 U984 ( .A(n1370), .B(n1369), .Y(n923) );
  INVX1 U985 ( .A(n923), .Y(n924) );
  AND2X2 U986 ( .A(n1383), .B(n1382), .Y(n925) );
  INVX1 U987 ( .A(n925), .Y(n926) );
  AND2X2 U988 ( .A(n1396), .B(n1395), .Y(n927) );
  INVX1 U989 ( .A(n927), .Y(n928) );
  AND2X2 U990 ( .A(n1486), .B(n1485), .Y(n929) );
  INVX1 U991 ( .A(n929), .Y(n930) );
  AND2X2 U992 ( .A(n1499), .B(n1498), .Y(n931) );
  INVX1 U993 ( .A(n931), .Y(n932) );
  BUFX2 U994 ( .A(n1338), .Y(n933) );
  BUFX2 U995 ( .A(n1351), .Y(n934) );
  BUFX2 U996 ( .A(n1364), .Y(n935) );
  BUFX2 U997 ( .A(n1377), .Y(n936) );
  BUFX2 U998 ( .A(n1390), .Y(n937) );
  BUFX2 U999 ( .A(n1403), .Y(n938) );
  BUFX2 U1000 ( .A(n1493), .Y(n939) );
  INVX1 U1001 ( .A(n970), .Y(n940) );
  INVX1 U1002 ( .A(n1500), .Y(n941) );
  INVX1 U1003 ( .A(n1501), .Y(n942) );
  BUFX2 U1004 ( .A(n1553), .Y(n970) );
  BUFX2 U1005 ( .A(n1839), .Y(err) );
  BUFX2 U1006 ( .A(n1336), .Y(n944) );
  BUFX2 U1007 ( .A(n1349), .Y(n945) );
  BUFX2 U1008 ( .A(n1362), .Y(n946) );
  BUFX2 U1009 ( .A(n1375), .Y(n947) );
  BUFX2 U1010 ( .A(n1388), .Y(n948) );
  BUFX2 U1011 ( .A(n1401), .Y(n949) );
  BUFX2 U1012 ( .A(n1491), .Y(n950) );
  INVX1 U1013 ( .A(n971), .Y(n951) );
  INVX1 U1014 ( .A(n1502), .Y(n952) );
  INVX1 U1015 ( .A(n1503), .Y(n953) );
  BUFX2 U1016 ( .A(n1515), .Y(n971) );
  BUFX2 U1017 ( .A(n1524), .Y(n972) );
  BUFX2 U1018 ( .A(n1542), .Y(n974) );
  BUFX2 U1019 ( .A(n1552), .Y(n975) );
  BUFX2 U1020 ( .A(n1562), .Y(n976) );
  BUFX2 U1021 ( .A(n1572), .Y(n977) );
  BUFX2 U1022 ( .A(n1581), .Y(n978) );
  BUFX2 U1023 ( .A(n1591), .Y(n979) );
  BUFX2 U1024 ( .A(n1611), .Y(n982) );
  BUFX2 U1025 ( .A(n1630), .Y(n985) );
  BUFX2 U1026 ( .A(n1651), .Y(n988) );
  BUFX2 U1027 ( .A(n1671), .Y(n991) );
  BUFX2 U1028 ( .A(n1680), .Y(n992) );
  BUFX2 U1029 ( .A(n1690), .Y(n993) );
  BUFX2 U1030 ( .A(n1699), .Y(n994) );
  BUFX2 U1031 ( .A(n1709), .Y(n995) );
  BUFX2 U1032 ( .A(n1718), .Y(n996) );
  BUFX2 U1033 ( .A(n1728), .Y(n997) );
  BUFX2 U1034 ( .A(n1737), .Y(n998) );
  BUFX2 U1035 ( .A(n1747), .Y(n999) );
  BUFX2 U1036 ( .A(n1766), .Y(n1002) );
  BUFX2 U1037 ( .A(n1786), .Y(n1005) );
  BUFX2 U1038 ( .A(n1806), .Y(n1008) );
  BUFX2 U1039 ( .A(n1819), .Y(n973) );
  AND2X1 U1040 ( .A(n1631), .B(n1319), .Y(n1818) );
  BUFX2 U1041 ( .A(n1838), .Y(n1011) );
  BUFX2 U1042 ( .A(n1601), .Y(n954) );
  BUFX2 U1043 ( .A(n1620), .Y(n955) );
  BUFX2 U1044 ( .A(n1641), .Y(n956) );
  BUFX2 U1045 ( .A(n1661), .Y(n957) );
  BUFX2 U1046 ( .A(n1756), .Y(n958) );
  BUFX2 U1047 ( .A(n1776), .Y(n959) );
  BUFX2 U1048 ( .A(n1796), .Y(n960) );
  BUFX2 U1049 ( .A(n1817), .Y(n961) );
  AND2X1 U1050 ( .A(enable), .B(n1014), .Y(n962) );
  INVX1 U1051 ( .A(n962), .Y(n963) );
  AND2X1 U1052 ( .A(n1514), .B(n1513), .Y(n964) );
  INVX1 U1053 ( .A(n964), .Y(n965) );
  INVX1 U1054 ( .A(n966), .Y(n967) );
  INVX1 U1055 ( .A(n968), .Y(n969) );
  AND2X1 U1056 ( .A(n951), .B(n1311), .Y(n1525) );
  INVX1 U1057 ( .A(rd), .Y(n1023) );
  INVX1 U1058 ( .A(wr), .Y(n1024) );
endmodule


module final_memory_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1842, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1050), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1051), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1052), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1053), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1054), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1055), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1056), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1057), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1058), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1059), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1060), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1061), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1062), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1063), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1064), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1065), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1066), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1067), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1068), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1069), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1070), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1071), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1072), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1073), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1074), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1075), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1076), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1077), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1078), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1079), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1080), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1081), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1082), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1083), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1084), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1085), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1087), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1088), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1089), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1090), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1091), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1092), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1093), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1094), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1095), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1096), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1097), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1098), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1099), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1100), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1101), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1102), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1103), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1104), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1105), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1106), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1107), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1108), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1109), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1110), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1111), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1112), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1113), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1114), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1115), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1116), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1117), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1118), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1119), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1120), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1121), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1122), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1123), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1124), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1125), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1126), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1127), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1128), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1129), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1130), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1131), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1132), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1133), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1134), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1135), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1136), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1137), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1138), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1139), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1140), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1141), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1142), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1143), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1144), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1145), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1146), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1147), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1148), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1149), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1150), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1151), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1152), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1153), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1154), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1155), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1156), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1157), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1158), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1159), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1160), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1161), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1162), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1163), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1164), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1165), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1166), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1167), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1168), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1169), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1170), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1171), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1172), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1173), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1174), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1175), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1176), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1177), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1178), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1179), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1180), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1181), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1182), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1183), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1184), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1185), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1186), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1187), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1188), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1189), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1190), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1191), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1192), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1193), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1194), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1195), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1196), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1197), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1198), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1199), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1200), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1201), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1202), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1203), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1204), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1205), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1206), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1207), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1208), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1209), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1210), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1211), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1212), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1213), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1214), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1215), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1216), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1217), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1218), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1219), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1220), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1221), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1222), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1223), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1224), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1225), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1226), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1227), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1228), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1229), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1230), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1231), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1232), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1233), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1234), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1235), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1236), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1237), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1238), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1239), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1240), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1241), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1242), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1243), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1244), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1245), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1246), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1247), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1248), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1249), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1250), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1251), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1252), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1253), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1254), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1255), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1256), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1257), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1258), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1259), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1260), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1261), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1262), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1263), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1264), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1265), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1266), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1267), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1268), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1269), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1270), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1271), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1272), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1273), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1274), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1275), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1276), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1277), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1278), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1279), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1280), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1281), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1282), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1283), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1284), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1285), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1286), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1287), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1288), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1289), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1290), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1291), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1292), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1293), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1294), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1296), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1297), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1298), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1299), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1300), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1301), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1302), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1303), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1304), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1305), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1306), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1307), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1308), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1309), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1310), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1311), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1312), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1313), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1481), .B(n1480), .Y(n1482) );
  AND2X2 U10 ( .A(n1476), .B(n1475), .Y(n1477) );
  AND2X2 U11 ( .A(n1470), .B(n1469), .Y(n1471) );
  AND2X2 U12 ( .A(n1465), .B(n1464), .Y(n1466) );
  AND2X2 U13 ( .A(n1459), .B(n1458), .Y(n1460) );
  AND2X2 U14 ( .A(n1454), .B(n1453), .Y(n1455) );
  AND2X2 U15 ( .A(n1448), .B(n1447), .Y(n1449) );
  AND2X2 U16 ( .A(n1443), .B(n1442), .Y(n1444) );
  AND2X2 U17 ( .A(n1437), .B(n1436), .Y(n1438) );
  AND2X2 U18 ( .A(n1432), .B(n1431), .Y(n1433) );
  AND2X2 U19 ( .A(n1426), .B(n1425), .Y(n1427) );
  AND2X2 U20 ( .A(n1421), .B(n1420), .Y(n1422) );
  AND2X2 U21 ( .A(n1415), .B(n1414), .Y(n1416) );
  AND2X2 U22 ( .A(n1410), .B(n1409), .Y(n1411) );
  AND2X2 U30 ( .A(n1330), .B(n1030), .Y(n1635) );
  AND2X2 U31 ( .A(n1329), .B(n1030), .Y(n1790) );
  AND2X2 U32 ( .A(n1330), .B(\addr_1c<0> ), .Y(n1655) );
  AND2X2 U33 ( .A(n1329), .B(\addr_1c<0> ), .Y(n1810) );
  AND2X2 U34 ( .A(n1324), .B(n1323), .Y(n1325) );
  AND2X2 U45 ( .A(n1317), .B(n1316), .Y(n1318) );
  NOR3X1 U94 ( .A(n1027), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1026), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1042), .C(n1840), .Y(n1313) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1840) );
  OAI21X1 U98 ( .A(n1011), .B(n1043), .C(n1839), .Y(n1312) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1839) );
  OAI21X1 U100 ( .A(n1011), .B(n1044), .C(n1838), .Y(n1311) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1838) );
  OAI21X1 U102 ( .A(n1011), .B(n1045), .C(n1837), .Y(n1310) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1837) );
  OAI21X1 U104 ( .A(n1011), .B(n1046), .C(n1836), .Y(n1309) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1836) );
  OAI21X1 U106 ( .A(n1011), .B(n1047), .C(n1835), .Y(n1308) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1835) );
  OAI21X1 U108 ( .A(n1011), .B(n1048), .C(n1834), .Y(n1307) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1834) );
  OAI21X1 U110 ( .A(n1011), .B(n1049), .C(n1833), .Y(n1306) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1833) );
  NAND3X1 U112 ( .A(n1832), .B(n1831), .C(n964), .Y(n1841) );
  OAI21X1 U113 ( .A(n6), .B(n1034), .C(n1830), .Y(n1305) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1830) );
  OAI21X1 U115 ( .A(n6), .B(n1035), .C(n1829), .Y(n1304) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1829) );
  OAI21X1 U117 ( .A(n6), .B(n1036), .C(n1828), .Y(n1303) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1828) );
  OAI21X1 U119 ( .A(n6), .B(n1037), .C(n1827), .Y(n1302) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1827) );
  OAI21X1 U121 ( .A(n6), .B(n1038), .C(n1826), .Y(n1301) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1826) );
  OAI21X1 U123 ( .A(n6), .B(n1039), .C(n1825), .Y(n1300) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1825) );
  OAI21X1 U125 ( .A(n6), .B(n1040), .C(n1824), .Y(n1299) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1824) );
  OAI21X1 U127 ( .A(n6), .B(n1041), .C(n1823), .Y(n1298) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1823) );
  OAI21X1 U130 ( .A(n1042), .B(n1010), .C(n1819), .Y(n1297) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1819) );
  OAI21X1 U132 ( .A(n1043), .B(n1009), .C(n1818), .Y(n1296) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1818) );
  OAI21X1 U134 ( .A(n1044), .B(n1009), .C(n1817), .Y(n1295) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1817) );
  OAI21X1 U136 ( .A(n1045), .B(n1009), .C(n1816), .Y(n1294) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1816) );
  OAI21X1 U138 ( .A(n1046), .B(n1009), .C(n1815), .Y(n1293) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1815) );
  OAI21X1 U140 ( .A(n1047), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1814) );
  OAI21X1 U142 ( .A(n1048), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1813) );
  OAI21X1 U144 ( .A(n1049), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1812) );
  NAND3X1 U146 ( .A(n1811), .B(n1832), .C(n1810), .Y(n1820) );
  OAI21X1 U147 ( .A(n1034), .B(n1008), .C(n1808), .Y(n1289) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1808) );
  OAI21X1 U149 ( .A(n1035), .B(n1008), .C(n1807), .Y(n1288) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1807) );
  OAI21X1 U151 ( .A(n1036), .B(n1008), .C(n1806), .Y(n1287) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1806) );
  OAI21X1 U153 ( .A(n1037), .B(n1008), .C(n1805), .Y(n1286) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1805) );
  OAI21X1 U155 ( .A(n1038), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1804) );
  OAI21X1 U157 ( .A(n1039), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1803) );
  OAI21X1 U159 ( .A(n1040), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1802) );
  OAI21X1 U161 ( .A(n1041), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1801) );
  NAND3X1 U163 ( .A(n973), .B(n1832), .C(n1800), .Y(n1809) );
  OAI21X1 U164 ( .A(n1042), .B(n1007), .C(n1798), .Y(n1281) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1798) );
  OAI21X1 U166 ( .A(n1043), .B(n1006), .C(n1797), .Y(n1280) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1797) );
  OAI21X1 U168 ( .A(n1044), .B(n1006), .C(n1796), .Y(n1279) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1796) );
  OAI21X1 U170 ( .A(n1045), .B(n1006), .C(n1795), .Y(n1278) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1795) );
  OAI21X1 U172 ( .A(n1046), .B(n1006), .C(n1794), .Y(n1277) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1794) );
  OAI21X1 U174 ( .A(n1047), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1793) );
  OAI21X1 U176 ( .A(n1048), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1792) );
  OAI21X1 U178 ( .A(n1049), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1791) );
  NAND3X1 U180 ( .A(n1811), .B(n1832), .C(n1790), .Y(n1799) );
  OAI21X1 U181 ( .A(n1034), .B(n1005), .C(n1788), .Y(n1273) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1788) );
  OAI21X1 U183 ( .A(n1035), .B(n1005), .C(n1787), .Y(n1272) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1787) );
  OAI21X1 U185 ( .A(n1036), .B(n1005), .C(n1786), .Y(n1271) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1786) );
  OAI21X1 U187 ( .A(n1037), .B(n1005), .C(n1785), .Y(n1270) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1785) );
  OAI21X1 U189 ( .A(n1038), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1784) );
  OAI21X1 U191 ( .A(n1039), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1783) );
  OAI21X1 U193 ( .A(n1040), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1782) );
  OAI21X1 U195 ( .A(n1041), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1781) );
  NAND3X1 U197 ( .A(n973), .B(n1832), .C(n1780), .Y(n1789) );
  OAI21X1 U198 ( .A(n1042), .B(n1004), .C(n1778), .Y(n1265) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1778) );
  OAI21X1 U200 ( .A(n1043), .B(n1003), .C(n1777), .Y(n1264) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1777) );
  OAI21X1 U202 ( .A(n1044), .B(n1003), .C(n1776), .Y(n1263) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1776) );
  OAI21X1 U204 ( .A(n1045), .B(n1003), .C(n1775), .Y(n1262) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1775) );
  OAI21X1 U206 ( .A(n1046), .B(n1003), .C(n1774), .Y(n1261) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1774) );
  OAI21X1 U208 ( .A(n1047), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1773) );
  OAI21X1 U210 ( .A(n1048), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1772) );
  OAI21X1 U212 ( .A(n1049), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1771) );
  NAND3X1 U214 ( .A(n1810), .B(n1013), .C(n1770), .Y(n1779) );
  OAI21X1 U215 ( .A(n1034), .B(n1002), .C(n1768), .Y(n1257) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1768) );
  OAI21X1 U217 ( .A(n1035), .B(n1002), .C(n1767), .Y(n1256) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1767) );
  OAI21X1 U219 ( .A(n1036), .B(n1002), .C(n1766), .Y(n1255) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1766) );
  OAI21X1 U221 ( .A(n1037), .B(n1002), .C(n1765), .Y(n1254) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1765) );
  OAI21X1 U223 ( .A(n1038), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1764) );
  OAI21X1 U225 ( .A(n1039), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1763) );
  OAI21X1 U227 ( .A(n1040), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1762) );
  OAI21X1 U229 ( .A(n1041), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1761) );
  NAND3X1 U231 ( .A(n973), .B(n1013), .C(n1760), .Y(n1769) );
  OAI21X1 U232 ( .A(n1042), .B(n1001), .C(n1758), .Y(n1249) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1758) );
  OAI21X1 U234 ( .A(n1043), .B(n1000), .C(n1757), .Y(n1248) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1757) );
  OAI21X1 U236 ( .A(n1044), .B(n1000), .C(n1756), .Y(n1247) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1756) );
  OAI21X1 U238 ( .A(n1045), .B(n1000), .C(n1755), .Y(n1246) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1755) );
  OAI21X1 U240 ( .A(n1046), .B(n1000), .C(n1754), .Y(n1245) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1754) );
  OAI21X1 U242 ( .A(n1047), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1753) );
  OAI21X1 U244 ( .A(n1048), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1752) );
  OAI21X1 U246 ( .A(n1049), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1751) );
  NAND3X1 U248 ( .A(n1790), .B(n1013), .C(n1770), .Y(n1759) );
  OAI21X1 U249 ( .A(n1034), .B(n999), .C(n1749), .Y(n1241) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1749) );
  OAI21X1 U251 ( .A(n1035), .B(n999), .C(n1748), .Y(n1240) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1748) );
  OAI21X1 U253 ( .A(n1036), .B(n999), .C(n1747), .Y(n1239) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1747) );
  OAI21X1 U255 ( .A(n1037), .B(n999), .C(n1746), .Y(n1238) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1746) );
  OAI21X1 U257 ( .A(n1038), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1745) );
  OAI21X1 U259 ( .A(n1039), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1744) );
  OAI21X1 U261 ( .A(n1040), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1743) );
  OAI21X1 U263 ( .A(n1041), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1742) );
  NAND3X1 U265 ( .A(n973), .B(n1013), .C(n1741), .Y(n1750) );
  OAI21X1 U266 ( .A(n1042), .B(n998), .C(n1739), .Y(n1233) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1739) );
  OAI21X1 U268 ( .A(n1043), .B(n998), .C(n1738), .Y(n1232) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1738) );
  OAI21X1 U270 ( .A(n1044), .B(n998), .C(n1737), .Y(n1231) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1737) );
  OAI21X1 U272 ( .A(n1045), .B(n998), .C(n1736), .Y(n1230) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1736) );
  OAI21X1 U274 ( .A(n1046), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1735) );
  OAI21X1 U276 ( .A(n1047), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1734) );
  OAI21X1 U278 ( .A(n1048), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1733) );
  OAI21X1 U280 ( .A(n1049), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1732) );
  NAND3X1 U282 ( .A(n1810), .B(n1013), .C(n969), .Y(n1740) );
  OAI21X1 U283 ( .A(n1034), .B(n997), .C(n1730), .Y(n1225) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1730) );
  OAI21X1 U285 ( .A(n1035), .B(n997), .C(n1729), .Y(n1224) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1729) );
  OAI21X1 U287 ( .A(n1036), .B(n997), .C(n1728), .Y(n1223) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1728) );
  OAI21X1 U289 ( .A(n1037), .B(n997), .C(n1727), .Y(n1222) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1727) );
  OAI21X1 U291 ( .A(n1038), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1726) );
  OAI21X1 U293 ( .A(n1039), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1725) );
  OAI21X1 U295 ( .A(n1040), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1724) );
  OAI21X1 U297 ( .A(n1041), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1723) );
  NAND3X1 U299 ( .A(n973), .B(n1013), .C(n1722), .Y(n1731) );
  OAI21X1 U300 ( .A(n1042), .B(n996), .C(n1720), .Y(n1217) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1720) );
  OAI21X1 U302 ( .A(n1043), .B(n996), .C(n1719), .Y(n1216) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1719) );
  OAI21X1 U304 ( .A(n1044), .B(n996), .C(n1718), .Y(n1215) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1718) );
  OAI21X1 U306 ( .A(n1045), .B(n996), .C(n1717), .Y(n1214) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1717) );
  OAI21X1 U308 ( .A(n1046), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1716) );
  OAI21X1 U310 ( .A(n1047), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1715) );
  OAI21X1 U312 ( .A(n1048), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1714) );
  OAI21X1 U314 ( .A(n1049), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1713) );
  NAND3X1 U316 ( .A(n1790), .B(n1013), .C(n969), .Y(n1721) );
  OAI21X1 U317 ( .A(n1034), .B(n995), .C(n1711), .Y(n1209) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1711) );
  OAI21X1 U319 ( .A(n1035), .B(n995), .C(n1710), .Y(n1208) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1710) );
  OAI21X1 U321 ( .A(n1036), .B(n995), .C(n1709), .Y(n1207) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1709) );
  OAI21X1 U323 ( .A(n1037), .B(n995), .C(n1708), .Y(n1206) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1708) );
  OAI21X1 U325 ( .A(n1038), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1707) );
  OAI21X1 U327 ( .A(n1039), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1706) );
  OAI21X1 U329 ( .A(n1040), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1705) );
  OAI21X1 U331 ( .A(n1041), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1704) );
  NAND3X1 U333 ( .A(n973), .B(n1013), .C(n1703), .Y(n1712) );
  OAI21X1 U334 ( .A(n1042), .B(n994), .C(n1701), .Y(n1201) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1701) );
  OAI21X1 U336 ( .A(n1043), .B(n994), .C(n1700), .Y(n1200) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1700) );
  OAI21X1 U338 ( .A(n1044), .B(n994), .C(n1699), .Y(n1199) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1699) );
  OAI21X1 U340 ( .A(n1045), .B(n994), .C(n1698), .Y(n1198) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1698) );
  OAI21X1 U342 ( .A(n1046), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1697) );
  OAI21X1 U344 ( .A(n1047), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1696) );
  OAI21X1 U346 ( .A(n1048), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1695) );
  OAI21X1 U348 ( .A(n1049), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1694) );
  NAND3X1 U350 ( .A(n1810), .B(n1013), .C(n967), .Y(n1702) );
  OAI21X1 U351 ( .A(n1034), .B(n993), .C(n1692), .Y(n1193) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1692) );
  OAI21X1 U353 ( .A(n1035), .B(n993), .C(n1691), .Y(n1192) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1691) );
  OAI21X1 U355 ( .A(n1036), .B(n993), .C(n1690), .Y(n1191) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1690) );
  OAI21X1 U357 ( .A(n1037), .B(n993), .C(n1689), .Y(n1190) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1689) );
  OAI21X1 U359 ( .A(n1038), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1688) );
  OAI21X1 U361 ( .A(n1039), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1687) );
  OAI21X1 U363 ( .A(n1040), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1686) );
  OAI21X1 U365 ( .A(n1041), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1685) );
  NAND3X1 U367 ( .A(n973), .B(n1013), .C(n1684), .Y(n1693) );
  OAI21X1 U368 ( .A(n1042), .B(n992), .C(n1682), .Y(n1185) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1682) );
  OAI21X1 U370 ( .A(n1043), .B(n992), .C(n1681), .Y(n1184) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1681) );
  OAI21X1 U372 ( .A(n1044), .B(n992), .C(n1680), .Y(n1183) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1680) );
  OAI21X1 U374 ( .A(n1045), .B(n992), .C(n1679), .Y(n1182) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1679) );
  OAI21X1 U376 ( .A(n1046), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1678) );
  OAI21X1 U378 ( .A(n1047), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1677) );
  OAI21X1 U380 ( .A(n1048), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1676) );
  OAI21X1 U382 ( .A(n1049), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1675) );
  NAND3X1 U384 ( .A(n1790), .B(n1013), .C(n967), .Y(n1683) );
  OAI21X1 U385 ( .A(n1034), .B(n991), .C(n1673), .Y(n1177) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1673) );
  OAI21X1 U387 ( .A(n1035), .B(n991), .C(n1672), .Y(n1176) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1672) );
  OAI21X1 U389 ( .A(n1036), .B(n991), .C(n1671), .Y(n1175) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1671) );
  OAI21X1 U391 ( .A(n1037), .B(n991), .C(n1670), .Y(n1174) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1670) );
  OAI21X1 U393 ( .A(n1038), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1669) );
  OAI21X1 U395 ( .A(n1039), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1668) );
  OAI21X1 U397 ( .A(n1040), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1667) );
  OAI21X1 U399 ( .A(n1041), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1666) );
  NAND3X1 U401 ( .A(n973), .B(n1013), .C(n1665), .Y(n1674) );
  OAI21X1 U402 ( .A(n1042), .B(n990), .C(n1663), .Y(n1169) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1663) );
  OAI21X1 U404 ( .A(n1043), .B(n989), .C(n1662), .Y(n1168) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1662) );
  OAI21X1 U406 ( .A(n1044), .B(n989), .C(n1661), .Y(n1167) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1661) );
  OAI21X1 U408 ( .A(n1045), .B(n989), .C(n1660), .Y(n1166) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1660) );
  OAI21X1 U410 ( .A(n1046), .B(n989), .C(n1659), .Y(n1165) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1659) );
  OAI21X1 U412 ( .A(n1047), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1658) );
  OAI21X1 U414 ( .A(n1048), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1657) );
  OAI21X1 U416 ( .A(n1049), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1656) );
  NAND3X1 U418 ( .A(n1811), .B(n1012), .C(n1655), .Y(n1664) );
  OAI21X1 U419 ( .A(n1034), .B(n988), .C(n1653), .Y(n1161) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1653) );
  OAI21X1 U421 ( .A(n1035), .B(n988), .C(n1652), .Y(n1160) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1652) );
  OAI21X1 U423 ( .A(n1036), .B(n988), .C(n1651), .Y(n1159) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1651) );
  OAI21X1 U425 ( .A(n1037), .B(n988), .C(n1650), .Y(n1158) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1650) );
  OAI21X1 U427 ( .A(n1038), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1649) );
  OAI21X1 U429 ( .A(n1039), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1648) );
  OAI21X1 U431 ( .A(n1040), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1647) );
  OAI21X1 U433 ( .A(n1041), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1646) );
  NAND3X1 U435 ( .A(n973), .B(n1012), .C(n1645), .Y(n1654) );
  OAI21X1 U436 ( .A(n1042), .B(n987), .C(n1643), .Y(n1153) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1643) );
  OAI21X1 U438 ( .A(n1043), .B(n986), .C(n1642), .Y(n1152) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1642) );
  OAI21X1 U440 ( .A(n1044), .B(n986), .C(n1641), .Y(n1151) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1641) );
  OAI21X1 U442 ( .A(n1045), .B(n986), .C(n1640), .Y(n1150) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1640) );
  OAI21X1 U444 ( .A(n1046), .B(n986), .C(n1639), .Y(n1149) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1639) );
  OAI21X1 U446 ( .A(n1047), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1638) );
  OAI21X1 U448 ( .A(n1048), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1637) );
  OAI21X1 U450 ( .A(n1049), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1636) );
  NAND3X1 U452 ( .A(n1811), .B(n1012), .C(n1635), .Y(n1644) );
  OAI21X1 U453 ( .A(n1034), .B(n985), .C(n1632), .Y(n1145) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1632) );
  OAI21X1 U455 ( .A(n1035), .B(n985), .C(n1631), .Y(n1144) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1631) );
  OAI21X1 U457 ( .A(n1036), .B(n985), .C(n1630), .Y(n1143) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1630) );
  OAI21X1 U459 ( .A(n1037), .B(n985), .C(n1629), .Y(n1142) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1629) );
  OAI21X1 U461 ( .A(n1038), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1628) );
  OAI21X1 U463 ( .A(n1039), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1627) );
  OAI21X1 U465 ( .A(n1040), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1626) );
  OAI21X1 U467 ( .A(n1041), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1625) );
  NAND3X1 U469 ( .A(n973), .B(n1012), .C(n1624), .Y(n1633) );
  OAI21X1 U470 ( .A(n1042), .B(n984), .C(n1622), .Y(n1137) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1622) );
  OAI21X1 U472 ( .A(n1043), .B(n983), .C(n1621), .Y(n1136) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1621) );
  OAI21X1 U474 ( .A(n1044), .B(n983), .C(n1620), .Y(n1135) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1620) );
  OAI21X1 U476 ( .A(n1045), .B(n983), .C(n1619), .Y(n1134) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1619) );
  OAI21X1 U478 ( .A(n1046), .B(n983), .C(n1618), .Y(n1133) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1618) );
  OAI21X1 U480 ( .A(n1047), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1617) );
  OAI21X1 U482 ( .A(n1048), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1616) );
  OAI21X1 U484 ( .A(n1049), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1615) );
  NAND3X1 U486 ( .A(n1770), .B(n1012), .C(n1655), .Y(n1623) );
  OAI21X1 U487 ( .A(n1034), .B(n982), .C(n1613), .Y(n1129) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1613) );
  OAI21X1 U489 ( .A(n1035), .B(n982), .C(n1612), .Y(n1128) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1612) );
  OAI21X1 U491 ( .A(n1036), .B(n982), .C(n1611), .Y(n1127) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1611) );
  OAI21X1 U493 ( .A(n1037), .B(n982), .C(n1610), .Y(n1126) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1610) );
  OAI21X1 U495 ( .A(n1038), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1609) );
  OAI21X1 U497 ( .A(n1039), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1608) );
  OAI21X1 U499 ( .A(n1040), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1607) );
  OAI21X1 U501 ( .A(n1041), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1606) );
  NAND3X1 U503 ( .A(n973), .B(n1012), .C(n1605), .Y(n1614) );
  OAI21X1 U504 ( .A(n1042), .B(n981), .C(n1603), .Y(n1121) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1603) );
  OAI21X1 U506 ( .A(n1043), .B(n980), .C(n1602), .Y(n1120) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1602) );
  OAI21X1 U508 ( .A(n1044), .B(n980), .C(n1601), .Y(n1119) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1601) );
  OAI21X1 U510 ( .A(n1045), .B(n980), .C(n1600), .Y(n1118) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1600) );
  OAI21X1 U512 ( .A(n1046), .B(n980), .C(n1599), .Y(n1117) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1599) );
  OAI21X1 U514 ( .A(n1047), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1598) );
  OAI21X1 U516 ( .A(n1048), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1597) );
  OAI21X1 U518 ( .A(n1049), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1596) );
  NAND3X1 U520 ( .A(n1770), .B(n1012), .C(n1635), .Y(n1604) );
  OAI21X1 U521 ( .A(n1034), .B(n979), .C(n1593), .Y(n1113) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1593) );
  OAI21X1 U523 ( .A(n1035), .B(n979), .C(n1592), .Y(n1112) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1592) );
  OAI21X1 U525 ( .A(n1036), .B(n979), .C(n1591), .Y(n1111) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1591) );
  OAI21X1 U527 ( .A(n1037), .B(n979), .C(n1590), .Y(n1110) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1590) );
  OAI21X1 U529 ( .A(n1038), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1589) );
  OAI21X1 U531 ( .A(n1039), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1588) );
  OAI21X1 U533 ( .A(n1040), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1587) );
  OAI21X1 U535 ( .A(n1041), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1586) );
  NAND3X1 U537 ( .A(n973), .B(n1012), .C(n1585), .Y(n1594) );
  OAI21X1 U538 ( .A(n1042), .B(n978), .C(n1583), .Y(n1105) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1583) );
  OAI21X1 U540 ( .A(n1043), .B(n978), .C(n1582), .Y(n1104) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1582) );
  OAI21X1 U542 ( .A(n1044), .B(n978), .C(n1581), .Y(n1103) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1581) );
  OAI21X1 U544 ( .A(n1045), .B(n978), .C(n1580), .Y(n1102) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1580) );
  OAI21X1 U546 ( .A(n1046), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1579) );
  OAI21X1 U548 ( .A(n1047), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1578) );
  OAI21X1 U550 ( .A(n1048), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1577) );
  OAI21X1 U552 ( .A(n1049), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1576) );
  NAND3X1 U554 ( .A(n969), .B(n1012), .C(n1655), .Y(n1584) );
  OAI21X1 U555 ( .A(n1034), .B(n977), .C(n1574), .Y(n1097) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1574) );
  OAI21X1 U557 ( .A(n1035), .B(n977), .C(n1573), .Y(n1096) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1573) );
  OAI21X1 U559 ( .A(n1036), .B(n977), .C(n1572), .Y(n1095) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1572) );
  OAI21X1 U561 ( .A(n1037), .B(n977), .C(n1571), .Y(n1094) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1571) );
  OAI21X1 U563 ( .A(n1038), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1570) );
  OAI21X1 U565 ( .A(n1039), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1569) );
  OAI21X1 U567 ( .A(n1040), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1568) );
  OAI21X1 U569 ( .A(n1041), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1567) );
  NAND3X1 U571 ( .A(n973), .B(n1012), .C(n1566), .Y(n1575) );
  OAI21X1 U572 ( .A(n1042), .B(n976), .C(n1564), .Y(n1089) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1564) );
  OAI21X1 U574 ( .A(n1043), .B(n976), .C(n1563), .Y(n1088) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1563) );
  OAI21X1 U576 ( .A(n1044), .B(n976), .C(n1562), .Y(n1087) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1562) );
  OAI21X1 U578 ( .A(n1045), .B(n976), .C(n1561), .Y(n1086) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1561) );
  OAI21X1 U580 ( .A(n1046), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1560) );
  OAI21X1 U582 ( .A(n1047), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1559) );
  OAI21X1 U584 ( .A(n1048), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1558) );
  OAI21X1 U586 ( .A(n1049), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1557) );
  NAND3X1 U588 ( .A(n969), .B(n1012), .C(n1635), .Y(n1565) );
  OAI21X1 U590 ( .A(n1034), .B(n975), .C(n1554), .Y(n1081) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1554) );
  OAI21X1 U592 ( .A(n1035), .B(n975), .C(n1553), .Y(n1080) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1553) );
  OAI21X1 U594 ( .A(n1036), .B(n975), .C(n1552), .Y(n1079) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1552) );
  OAI21X1 U596 ( .A(n1037), .B(n975), .C(n1551), .Y(n1078) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1551) );
  OAI21X1 U598 ( .A(n1038), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1550) );
  OAI21X1 U600 ( .A(n1039), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1549) );
  OAI21X1 U602 ( .A(n1040), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1548) );
  OAI21X1 U604 ( .A(n1041), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1547) );
  NAND3X1 U606 ( .A(n973), .B(n1012), .C(n1546), .Y(n1555) );
  OAI21X1 U607 ( .A(n1042), .B(n974), .C(n1544), .Y(n1073) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1544) );
  OAI21X1 U609 ( .A(n1043), .B(n974), .C(n1543), .Y(n1072) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1543) );
  OAI21X1 U611 ( .A(n1044), .B(n974), .C(n1542), .Y(n1071) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1542) );
  OAI21X1 U613 ( .A(n1045), .B(n974), .C(n1541), .Y(n1070) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1541) );
  OAI21X1 U615 ( .A(n1046), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1540) );
  OAI21X1 U617 ( .A(n1047), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1539) );
  OAI21X1 U619 ( .A(n1048), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1538) );
  OAI21X1 U621 ( .A(n1049), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1537) );
  NAND3X1 U623 ( .A(n967), .B(n1012), .C(n1655), .Y(n1545) );
  OAI21X1 U624 ( .A(n1034), .B(n8), .C(n1536), .Y(n1065) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1536) );
  OAI21X1 U626 ( .A(n1035), .B(n8), .C(n1535), .Y(n1064) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1535) );
  OAI21X1 U628 ( .A(n1036), .B(n8), .C(n1534), .Y(n1063) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1534) );
  OAI21X1 U630 ( .A(n1037), .B(n8), .C(n1533), .Y(n1062) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1533) );
  OAI21X1 U632 ( .A(n1038), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1532) );
  OAI21X1 U634 ( .A(n1039), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1531) );
  OAI21X1 U636 ( .A(n1040), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1530) );
  OAI21X1 U638 ( .A(n1041), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1529) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1822) );
  OAI21X1 U642 ( .A(n1042), .B(n972), .C(n1526), .Y(n1057) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1526) );
  OAI21X1 U644 ( .A(n1043), .B(n972), .C(n1525), .Y(n1056) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1525) );
  OAI21X1 U646 ( .A(n1044), .B(n972), .C(n1524), .Y(n1055) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1524) );
  OAI21X1 U648 ( .A(n1045), .B(n972), .C(n1523), .Y(n1054) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1523) );
  OAI21X1 U650 ( .A(n1046), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1522) );
  OAI21X1 U652 ( .A(n1047), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1521) );
  OAI21X1 U654 ( .A(n1048), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1520) );
  OAI21X1 U656 ( .A(n1049), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1519) );
  NAND3X1 U658 ( .A(n967), .B(n1013), .C(n1635), .Y(n1527) );
  NOR3X1 U661 ( .A(n1515), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1516) );
  NOR3X1 U662 ( .A(n1514), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1517) );
  AOI21X1 U663 ( .A(n461), .B(n1513), .C(n963), .Y(n1842) );
  OAI21X1 U665 ( .A(rd), .B(n1512), .C(wr), .Y(n1513) );
  NAND3X1 U667 ( .A(n1511), .B(n1029), .C(n1510), .Y(n1512) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1510) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1511) );
  AOI21X1 U670 ( .A(n448), .B(n1508), .C(n1028), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1507), .C(n4), .Y(n1508) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1790), .C(\mem<0><1> ), .D(n1635), .Y(
        n1505) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1810), .C(\mem<2><1> ), .D(n1655), .Y(
        n1506) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1790), .C(\mem<4><1> ), .D(n1635), .Y(
        n1503) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1810), .C(\mem<6><1> ), .D(n1655), .Y(
        n1504) );
  AOI22X1 U678 ( .A(n1595), .B(n892), .C(n1634), .D(n932), .Y(n1509) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1790), .C(\mem<12><1> ), .D(n1635), .Y(
        n1501) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1810), .C(\mem<14><1> ), .D(n1655), .Y(
        n1502) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1790), .C(\mem<8><1> ), .D(n1635), .Y(
        n1499) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1810), .C(\mem<10><1> ), .D(n1655), .Y(
        n1500) );
  AOI21X1 U685 ( .A(n447), .B(n1497), .C(n1028), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1495), .C(n949), .Y(n1497) );
  AOI21X1 U687 ( .A(n1493), .B(n1492), .C(n971), .Y(n1494) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1790), .C(\mem<0><0> ), .D(n1635), .Y(
        n1492) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1810), .C(\mem<2><0> ), .D(n1655), .Y(
        n1493) );
  AOI21X1 U690 ( .A(n1491), .B(n1490), .C(n970), .Y(n1496) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1790), .C(\mem<4><0> ), .D(n1635), .Y(
        n1490) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1810), .C(\mem<6><0> ), .D(n1655), .Y(
        n1491) );
  AOI22X1 U693 ( .A(n1595), .B(n890), .C(n1634), .D(n930), .Y(n1498) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1790), .C(\mem<12><0> ), .D(n1635), .Y(
        n1488) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1810), .C(\mem<14><0> ), .D(n1655), .Y(
        n1489) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1790), .C(\mem<8><0> ), .D(n1635), .Y(
        n1486) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1810), .C(\mem<10><0> ), .D(n1655), .Y(
        n1487) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1485) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1684), .C(\mem<19><7> ), .D(n1703), .Y(
        n1480) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1722), .C(\mem<23><7> ), .D(n1741), .Y(
        n1481) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1760), .C(\mem<27><7> ), .D(n1780), .Y(
        n1483) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1800), .C(\mem<31><7> ), .D(n1821), .Y(
        n1484) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1528), .C(\mem<3><7> ), .D(n1546), .Y(
        n1475) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1566), .C(\mem<7><7> ), .D(n1585), .Y(
        n1476) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1605), .C(\mem<11><7> ), .D(n1624), .Y(
        n1478) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1645), .C(\mem<15><7> ), .D(n1665), .Y(
        n1479) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1474) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1684), .C(\mem<19><6> ), .D(n1703), .Y(
        n1469) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1722), .C(\mem<23><6> ), .D(n1741), .Y(
        n1470) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1760), .C(\mem<27><6> ), .D(n1780), .Y(
        n1472) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1800), .C(\mem<31><6> ), .D(n1821), .Y(
        n1473) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1528), .C(\mem<3><6> ), .D(n1546), .Y(
        n1464) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1566), .C(\mem<7><6> ), .D(n1585), .Y(
        n1465) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1605), .C(\mem<11><6> ), .D(n1624), .Y(
        n1467) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1645), .C(\mem<15><6> ), .D(n1665), .Y(
        n1468) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1463) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1684), .C(\mem<19><5> ), .D(n1703), .Y(
        n1458) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1722), .C(\mem<23><5> ), .D(n1741), .Y(
        n1459) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1760), .C(\mem<27><5> ), .D(n1780), .Y(
        n1461) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1800), .C(\mem<31><5> ), .D(n1821), .Y(
        n1462) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1528), .C(\mem<3><5> ), .D(n1546), .Y(
        n1453) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1566), .C(\mem<7><5> ), .D(n1585), .Y(
        n1454) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1605), .C(\mem<11><5> ), .D(n1624), .Y(
        n1456) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1645), .C(\mem<15><5> ), .D(n1665), .Y(
        n1457) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1452) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1684), .C(\mem<19><4> ), .D(n1703), .Y(
        n1447) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1722), .C(\mem<23><4> ), .D(n1741), .Y(
        n1448) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1760), .C(\mem<27><4> ), .D(n1780), .Y(
        n1450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1800), .C(\mem<31><4> ), .D(n1821), .Y(
        n1451) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1528), .C(\mem<3><4> ), .D(n1546), .Y(
        n1442) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1566), .C(\mem<7><4> ), .D(n1585), .Y(
        n1443) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1605), .C(\mem<11><4> ), .D(n1624), .Y(
        n1445) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1645), .C(\mem<15><4> ), .D(n1665), .Y(
        n1446) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1441) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1684), .C(\mem<19><3> ), .D(n1703), .Y(
        n1436) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1722), .C(\mem<23><3> ), .D(n1741), .Y(
        n1437) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1760), .C(\mem<27><3> ), .D(n1780), .Y(
        n1439) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1800), .C(\mem<31><3> ), .D(n1821), .Y(
        n1440) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1528), .C(\mem<3><3> ), .D(n1546), .Y(
        n1431) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1566), .C(\mem<7><3> ), .D(n1585), .Y(
        n1432) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1605), .C(\mem<11><3> ), .D(n1624), .Y(
        n1434) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1645), .C(\mem<15><3> ), .D(n1665), .Y(
        n1435) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1430) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1684), .C(\mem<19><2> ), .D(n1703), .Y(
        n1425) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1722), .C(\mem<23><2> ), .D(n1741), .Y(
        n1426) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1760), .C(\mem<27><2> ), .D(n1780), .Y(
        n1428) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1800), .C(\mem<31><2> ), .D(n1821), .Y(
        n1429) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1528), .C(\mem<3><2> ), .D(n1546), .Y(
        n1420) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1566), .C(\mem<7><2> ), .D(n1585), .Y(
        n1421) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1605), .C(\mem<11><2> ), .D(n1624), .Y(
        n1423) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1645), .C(\mem<15><2> ), .D(n1665), .Y(
        n1424) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1419) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1684), .C(\mem<19><1> ), .D(n1703), .Y(
        n1414) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1722), .C(\mem<23><1> ), .D(n1741), .Y(
        n1415) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1760), .C(\mem<27><1> ), .D(n1780), .Y(
        n1417) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1800), .C(\mem<31><1> ), .D(n1821), .Y(
        n1418) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1528), .C(\mem<3><1> ), .D(n1546), .Y(
        n1409) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1566), .C(\mem<7><1> ), .D(n1585), .Y(
        n1410) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1605), .C(\mem<11><1> ), .D(n1624), .Y(
        n1412) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1645), .C(\mem<15><1> ), .D(n1665), .Y(
        n1413) );
  AOI21X1 U777 ( .A(n435), .B(n1407), .C(n1028), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1405), .C(n948), .Y(n1407) );
  AOI21X1 U779 ( .A(n1403), .B(n1402), .C(n971), .Y(n1404) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1790), .C(\mem<0><7> ), .D(n1635), .Y(
        n1402) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1810), .C(\mem<2><7> ), .D(n1655), .Y(
        n1403) );
  AOI21X1 U782 ( .A(n1401), .B(n1400), .C(n970), .Y(n1406) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1790), .C(\mem<4><7> ), .D(n1635), .Y(
        n1400) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1810), .C(\mem<6><7> ), .D(n1655), .Y(
        n1401) );
  AOI22X1 U785 ( .A(n1595), .B(n888), .C(n1634), .D(n928), .Y(n1408) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1790), .C(\mem<12><7> ), .D(n1635), .Y(
        n1398) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1810), .C(\mem<14><7> ), .D(n1655), .Y(
        n1399) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1790), .C(\mem<8><7> ), .D(n1635), .Y(
        n1396) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1810), .C(\mem<10><7> ), .D(n1655), .Y(
        n1397) );
  AOI21X1 U792 ( .A(n434), .B(n1394), .C(n1028), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1392), .C(n947), .Y(n1394) );
  AOI21X1 U794 ( .A(n1390), .B(n1389), .C(n971), .Y(n1391) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1790), .C(\mem<0><6> ), .D(n1635), .Y(
        n1389) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1810), .C(\mem<2><6> ), .D(n1655), .Y(
        n1390) );
  AOI21X1 U797 ( .A(n1388), .B(n1387), .C(n970), .Y(n1393) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1790), .C(\mem<4><6> ), .D(n1635), .Y(
        n1387) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1810), .C(\mem<6><6> ), .D(n1655), .Y(
        n1388) );
  AOI22X1 U800 ( .A(n1595), .B(n886), .C(n1634), .D(n926), .Y(n1395) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1790), .C(\mem<12><6> ), .D(n1635), .Y(
        n1385) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1810), .C(\mem<14><6> ), .D(n1655), .Y(
        n1386) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1790), .C(\mem<8><6> ), .D(n1635), .Y(
        n1383) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1810), .C(\mem<10><6> ), .D(n1655), .Y(
        n1384) );
  AOI21X1 U807 ( .A(n422), .B(n1381), .C(n1028), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1379), .C(n946), .Y(n1381) );
  AOI21X1 U809 ( .A(n1377), .B(n1376), .C(n971), .Y(n1378) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1790), .C(\mem<0><5> ), .D(n1635), .Y(
        n1376) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1810), .C(\mem<2><5> ), .D(n1655), .Y(
        n1377) );
  AOI21X1 U812 ( .A(n1375), .B(n1374), .C(n970), .Y(n1380) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1790), .C(\mem<4><5> ), .D(n1635), .Y(
        n1374) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1810), .C(\mem<6><5> ), .D(n1655), .Y(
        n1375) );
  AOI22X1 U815 ( .A(n1595), .B(n884), .C(n1634), .D(n924), .Y(n1382) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1790), .C(\mem<12><5> ), .D(n1635), .Y(
        n1372) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1810), .C(\mem<14><5> ), .D(n1655), .Y(
        n1373) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1790), .C(\mem<8><5> ), .D(n1635), .Y(
        n1370) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1810), .C(\mem<10><5> ), .D(n1655), .Y(
        n1371) );
  AOI21X1 U822 ( .A(n421), .B(n1368), .C(n1028), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1366), .C(n945), .Y(n1368) );
  AOI21X1 U824 ( .A(n1364), .B(n1363), .C(n971), .Y(n1365) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1790), .C(\mem<0><4> ), .D(n1635), .Y(
        n1363) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1810), .C(\mem<2><4> ), .D(n1655), .Y(
        n1364) );
  AOI21X1 U827 ( .A(n1362), .B(n1361), .C(n970), .Y(n1367) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1790), .C(\mem<4><4> ), .D(n1635), .Y(
        n1361) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1810), .C(\mem<6><4> ), .D(n1655), .Y(
        n1362) );
  AOI22X1 U830 ( .A(n1595), .B(n882), .C(n1634), .D(n922), .Y(n1369) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1790), .C(\mem<12><4> ), .D(n1635), .Y(
        n1359) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1810), .C(\mem<14><4> ), .D(n1655), .Y(
        n1360) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1790), .C(\mem<8><4> ), .D(n1635), .Y(
        n1357) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1810), .C(\mem<10><4> ), .D(n1655), .Y(
        n1358) );
  AOI21X1 U837 ( .A(n409), .B(n1355), .C(n1028), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1353), .C(n944), .Y(n1355) );
  AOI21X1 U839 ( .A(n1351), .B(n1350), .C(n971), .Y(n1352) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1790), .C(\mem<0><3> ), .D(n1635), .Y(
        n1350) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1810), .C(\mem<2><3> ), .D(n1655), .Y(
        n1351) );
  AOI21X1 U842 ( .A(n1349), .B(n1348), .C(n970), .Y(n1354) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1790), .C(\mem<4><3> ), .D(n1635), .Y(
        n1348) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1810), .C(\mem<6><3> ), .D(n1655), .Y(
        n1349) );
  AOI22X1 U845 ( .A(n1595), .B(n880), .C(n1634), .D(n920), .Y(n1356) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1790), .C(\mem<12><3> ), .D(n1635), .Y(
        n1346) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1810), .C(\mem<14><3> ), .D(n1655), .Y(
        n1347) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1790), .C(\mem<8><3> ), .D(n1635), .Y(
        n1344) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1810), .C(\mem<10><3> ), .D(n1655), .Y(
        n1345) );
  AOI21X1 U852 ( .A(n408), .B(n1342), .C(n1028), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1340), .C(n943), .Y(n1342) );
  AOI21X1 U854 ( .A(n1338), .B(n1337), .C(n971), .Y(n1339) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1790), .C(\mem<0><2> ), .D(n1635), .Y(
        n1337) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1810), .C(\mem<2><2> ), .D(n1655), .Y(
        n1338) );
  AOI21X1 U857 ( .A(n1336), .B(n1335), .C(n970), .Y(n1341) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1790), .C(\mem<4><2> ), .D(n1635), .Y(
        n1335) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1810), .C(\mem<6><2> ), .D(n1655), .Y(
        n1336) );
  AOI22X1 U860 ( .A(n1595), .B(n878), .C(n1634), .D(n918), .Y(n1343) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1790), .C(\mem<12><2> ), .D(n1635), .Y(
        n1333) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1810), .C(\mem<14><2> ), .D(n1655), .Y(
        n1334) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1790), .C(\mem<8><2> ), .D(n1635), .Y(
        n1331) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1810), .C(\mem<10><2> ), .D(n1655), .Y(
        n1332) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1330) );
  NOR2X1 U868 ( .A(n1033), .B(\addr_1c<4> ), .Y(n1329) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1328) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1684), .C(\mem<19><0> ), .D(n1703), .Y(
        n1323) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1722), .C(\mem<23><0> ), .D(n1741), .Y(
        n1324) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1760), .C(\mem<27><0> ), .D(n1780), .Y(
        n1326) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1800), .C(\mem<31><0> ), .D(n1821), .Y(
        n1327) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1528), .C(\mem<3><0> ), .D(n1546), .Y(
        n1316) );
  NAND2X1 U877 ( .A(n1031), .B(n1032), .Y(n1518) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1566), .C(\mem<7><0> ), .D(n1585), .Y(
        n1317) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1032), .Y(n1556) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1605), .C(\mem<11><0> ), .D(n1624), .Y(
        n1319) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1645), .C(\mem<15><0> ), .D(n1665), .Y(
        n1320) );
  dff_101 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1015) );
  dff_100 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1016) );
  dff_99 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1016)
         );
  dff_98 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1016)
         );
  dff_97 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1016)
         );
  dff_96 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1016)
         );
  dff_95 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1016)
         );
  dff_94 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1016)
         );
  dff_93 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1016)
         );
  dff_92 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1016)
         );
  dff_91 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1015)
         );
  dff_90 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1015)
         );
  dff_89 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1015) );
  dff_88 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1015) );
  dff_87 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1015) );
  dff_86 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1015) );
  dff_85 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1015) );
  dff_84 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1015) );
  dff_83 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1015) );
  dff_82 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1015) );
  dff_81 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1015) );
  dff_80 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1015) );
  dff_79 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1015) );
  dff_78 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1015) );
  dff_77 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1015) );
  dff_76 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1015) );
  dff_75 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1015) );
  dff_74 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1015) );
  dff_73 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1015) );
  dff_72 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1015) );
  dff_71 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1015) );
  dff_70 \reg2[0]  ( .q(\data_out<0> ), .d(n1025), .clk(clk), .rst(n1016) );
  dff_69 \reg2[1]  ( .q(\data_out<1> ), .d(n1024), .clk(clk), .rst(n1016) );
  dff_68 \reg2[2]  ( .q(\data_out<2> ), .d(n1023), .clk(clk), .rst(n1016) );
  dff_67 \reg2[3]  ( .q(\data_out<3> ), .d(n1022), .clk(clk), .rst(n1016) );
  dff_66 \reg2[4]  ( .q(\data_out<4> ), .d(n1021), .clk(clk), .rst(n1016) );
  dff_65 \reg2[5]  ( .q(\data_out<5> ), .d(n1020), .clk(clk), .rst(n1016) );
  dff_64 \reg2[6]  ( .q(\data_out<6> ), .d(n1019), .clk(clk), .rst(n1015) );
  dff_63 \reg2[7]  ( .q(\data_out<7> ), .d(n1018), .clk(clk), .rst(n1015) );
  dff_62 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1015) );
  dff_61 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1015) );
  dff_60 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1015) );
  dff_59 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1015) );
  dff_58 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1015) );
  dff_57 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1015) );
  dff_56 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1015) );
  dff_55 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1015) );
  dff_54 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1015) );
  dff_53 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1015) );
  dff_52 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1015) );
  dff_51 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1016) );
  OR2X1 U2 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1514) );
  AND2X1 U3 ( .A(\addr_1c<4> ), .B(n1528), .Y(n1831) );
  INVX1 U4 ( .A(\addr_1c<3> ), .Y(n1033) );
  INVX1 U5 ( .A(\addr_1c<2> ), .Y(n1032) );
  INVX1 U6 ( .A(wr1), .Y(n1029) );
  OR2X1 U7 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1515) );
  INVX1 U8 ( .A(\addr_1c<0> ), .Y(n1030) );
  AND2X1 U23 ( .A(n1030), .B(n1033), .Y(n1314) );
  AND2X1 U24 ( .A(\addr_1c<0> ), .B(n1033), .Y(n1315) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1322) );
  AND2X1 U26 ( .A(\addr_1c<3> ), .B(n1030), .Y(n1321) );
  INVX1 U27 ( .A(\addr_1c<1> ), .Y(n1031) );
  AND2X1 U28 ( .A(n1595), .B(n1322), .Y(n1780) );
  AND2X1 U29 ( .A(n1595), .B(n1321), .Y(n1760) );
  AND2X1 U35 ( .A(n940), .B(n1322), .Y(n1741) );
  AND2X1 U36 ( .A(n940), .B(n1321), .Y(n1722) );
  AND2X1 U37 ( .A(n1322), .B(n950), .Y(n1703) );
  AND2X1 U38 ( .A(n1321), .B(n950), .Y(n1684) );
  AND2X1 U39 ( .A(n1315), .B(n1595), .Y(n1624) );
  AND2X1 U40 ( .A(n1595), .B(n1314), .Y(n1605) );
  AND2X1 U41 ( .A(n1315), .B(n940), .Y(n1585) );
  AND2X1 U42 ( .A(n940), .B(n1314), .Y(n1566) );
  OR2X1 U43 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U44 ( .A(n1315), .B(n950), .Y(n1546) );
  OR2X1 U46 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U47 ( .A(n1634), .B(n1314), .Y(n1645) );
  AND2X1 U48 ( .A(n1315), .B(n1634), .Y(n1665) );
  AND2X1 U49 ( .A(n1321), .B(n1634), .Y(n1800) );
  AND2X1 U50 ( .A(\addr_1c<2> ), .B(n1031), .Y(n1595) );
  AND2X1 U51 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1634) );
  BUFX2 U52 ( .A(n961), .Y(n1010) );
  BUFX2 U53 ( .A(n961), .Y(n1009) );
  BUFX2 U54 ( .A(n960), .Y(n1007) );
  BUFX2 U55 ( .A(n960), .Y(n1006) );
  BUFX2 U56 ( .A(n959), .Y(n1004) );
  BUFX2 U57 ( .A(n959), .Y(n1003) );
  BUFX2 U58 ( .A(n958), .Y(n1001) );
  BUFX2 U59 ( .A(n958), .Y(n1000) );
  BUFX2 U60 ( .A(n957), .Y(n990) );
  BUFX2 U61 ( .A(n957), .Y(n989) );
  BUFX2 U62 ( .A(n956), .Y(n987) );
  BUFX2 U63 ( .A(n956), .Y(n986) );
  BUFX2 U64 ( .A(n955), .Y(n984) );
  BUFX2 U65 ( .A(n955), .Y(n983) );
  BUFX2 U66 ( .A(n954), .Y(n981) );
  BUFX2 U67 ( .A(n954), .Y(n980) );
  INVX1 U68 ( .A(\data_in_1c<0> ), .Y(n1034) );
  INVX1 U69 ( .A(\data_in_1c<1> ), .Y(n1035) );
  INVX1 U70 ( .A(\data_in_1c<2> ), .Y(n1036) );
  INVX1 U71 ( .A(\data_in_1c<3> ), .Y(n1037) );
  INVX1 U72 ( .A(\data_in_1c<4> ), .Y(n1038) );
  INVX1 U73 ( .A(\data_in_1c<5> ), .Y(n1039) );
  INVX1 U74 ( .A(\data_in_1c<6> ), .Y(n1040) );
  INVX1 U75 ( .A(\data_in_1c<7> ), .Y(n1041) );
  INVX1 U76 ( .A(\data_in_1c<8> ), .Y(n1042) );
  INVX1 U77 ( .A(\data_in_1c<9> ), .Y(n1043) );
  INVX1 U78 ( .A(\data_in_1c<10> ), .Y(n1044) );
  INVX1 U79 ( .A(\data_in_1c<11> ), .Y(n1045) );
  INVX1 U80 ( .A(\data_in_1c<12> ), .Y(n1046) );
  INVX1 U81 ( .A(\data_in_1c<13> ), .Y(n1047) );
  INVX1 U82 ( .A(\data_in_1c<14> ), .Y(n1048) );
  INVX1 U83 ( .A(\data_in_1c<15> ), .Y(n1049) );
  AND2X1 U84 ( .A(n1831), .B(\mem<32><0> ), .Y(n1495) );
  AND2X1 U85 ( .A(n1831), .B(\mem<32><1> ), .Y(n1507) );
  AND2X1 U86 ( .A(n1831), .B(\mem<32><2> ), .Y(n1340) );
  AND2X1 U87 ( .A(n1831), .B(\mem<32><3> ), .Y(n1353) );
  AND2X1 U88 ( .A(n1831), .B(\mem<32><4> ), .Y(n1366) );
  AND2X1 U89 ( .A(n1831), .B(\mem<32><5> ), .Y(n1379) );
  AND2X1 U90 ( .A(n1831), .B(\mem<32><6> ), .Y(n1392) );
  AND2X1 U91 ( .A(n1831), .B(\mem<32><7> ), .Y(n1405) );
  INVX1 U92 ( .A(rd1), .Y(n1028) );
  INVX1 U93 ( .A(n1328), .Y(n1025) );
  INVX1 U129 ( .A(n1419), .Y(n1024) );
  INVX1 U589 ( .A(n1430), .Y(n1023) );
  INVX1 U640 ( .A(n1441), .Y(n1022) );
  INVX1 U659 ( .A(n1452), .Y(n1021) );
  INVX1 U660 ( .A(n1463), .Y(n1020) );
  INVX1 U664 ( .A(n1474), .Y(n1019) );
  INVX1 U666 ( .A(n1485), .Y(n1018) );
  INVX2 U672 ( .A(n1017), .Y(n1015) );
  INVX1 U675 ( .A(n1832), .Y(n1014) );
  AND2X1 U679 ( .A(wr1), .B(n1017), .Y(n1832) );
  INVX1 U682 ( .A(rst), .Y(n1017) );
  AND2X1 U694 ( .A(n1634), .B(n964), .Y(n1811) );
  INVX1 U697 ( .A(n1014), .Y(n1012) );
  AND2X1 U701 ( .A(n1595), .B(n964), .Y(n1770) );
  INVX1 U706 ( .A(n1014), .Y(n1013) );
  AND2X1 U712 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U717 ( .A(n1), .Y(n2) );
  AND2X1 U723 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U728 ( .A(n3), .Y(n4) );
  AND2X1 U734 ( .A(n1821), .B(n189), .Y(n5) );
  INVX1 U739 ( .A(n5), .Y(n6) );
  AND2X1 U745 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U750 ( .A(n7), .Y(n8) );
  OR2X1 U756 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U761 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U767 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U772 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U786 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U789 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U801 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U804 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U816 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U819 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U831 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U834 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U846 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U849 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U861 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U864 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U870 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U875 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U882 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U883 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U884 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U885 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U886 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U887 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U888 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U889 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U890 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U891 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U892 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U893 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U894 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U895 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U896 ( .A(n973), .B(n1832), .Y(n189) );
  AND2X1 U897 ( .A(n1832), .B(n1528), .Y(n289) );
  INVX1 U898 ( .A(n1017), .Y(n1016) );
  AND2X1 U899 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U900 ( .A(n348), .Y(n372) );
  AND2X1 U901 ( .A(n950), .B(n952), .Y(n379) );
  INVX1 U902 ( .A(n379), .Y(n381) );
  AND2X1 U903 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U904 ( .A(n386), .Y(n387) );
  AND2X1 U905 ( .A(n950), .B(n951), .Y(n401) );
  INVX1 U906 ( .A(n401), .Y(n402) );
  BUFX2 U907 ( .A(n1343), .Y(n408) );
  BUFX2 U908 ( .A(n1356), .Y(n409) );
  BUFX2 U909 ( .A(n1369), .Y(n421) );
  BUFX2 U910 ( .A(n1382), .Y(n422) );
  BUFX2 U911 ( .A(n1395), .Y(n434) );
  BUFX2 U912 ( .A(n1408), .Y(n435) );
  BUFX2 U913 ( .A(n1498), .Y(n447) );
  BUFX2 U914 ( .A(n1509), .Y(n448) );
  AND2X2 U915 ( .A(rd), .B(n1512), .Y(n460) );
  INVX1 U916 ( .A(n460), .Y(n461) );
  INVX1 U917 ( .A(n1318), .Y(n473) );
  INVX1 U918 ( .A(n1319), .Y(n474) );
  INVX1 U919 ( .A(n1320), .Y(n486) );
  INVX1 U920 ( .A(n1411), .Y(n487) );
  INVX1 U921 ( .A(n1412), .Y(n507) );
  INVX1 U922 ( .A(n1413), .Y(n508) );
  INVX1 U923 ( .A(n1422), .Y(n522) );
  INVX1 U924 ( .A(n1423), .Y(n523) );
  INVX1 U925 ( .A(n1424), .Y(n537) );
  INVX1 U926 ( .A(n1433), .Y(n538) );
  INVX1 U927 ( .A(n1434), .Y(n552) );
  INVX1 U928 ( .A(n1435), .Y(n553) );
  INVX1 U929 ( .A(n1444), .Y(n567) );
  INVX1 U930 ( .A(n1445), .Y(n568) );
  INVX1 U931 ( .A(n1446), .Y(n582) );
  INVX1 U932 ( .A(n1455), .Y(n583) );
  INVX1 U933 ( .A(n1456), .Y(n591) );
  INVX1 U934 ( .A(n1457), .Y(n592) );
  INVX1 U935 ( .A(n1466), .Y(n871) );
  INVX1 U936 ( .A(n1467), .Y(n872) );
  INVX1 U937 ( .A(n1468), .Y(n873) );
  INVX1 U938 ( .A(n1477), .Y(n874) );
  INVX1 U939 ( .A(n1478), .Y(n875) );
  INVX1 U940 ( .A(n1479), .Y(n876) );
  AND2X2 U941 ( .A(n1332), .B(n1331), .Y(n877) );
  INVX1 U942 ( .A(n877), .Y(n878) );
  AND2X2 U943 ( .A(n1345), .B(n1344), .Y(n879) );
  INVX1 U944 ( .A(n879), .Y(n880) );
  AND2X2 U945 ( .A(n1358), .B(n1357), .Y(n881) );
  INVX1 U946 ( .A(n881), .Y(n882) );
  AND2X2 U947 ( .A(n1371), .B(n1370), .Y(n883) );
  INVX1 U948 ( .A(n883), .Y(n884) );
  AND2X2 U949 ( .A(n1384), .B(n1383), .Y(n885) );
  INVX1 U950 ( .A(n885), .Y(n886) );
  AND2X2 U951 ( .A(n1397), .B(n1396), .Y(n887) );
  INVX1 U952 ( .A(n887), .Y(n888) );
  AND2X2 U953 ( .A(n1487), .B(n1486), .Y(n889) );
  INVX1 U954 ( .A(n889), .Y(n890) );
  AND2X2 U955 ( .A(n1500), .B(n1499), .Y(n891) );
  INVX1 U956 ( .A(n891), .Y(n892) );
  INVX1 U957 ( .A(n1325), .Y(n893) );
  INVX1 U958 ( .A(n1326), .Y(n894) );
  INVX1 U959 ( .A(n1327), .Y(n895) );
  INVX1 U960 ( .A(n1416), .Y(n896) );
  INVX1 U961 ( .A(n1417), .Y(n897) );
  INVX1 U962 ( .A(n1418), .Y(n898) );
  INVX1 U963 ( .A(n1427), .Y(n899) );
  INVX1 U964 ( .A(n1428), .Y(n900) );
  INVX1 U965 ( .A(n1429), .Y(n901) );
  INVX1 U966 ( .A(n1438), .Y(n902) );
  INVX1 U967 ( .A(n1439), .Y(n903) );
  INVX1 U968 ( .A(n1440), .Y(n904) );
  INVX1 U969 ( .A(n1449), .Y(n905) );
  INVX1 U970 ( .A(n1450), .Y(n906) );
  INVX1 U971 ( .A(n1451), .Y(n907) );
  INVX1 U972 ( .A(n1460), .Y(n908) );
  INVX1 U973 ( .A(n1461), .Y(n909) );
  INVX1 U974 ( .A(n1462), .Y(n910) );
  INVX1 U975 ( .A(n1471), .Y(n911) );
  INVX1 U976 ( .A(n1472), .Y(n912) );
  INVX1 U977 ( .A(n1473), .Y(n913) );
  INVX1 U978 ( .A(n1482), .Y(n914) );
  INVX1 U979 ( .A(n1483), .Y(n915) );
  INVX1 U980 ( .A(n1484), .Y(n916) );
  AND2X2 U981 ( .A(n1334), .B(n1333), .Y(n917) );
  INVX1 U982 ( .A(n917), .Y(n918) );
  AND2X2 U983 ( .A(n1347), .B(n1346), .Y(n919) );
  INVX1 U984 ( .A(n919), .Y(n920) );
  AND2X2 U985 ( .A(n1360), .B(n1359), .Y(n921) );
  INVX1 U986 ( .A(n921), .Y(n922) );
  AND2X2 U987 ( .A(n1373), .B(n1372), .Y(n923) );
  INVX1 U988 ( .A(n923), .Y(n924) );
  AND2X2 U989 ( .A(n1386), .B(n1385), .Y(n925) );
  INVX1 U990 ( .A(n925), .Y(n926) );
  AND2X2 U991 ( .A(n1399), .B(n1398), .Y(n927) );
  INVX1 U992 ( .A(n927), .Y(n928) );
  AND2X2 U993 ( .A(n1489), .B(n1488), .Y(n929) );
  INVX1 U994 ( .A(n929), .Y(n930) );
  AND2X2 U995 ( .A(n1502), .B(n1501), .Y(n931) );
  INVX1 U996 ( .A(n931), .Y(n932) );
  BUFX2 U997 ( .A(n1341), .Y(n933) );
  BUFX2 U998 ( .A(n1354), .Y(n934) );
  BUFX2 U999 ( .A(n1367), .Y(n935) );
  BUFX2 U1000 ( .A(n1380), .Y(n936) );
  BUFX2 U1001 ( .A(n1393), .Y(n937) );
  BUFX2 U1002 ( .A(n1406), .Y(n938) );
  BUFX2 U1003 ( .A(n1496), .Y(n939) );
  INVX1 U1004 ( .A(n970), .Y(n940) );
  INVX1 U1005 ( .A(n1503), .Y(n941) );
  INVX1 U1006 ( .A(n1504), .Y(n942) );
  BUFX2 U1007 ( .A(n1556), .Y(n970) );
  BUFX2 U1008 ( .A(n1339), .Y(n943) );
  BUFX2 U1009 ( .A(n1352), .Y(n944) );
  BUFX2 U1010 ( .A(n1365), .Y(n945) );
  BUFX2 U1011 ( .A(n1378), .Y(n946) );
  BUFX2 U1012 ( .A(n1391), .Y(n947) );
  BUFX2 U1013 ( .A(n1404), .Y(n948) );
  BUFX2 U1014 ( .A(n1494), .Y(n949) );
  INVX1 U1015 ( .A(n971), .Y(n950) );
  INVX1 U1016 ( .A(n1505), .Y(n951) );
  INVX1 U1017 ( .A(n1506), .Y(n952) );
  BUFX2 U1018 ( .A(n1518), .Y(n971) );
  BUFX2 U1019 ( .A(n1842), .Y(err) );
  BUFX2 U1020 ( .A(n1527), .Y(n972) );
  BUFX2 U1021 ( .A(n1545), .Y(n974) );
  BUFX2 U1022 ( .A(n1555), .Y(n975) );
  BUFX2 U1023 ( .A(n1565), .Y(n976) );
  BUFX2 U1024 ( .A(n1575), .Y(n977) );
  BUFX2 U1025 ( .A(n1584), .Y(n978) );
  BUFX2 U1026 ( .A(n1594), .Y(n979) );
  BUFX2 U1027 ( .A(n1614), .Y(n982) );
  BUFX2 U1028 ( .A(n1633), .Y(n985) );
  BUFX2 U1029 ( .A(n1654), .Y(n988) );
  BUFX2 U1030 ( .A(n1674), .Y(n991) );
  BUFX2 U1031 ( .A(n1683), .Y(n992) );
  BUFX2 U1032 ( .A(n1693), .Y(n993) );
  BUFX2 U1033 ( .A(n1702), .Y(n994) );
  BUFX2 U1034 ( .A(n1712), .Y(n995) );
  BUFX2 U1035 ( .A(n1721), .Y(n996) );
  BUFX2 U1036 ( .A(n1731), .Y(n997) );
  BUFX2 U1037 ( .A(n1740), .Y(n998) );
  BUFX2 U1038 ( .A(n1750), .Y(n999) );
  BUFX2 U1039 ( .A(n1769), .Y(n1002) );
  BUFX2 U1040 ( .A(n1789), .Y(n1005) );
  BUFX2 U1041 ( .A(n1809), .Y(n1008) );
  BUFX2 U1042 ( .A(n1822), .Y(n973) );
  AND2X1 U1043 ( .A(n1634), .B(n1322), .Y(n1821) );
  BUFX2 U1044 ( .A(n1841), .Y(n1011) );
  BUFX2 U1045 ( .A(n1604), .Y(n954) );
  BUFX2 U1046 ( .A(n1623), .Y(n955) );
  BUFX2 U1047 ( .A(n1644), .Y(n956) );
  BUFX2 U1048 ( .A(n1664), .Y(n957) );
  BUFX2 U1049 ( .A(n1759), .Y(n958) );
  BUFX2 U1050 ( .A(n1779), .Y(n959) );
  BUFX2 U1051 ( .A(n1799), .Y(n960) );
  BUFX2 U1052 ( .A(n1820), .Y(n961) );
  AND2X1 U1053 ( .A(enable), .B(n1017), .Y(n962) );
  INVX1 U1054 ( .A(n962), .Y(n963) );
  AND2X1 U1055 ( .A(n1517), .B(n1516), .Y(n964) );
  INVX1 U1056 ( .A(n964), .Y(n965) );
  INVX1 U1057 ( .A(n966), .Y(n967) );
  INVX1 U1058 ( .A(n968), .Y(n969) );
  AND2X1 U1059 ( .A(n950), .B(n1314), .Y(n1528) );
  INVX1 U1060 ( .A(rd), .Y(n1026) );
  INVX1 U1061 ( .A(wr), .Y(n1027) );
endmodule


module final_memory_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1842, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1050), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1051), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1052), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1053), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1054), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1055), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1056), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1057), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1058), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1059), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1060), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1061), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1062), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1063), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1064), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1065), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1066), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1067), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1068), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1069), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1070), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1071), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1072), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1073), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1074), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1075), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1076), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1077), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1078), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1079), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1080), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1081), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1082), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1083), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1084), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1085), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1087), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1088), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1089), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1090), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1091), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1092), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1093), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1094), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1095), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1096), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1097), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1098), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1099), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1100), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1101), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1102), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1103), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1104), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1105), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1106), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1107), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1108), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1109), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1110), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1111), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1112), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1113), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1114), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1115), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1116), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1117), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1118), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1119), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1120), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1121), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1122), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1123), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1124), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1125), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1126), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1127), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1128), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1129), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1130), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1131), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1132), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1133), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1134), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1135), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1136), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1137), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1138), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1139), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1140), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1141), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1142), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1143), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1144), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1145), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1146), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1147), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1148), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1149), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1150), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1151), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1152), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1153), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1154), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1155), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1156), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1157), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1158), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1159), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1160), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1161), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1162), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1163), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1164), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1165), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1166), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1167), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1168), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1169), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1170), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1171), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1172), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1173), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1174), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1175), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1176), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1177), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1178), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1179), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1180), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1181), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1182), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1183), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1184), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1185), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1186), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1187), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1188), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1189), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1190), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1191), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1192), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1193), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1194), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1195), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1196), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1197), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1198), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1199), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1200), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1201), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1202), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1203), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1204), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1205), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1206), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1207), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1208), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1209), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1210), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1211), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1212), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1213), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1214), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1215), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1216), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1217), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1218), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1219), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1220), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1221), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1222), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1223), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1224), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1225), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1226), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1227), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1228), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1229), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1230), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1231), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1232), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1233), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1234), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1235), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1236), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1237), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1238), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1239), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1240), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1241), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1242), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1243), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1244), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1245), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1246), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1247), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1248), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1249), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1250), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1251), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1252), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1253), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1254), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1255), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1256), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1257), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1258), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1259), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1260), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1261), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1262), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1263), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1264), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1265), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1266), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1267), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1268), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1269), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1270), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1271), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1272), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1273), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1274), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1275), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1276), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1277), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1278), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1279), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1280), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1281), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1282), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1283), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1284), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1285), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1286), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1287), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1288), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1289), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1290), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1291), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1292), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1293), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1294), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1296), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1297), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1298), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1299), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1300), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1301), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1302), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1303), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1304), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1305), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1306), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1307), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1308), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1309), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1310), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1311), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1312), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1313), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1481), .B(n1480), .Y(n1482) );
  AND2X2 U10 ( .A(n1476), .B(n1475), .Y(n1477) );
  AND2X2 U11 ( .A(n1470), .B(n1469), .Y(n1471) );
  AND2X2 U12 ( .A(n1465), .B(n1464), .Y(n1466) );
  AND2X2 U13 ( .A(n1459), .B(n1458), .Y(n1460) );
  AND2X2 U14 ( .A(n1454), .B(n1453), .Y(n1455) );
  AND2X2 U15 ( .A(n1448), .B(n1447), .Y(n1449) );
  AND2X2 U16 ( .A(n1443), .B(n1442), .Y(n1444) );
  AND2X2 U17 ( .A(n1437), .B(n1436), .Y(n1438) );
  AND2X2 U18 ( .A(n1432), .B(n1431), .Y(n1433) );
  AND2X2 U19 ( .A(n1426), .B(n1425), .Y(n1427) );
  AND2X2 U20 ( .A(n1421), .B(n1420), .Y(n1422) );
  AND2X2 U21 ( .A(n1415), .B(n1414), .Y(n1416) );
  AND2X2 U22 ( .A(n1410), .B(n1409), .Y(n1411) );
  AND2X2 U30 ( .A(n1330), .B(n1030), .Y(n1635) );
  AND2X2 U31 ( .A(n1329), .B(n1030), .Y(n1790) );
  AND2X2 U32 ( .A(n1330), .B(\addr_1c<0> ), .Y(n1655) );
  AND2X2 U33 ( .A(n1329), .B(\addr_1c<0> ), .Y(n1810) );
  AND2X2 U34 ( .A(n1324), .B(n1323), .Y(n1325) );
  AND2X2 U45 ( .A(n1317), .B(n1316), .Y(n1318) );
  NOR3X1 U94 ( .A(n1027), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1026), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1042), .C(n1840), .Y(n1313) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1840) );
  OAI21X1 U98 ( .A(n1011), .B(n1043), .C(n1839), .Y(n1312) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1839) );
  OAI21X1 U100 ( .A(n1011), .B(n1044), .C(n1838), .Y(n1311) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1838) );
  OAI21X1 U102 ( .A(n1011), .B(n1045), .C(n1837), .Y(n1310) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1837) );
  OAI21X1 U104 ( .A(n1011), .B(n1046), .C(n1836), .Y(n1309) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1836) );
  OAI21X1 U106 ( .A(n1011), .B(n1047), .C(n1835), .Y(n1308) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1835) );
  OAI21X1 U108 ( .A(n1011), .B(n1048), .C(n1834), .Y(n1307) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1834) );
  OAI21X1 U110 ( .A(n1011), .B(n1049), .C(n1833), .Y(n1306) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1833) );
  NAND3X1 U112 ( .A(n1832), .B(n1831), .C(n964), .Y(n1841) );
  OAI21X1 U113 ( .A(n6), .B(n1034), .C(n1830), .Y(n1305) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1830) );
  OAI21X1 U115 ( .A(n6), .B(n1035), .C(n1829), .Y(n1304) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1829) );
  OAI21X1 U117 ( .A(n6), .B(n1036), .C(n1828), .Y(n1303) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1828) );
  OAI21X1 U119 ( .A(n6), .B(n1037), .C(n1827), .Y(n1302) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1827) );
  OAI21X1 U121 ( .A(n6), .B(n1038), .C(n1826), .Y(n1301) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1826) );
  OAI21X1 U123 ( .A(n6), .B(n1039), .C(n1825), .Y(n1300) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1825) );
  OAI21X1 U125 ( .A(n6), .B(n1040), .C(n1824), .Y(n1299) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1824) );
  OAI21X1 U127 ( .A(n6), .B(n1041), .C(n1823), .Y(n1298) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1823) );
  OAI21X1 U130 ( .A(n1042), .B(n1010), .C(n1819), .Y(n1297) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1819) );
  OAI21X1 U132 ( .A(n1043), .B(n1009), .C(n1818), .Y(n1296) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1818) );
  OAI21X1 U134 ( .A(n1044), .B(n1009), .C(n1817), .Y(n1295) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1817) );
  OAI21X1 U136 ( .A(n1045), .B(n1009), .C(n1816), .Y(n1294) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1816) );
  OAI21X1 U138 ( .A(n1046), .B(n1009), .C(n1815), .Y(n1293) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1815) );
  OAI21X1 U140 ( .A(n1047), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1814) );
  OAI21X1 U142 ( .A(n1048), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1813) );
  OAI21X1 U144 ( .A(n1049), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1812) );
  NAND3X1 U146 ( .A(n1811), .B(n1832), .C(n1810), .Y(n1820) );
  OAI21X1 U147 ( .A(n1034), .B(n1008), .C(n1808), .Y(n1289) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1808) );
  OAI21X1 U149 ( .A(n1035), .B(n1008), .C(n1807), .Y(n1288) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1807) );
  OAI21X1 U151 ( .A(n1036), .B(n1008), .C(n1806), .Y(n1287) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1806) );
  OAI21X1 U153 ( .A(n1037), .B(n1008), .C(n1805), .Y(n1286) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1805) );
  OAI21X1 U155 ( .A(n1038), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1804) );
  OAI21X1 U157 ( .A(n1039), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1803) );
  OAI21X1 U159 ( .A(n1040), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1802) );
  OAI21X1 U161 ( .A(n1041), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1801) );
  NAND3X1 U163 ( .A(n973), .B(n1832), .C(n1800), .Y(n1809) );
  OAI21X1 U164 ( .A(n1042), .B(n1007), .C(n1798), .Y(n1281) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1798) );
  OAI21X1 U166 ( .A(n1043), .B(n1006), .C(n1797), .Y(n1280) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1797) );
  OAI21X1 U168 ( .A(n1044), .B(n1006), .C(n1796), .Y(n1279) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1796) );
  OAI21X1 U170 ( .A(n1045), .B(n1006), .C(n1795), .Y(n1278) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1795) );
  OAI21X1 U172 ( .A(n1046), .B(n1006), .C(n1794), .Y(n1277) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1794) );
  OAI21X1 U174 ( .A(n1047), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1793) );
  OAI21X1 U176 ( .A(n1048), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1792) );
  OAI21X1 U178 ( .A(n1049), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1791) );
  NAND3X1 U180 ( .A(n1811), .B(n1832), .C(n1790), .Y(n1799) );
  OAI21X1 U181 ( .A(n1034), .B(n1005), .C(n1788), .Y(n1273) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1788) );
  OAI21X1 U183 ( .A(n1035), .B(n1005), .C(n1787), .Y(n1272) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1787) );
  OAI21X1 U185 ( .A(n1036), .B(n1005), .C(n1786), .Y(n1271) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1786) );
  OAI21X1 U187 ( .A(n1037), .B(n1005), .C(n1785), .Y(n1270) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1785) );
  OAI21X1 U189 ( .A(n1038), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1784) );
  OAI21X1 U191 ( .A(n1039), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1783) );
  OAI21X1 U193 ( .A(n1040), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1782) );
  OAI21X1 U195 ( .A(n1041), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1781) );
  NAND3X1 U197 ( .A(n973), .B(n1832), .C(n1780), .Y(n1789) );
  OAI21X1 U198 ( .A(n1042), .B(n1004), .C(n1778), .Y(n1265) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1778) );
  OAI21X1 U200 ( .A(n1043), .B(n1003), .C(n1777), .Y(n1264) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1777) );
  OAI21X1 U202 ( .A(n1044), .B(n1003), .C(n1776), .Y(n1263) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1776) );
  OAI21X1 U204 ( .A(n1045), .B(n1003), .C(n1775), .Y(n1262) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1775) );
  OAI21X1 U206 ( .A(n1046), .B(n1003), .C(n1774), .Y(n1261) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1774) );
  OAI21X1 U208 ( .A(n1047), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1773) );
  OAI21X1 U210 ( .A(n1048), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1772) );
  OAI21X1 U212 ( .A(n1049), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1771) );
  NAND3X1 U214 ( .A(n1810), .B(n1013), .C(n1770), .Y(n1779) );
  OAI21X1 U215 ( .A(n1034), .B(n1002), .C(n1768), .Y(n1257) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1768) );
  OAI21X1 U217 ( .A(n1035), .B(n1002), .C(n1767), .Y(n1256) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1767) );
  OAI21X1 U219 ( .A(n1036), .B(n1002), .C(n1766), .Y(n1255) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1766) );
  OAI21X1 U221 ( .A(n1037), .B(n1002), .C(n1765), .Y(n1254) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1765) );
  OAI21X1 U223 ( .A(n1038), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1764) );
  OAI21X1 U225 ( .A(n1039), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1763) );
  OAI21X1 U227 ( .A(n1040), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1762) );
  OAI21X1 U229 ( .A(n1041), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1761) );
  NAND3X1 U231 ( .A(n973), .B(n1013), .C(n1760), .Y(n1769) );
  OAI21X1 U232 ( .A(n1042), .B(n1001), .C(n1758), .Y(n1249) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1758) );
  OAI21X1 U234 ( .A(n1043), .B(n1000), .C(n1757), .Y(n1248) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1757) );
  OAI21X1 U236 ( .A(n1044), .B(n1000), .C(n1756), .Y(n1247) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1756) );
  OAI21X1 U238 ( .A(n1045), .B(n1000), .C(n1755), .Y(n1246) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1755) );
  OAI21X1 U240 ( .A(n1046), .B(n1000), .C(n1754), .Y(n1245) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1754) );
  OAI21X1 U242 ( .A(n1047), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1753) );
  OAI21X1 U244 ( .A(n1048), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1752) );
  OAI21X1 U246 ( .A(n1049), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1751) );
  NAND3X1 U248 ( .A(n1790), .B(n1013), .C(n1770), .Y(n1759) );
  OAI21X1 U249 ( .A(n1034), .B(n999), .C(n1749), .Y(n1241) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1749) );
  OAI21X1 U251 ( .A(n1035), .B(n999), .C(n1748), .Y(n1240) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1748) );
  OAI21X1 U253 ( .A(n1036), .B(n999), .C(n1747), .Y(n1239) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1747) );
  OAI21X1 U255 ( .A(n1037), .B(n999), .C(n1746), .Y(n1238) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1746) );
  OAI21X1 U257 ( .A(n1038), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1745) );
  OAI21X1 U259 ( .A(n1039), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1744) );
  OAI21X1 U261 ( .A(n1040), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1743) );
  OAI21X1 U263 ( .A(n1041), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1742) );
  NAND3X1 U265 ( .A(n973), .B(n1013), .C(n1741), .Y(n1750) );
  OAI21X1 U266 ( .A(n1042), .B(n998), .C(n1739), .Y(n1233) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1739) );
  OAI21X1 U268 ( .A(n1043), .B(n998), .C(n1738), .Y(n1232) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1738) );
  OAI21X1 U270 ( .A(n1044), .B(n998), .C(n1737), .Y(n1231) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1737) );
  OAI21X1 U272 ( .A(n1045), .B(n998), .C(n1736), .Y(n1230) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1736) );
  OAI21X1 U274 ( .A(n1046), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1735) );
  OAI21X1 U276 ( .A(n1047), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1734) );
  OAI21X1 U278 ( .A(n1048), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1733) );
  OAI21X1 U280 ( .A(n1049), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1732) );
  NAND3X1 U282 ( .A(n1810), .B(n1013), .C(n969), .Y(n1740) );
  OAI21X1 U283 ( .A(n1034), .B(n997), .C(n1730), .Y(n1225) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1730) );
  OAI21X1 U285 ( .A(n1035), .B(n997), .C(n1729), .Y(n1224) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1729) );
  OAI21X1 U287 ( .A(n1036), .B(n997), .C(n1728), .Y(n1223) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1728) );
  OAI21X1 U289 ( .A(n1037), .B(n997), .C(n1727), .Y(n1222) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1727) );
  OAI21X1 U291 ( .A(n1038), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1726) );
  OAI21X1 U293 ( .A(n1039), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1725) );
  OAI21X1 U295 ( .A(n1040), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1724) );
  OAI21X1 U297 ( .A(n1041), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1723) );
  NAND3X1 U299 ( .A(n973), .B(n1013), .C(n1722), .Y(n1731) );
  OAI21X1 U300 ( .A(n1042), .B(n996), .C(n1720), .Y(n1217) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1720) );
  OAI21X1 U302 ( .A(n1043), .B(n996), .C(n1719), .Y(n1216) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1719) );
  OAI21X1 U304 ( .A(n1044), .B(n996), .C(n1718), .Y(n1215) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1718) );
  OAI21X1 U306 ( .A(n1045), .B(n996), .C(n1717), .Y(n1214) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1717) );
  OAI21X1 U308 ( .A(n1046), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1716) );
  OAI21X1 U310 ( .A(n1047), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1715) );
  OAI21X1 U312 ( .A(n1048), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1714) );
  OAI21X1 U314 ( .A(n1049), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1713) );
  NAND3X1 U316 ( .A(n1790), .B(n1013), .C(n969), .Y(n1721) );
  OAI21X1 U317 ( .A(n1034), .B(n995), .C(n1711), .Y(n1209) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1711) );
  OAI21X1 U319 ( .A(n1035), .B(n995), .C(n1710), .Y(n1208) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1710) );
  OAI21X1 U321 ( .A(n1036), .B(n995), .C(n1709), .Y(n1207) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1709) );
  OAI21X1 U323 ( .A(n1037), .B(n995), .C(n1708), .Y(n1206) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1708) );
  OAI21X1 U325 ( .A(n1038), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1707) );
  OAI21X1 U327 ( .A(n1039), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1706) );
  OAI21X1 U329 ( .A(n1040), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1705) );
  OAI21X1 U331 ( .A(n1041), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1704) );
  NAND3X1 U333 ( .A(n973), .B(n1013), .C(n1703), .Y(n1712) );
  OAI21X1 U334 ( .A(n1042), .B(n994), .C(n1701), .Y(n1201) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1701) );
  OAI21X1 U336 ( .A(n1043), .B(n994), .C(n1700), .Y(n1200) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1700) );
  OAI21X1 U338 ( .A(n1044), .B(n994), .C(n1699), .Y(n1199) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1699) );
  OAI21X1 U340 ( .A(n1045), .B(n994), .C(n1698), .Y(n1198) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1698) );
  OAI21X1 U342 ( .A(n1046), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1697) );
  OAI21X1 U344 ( .A(n1047), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1696) );
  OAI21X1 U346 ( .A(n1048), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1695) );
  OAI21X1 U348 ( .A(n1049), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1694) );
  NAND3X1 U350 ( .A(n1810), .B(n1013), .C(n967), .Y(n1702) );
  OAI21X1 U351 ( .A(n1034), .B(n993), .C(n1692), .Y(n1193) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1692) );
  OAI21X1 U353 ( .A(n1035), .B(n993), .C(n1691), .Y(n1192) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1691) );
  OAI21X1 U355 ( .A(n1036), .B(n993), .C(n1690), .Y(n1191) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1690) );
  OAI21X1 U357 ( .A(n1037), .B(n993), .C(n1689), .Y(n1190) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1689) );
  OAI21X1 U359 ( .A(n1038), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1688) );
  OAI21X1 U361 ( .A(n1039), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1687) );
  OAI21X1 U363 ( .A(n1040), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1686) );
  OAI21X1 U365 ( .A(n1041), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1685) );
  NAND3X1 U367 ( .A(n973), .B(n1013), .C(n1684), .Y(n1693) );
  OAI21X1 U368 ( .A(n1042), .B(n992), .C(n1682), .Y(n1185) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1682) );
  OAI21X1 U370 ( .A(n1043), .B(n992), .C(n1681), .Y(n1184) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1681) );
  OAI21X1 U372 ( .A(n1044), .B(n992), .C(n1680), .Y(n1183) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1680) );
  OAI21X1 U374 ( .A(n1045), .B(n992), .C(n1679), .Y(n1182) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1679) );
  OAI21X1 U376 ( .A(n1046), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1678) );
  OAI21X1 U378 ( .A(n1047), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1677) );
  OAI21X1 U380 ( .A(n1048), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1676) );
  OAI21X1 U382 ( .A(n1049), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1675) );
  NAND3X1 U384 ( .A(n1790), .B(n1013), .C(n967), .Y(n1683) );
  OAI21X1 U385 ( .A(n1034), .B(n991), .C(n1673), .Y(n1177) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1673) );
  OAI21X1 U387 ( .A(n1035), .B(n991), .C(n1672), .Y(n1176) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1672) );
  OAI21X1 U389 ( .A(n1036), .B(n991), .C(n1671), .Y(n1175) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1671) );
  OAI21X1 U391 ( .A(n1037), .B(n991), .C(n1670), .Y(n1174) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1670) );
  OAI21X1 U393 ( .A(n1038), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1669) );
  OAI21X1 U395 ( .A(n1039), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1668) );
  OAI21X1 U397 ( .A(n1040), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1667) );
  OAI21X1 U399 ( .A(n1041), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1666) );
  NAND3X1 U401 ( .A(n973), .B(n1013), .C(n1665), .Y(n1674) );
  OAI21X1 U402 ( .A(n1042), .B(n990), .C(n1663), .Y(n1169) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1663) );
  OAI21X1 U404 ( .A(n1043), .B(n989), .C(n1662), .Y(n1168) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1662) );
  OAI21X1 U406 ( .A(n1044), .B(n989), .C(n1661), .Y(n1167) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1661) );
  OAI21X1 U408 ( .A(n1045), .B(n989), .C(n1660), .Y(n1166) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1660) );
  OAI21X1 U410 ( .A(n1046), .B(n989), .C(n1659), .Y(n1165) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1659) );
  OAI21X1 U412 ( .A(n1047), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1658) );
  OAI21X1 U414 ( .A(n1048), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1657) );
  OAI21X1 U416 ( .A(n1049), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1656) );
  NAND3X1 U418 ( .A(n1811), .B(n1012), .C(n1655), .Y(n1664) );
  OAI21X1 U419 ( .A(n1034), .B(n988), .C(n1653), .Y(n1161) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1653) );
  OAI21X1 U421 ( .A(n1035), .B(n988), .C(n1652), .Y(n1160) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1652) );
  OAI21X1 U423 ( .A(n1036), .B(n988), .C(n1651), .Y(n1159) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1651) );
  OAI21X1 U425 ( .A(n1037), .B(n988), .C(n1650), .Y(n1158) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1650) );
  OAI21X1 U427 ( .A(n1038), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1649) );
  OAI21X1 U429 ( .A(n1039), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1648) );
  OAI21X1 U431 ( .A(n1040), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1647) );
  OAI21X1 U433 ( .A(n1041), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1646) );
  NAND3X1 U435 ( .A(n973), .B(n1012), .C(n1645), .Y(n1654) );
  OAI21X1 U436 ( .A(n1042), .B(n987), .C(n1643), .Y(n1153) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1643) );
  OAI21X1 U438 ( .A(n1043), .B(n986), .C(n1642), .Y(n1152) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1642) );
  OAI21X1 U440 ( .A(n1044), .B(n986), .C(n1641), .Y(n1151) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1641) );
  OAI21X1 U442 ( .A(n1045), .B(n986), .C(n1640), .Y(n1150) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1640) );
  OAI21X1 U444 ( .A(n1046), .B(n986), .C(n1639), .Y(n1149) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1639) );
  OAI21X1 U446 ( .A(n1047), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1638) );
  OAI21X1 U448 ( .A(n1048), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1637) );
  OAI21X1 U450 ( .A(n1049), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1636) );
  NAND3X1 U452 ( .A(n1811), .B(n1012), .C(n1635), .Y(n1644) );
  OAI21X1 U453 ( .A(n1034), .B(n985), .C(n1632), .Y(n1145) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1632) );
  OAI21X1 U455 ( .A(n1035), .B(n985), .C(n1631), .Y(n1144) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1631) );
  OAI21X1 U457 ( .A(n1036), .B(n985), .C(n1630), .Y(n1143) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1630) );
  OAI21X1 U459 ( .A(n1037), .B(n985), .C(n1629), .Y(n1142) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1629) );
  OAI21X1 U461 ( .A(n1038), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1628) );
  OAI21X1 U463 ( .A(n1039), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1627) );
  OAI21X1 U465 ( .A(n1040), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1626) );
  OAI21X1 U467 ( .A(n1041), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1625) );
  NAND3X1 U469 ( .A(n973), .B(n1012), .C(n1624), .Y(n1633) );
  OAI21X1 U470 ( .A(n1042), .B(n984), .C(n1622), .Y(n1137) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1622) );
  OAI21X1 U472 ( .A(n1043), .B(n983), .C(n1621), .Y(n1136) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1621) );
  OAI21X1 U474 ( .A(n1044), .B(n983), .C(n1620), .Y(n1135) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1620) );
  OAI21X1 U476 ( .A(n1045), .B(n983), .C(n1619), .Y(n1134) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1619) );
  OAI21X1 U478 ( .A(n1046), .B(n983), .C(n1618), .Y(n1133) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1618) );
  OAI21X1 U480 ( .A(n1047), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1617) );
  OAI21X1 U482 ( .A(n1048), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1616) );
  OAI21X1 U484 ( .A(n1049), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1615) );
  NAND3X1 U486 ( .A(n1770), .B(n1012), .C(n1655), .Y(n1623) );
  OAI21X1 U487 ( .A(n1034), .B(n982), .C(n1613), .Y(n1129) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1613) );
  OAI21X1 U489 ( .A(n1035), .B(n982), .C(n1612), .Y(n1128) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1612) );
  OAI21X1 U491 ( .A(n1036), .B(n982), .C(n1611), .Y(n1127) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1611) );
  OAI21X1 U493 ( .A(n1037), .B(n982), .C(n1610), .Y(n1126) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1610) );
  OAI21X1 U495 ( .A(n1038), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1609) );
  OAI21X1 U497 ( .A(n1039), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1608) );
  OAI21X1 U499 ( .A(n1040), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1607) );
  OAI21X1 U501 ( .A(n1041), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1606) );
  NAND3X1 U503 ( .A(n973), .B(n1012), .C(n1605), .Y(n1614) );
  OAI21X1 U504 ( .A(n1042), .B(n981), .C(n1603), .Y(n1121) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1603) );
  OAI21X1 U506 ( .A(n1043), .B(n980), .C(n1602), .Y(n1120) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1602) );
  OAI21X1 U508 ( .A(n1044), .B(n980), .C(n1601), .Y(n1119) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1601) );
  OAI21X1 U510 ( .A(n1045), .B(n980), .C(n1600), .Y(n1118) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1600) );
  OAI21X1 U512 ( .A(n1046), .B(n980), .C(n1599), .Y(n1117) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1599) );
  OAI21X1 U514 ( .A(n1047), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1598) );
  OAI21X1 U516 ( .A(n1048), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1597) );
  OAI21X1 U518 ( .A(n1049), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1596) );
  NAND3X1 U520 ( .A(n1770), .B(n1012), .C(n1635), .Y(n1604) );
  OAI21X1 U521 ( .A(n1034), .B(n979), .C(n1593), .Y(n1113) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1593) );
  OAI21X1 U523 ( .A(n1035), .B(n979), .C(n1592), .Y(n1112) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1592) );
  OAI21X1 U525 ( .A(n1036), .B(n979), .C(n1591), .Y(n1111) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1591) );
  OAI21X1 U527 ( .A(n1037), .B(n979), .C(n1590), .Y(n1110) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1590) );
  OAI21X1 U529 ( .A(n1038), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1589) );
  OAI21X1 U531 ( .A(n1039), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1588) );
  OAI21X1 U533 ( .A(n1040), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1587) );
  OAI21X1 U535 ( .A(n1041), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1586) );
  NAND3X1 U537 ( .A(n973), .B(n1012), .C(n1585), .Y(n1594) );
  OAI21X1 U538 ( .A(n1042), .B(n978), .C(n1583), .Y(n1105) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1583) );
  OAI21X1 U540 ( .A(n1043), .B(n978), .C(n1582), .Y(n1104) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1582) );
  OAI21X1 U542 ( .A(n1044), .B(n978), .C(n1581), .Y(n1103) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1581) );
  OAI21X1 U544 ( .A(n1045), .B(n978), .C(n1580), .Y(n1102) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1580) );
  OAI21X1 U546 ( .A(n1046), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1579) );
  OAI21X1 U548 ( .A(n1047), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1578) );
  OAI21X1 U550 ( .A(n1048), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1577) );
  OAI21X1 U552 ( .A(n1049), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1576) );
  NAND3X1 U554 ( .A(n969), .B(n1012), .C(n1655), .Y(n1584) );
  OAI21X1 U555 ( .A(n1034), .B(n977), .C(n1574), .Y(n1097) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1574) );
  OAI21X1 U557 ( .A(n1035), .B(n977), .C(n1573), .Y(n1096) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1573) );
  OAI21X1 U559 ( .A(n1036), .B(n977), .C(n1572), .Y(n1095) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1572) );
  OAI21X1 U561 ( .A(n1037), .B(n977), .C(n1571), .Y(n1094) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1571) );
  OAI21X1 U563 ( .A(n1038), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1570) );
  OAI21X1 U565 ( .A(n1039), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1569) );
  OAI21X1 U567 ( .A(n1040), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1568) );
  OAI21X1 U569 ( .A(n1041), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1567) );
  NAND3X1 U571 ( .A(n973), .B(n1012), .C(n1566), .Y(n1575) );
  OAI21X1 U572 ( .A(n1042), .B(n976), .C(n1564), .Y(n1089) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1564) );
  OAI21X1 U574 ( .A(n1043), .B(n976), .C(n1563), .Y(n1088) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1563) );
  OAI21X1 U576 ( .A(n1044), .B(n976), .C(n1562), .Y(n1087) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1562) );
  OAI21X1 U578 ( .A(n1045), .B(n976), .C(n1561), .Y(n1086) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1561) );
  OAI21X1 U580 ( .A(n1046), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1560) );
  OAI21X1 U582 ( .A(n1047), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1559) );
  OAI21X1 U584 ( .A(n1048), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1558) );
  OAI21X1 U586 ( .A(n1049), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1557) );
  NAND3X1 U588 ( .A(n969), .B(n1012), .C(n1635), .Y(n1565) );
  OAI21X1 U590 ( .A(n1034), .B(n975), .C(n1554), .Y(n1081) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1554) );
  OAI21X1 U592 ( .A(n1035), .B(n975), .C(n1553), .Y(n1080) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1553) );
  OAI21X1 U594 ( .A(n1036), .B(n975), .C(n1552), .Y(n1079) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1552) );
  OAI21X1 U596 ( .A(n1037), .B(n975), .C(n1551), .Y(n1078) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1551) );
  OAI21X1 U598 ( .A(n1038), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1550) );
  OAI21X1 U600 ( .A(n1039), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1549) );
  OAI21X1 U602 ( .A(n1040), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1548) );
  OAI21X1 U604 ( .A(n1041), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1547) );
  NAND3X1 U606 ( .A(n973), .B(n1012), .C(n1546), .Y(n1555) );
  OAI21X1 U607 ( .A(n1042), .B(n974), .C(n1544), .Y(n1073) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1544) );
  OAI21X1 U609 ( .A(n1043), .B(n974), .C(n1543), .Y(n1072) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1543) );
  OAI21X1 U611 ( .A(n1044), .B(n974), .C(n1542), .Y(n1071) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1542) );
  OAI21X1 U613 ( .A(n1045), .B(n974), .C(n1541), .Y(n1070) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1541) );
  OAI21X1 U615 ( .A(n1046), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1540) );
  OAI21X1 U617 ( .A(n1047), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1539) );
  OAI21X1 U619 ( .A(n1048), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1538) );
  OAI21X1 U621 ( .A(n1049), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1537) );
  NAND3X1 U623 ( .A(n967), .B(n1012), .C(n1655), .Y(n1545) );
  OAI21X1 U624 ( .A(n1034), .B(n8), .C(n1536), .Y(n1065) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1536) );
  OAI21X1 U626 ( .A(n1035), .B(n8), .C(n1535), .Y(n1064) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1535) );
  OAI21X1 U628 ( .A(n1036), .B(n8), .C(n1534), .Y(n1063) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1534) );
  OAI21X1 U630 ( .A(n1037), .B(n8), .C(n1533), .Y(n1062) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1533) );
  OAI21X1 U632 ( .A(n1038), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1532) );
  OAI21X1 U634 ( .A(n1039), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1531) );
  OAI21X1 U636 ( .A(n1040), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1530) );
  OAI21X1 U638 ( .A(n1041), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1529) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1822) );
  OAI21X1 U642 ( .A(n1042), .B(n972), .C(n1526), .Y(n1057) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1526) );
  OAI21X1 U644 ( .A(n1043), .B(n972), .C(n1525), .Y(n1056) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1525) );
  OAI21X1 U646 ( .A(n1044), .B(n972), .C(n1524), .Y(n1055) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1524) );
  OAI21X1 U648 ( .A(n1045), .B(n972), .C(n1523), .Y(n1054) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1523) );
  OAI21X1 U650 ( .A(n1046), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1522) );
  OAI21X1 U652 ( .A(n1047), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1521) );
  OAI21X1 U654 ( .A(n1048), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1520) );
  OAI21X1 U656 ( .A(n1049), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1519) );
  NAND3X1 U658 ( .A(n967), .B(n1013), .C(n1635), .Y(n1527) );
  NOR3X1 U661 ( .A(n1515), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1516) );
  NOR3X1 U662 ( .A(n1514), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1517) );
  AOI21X1 U663 ( .A(n461), .B(n1513), .C(n963), .Y(n1842) );
  OAI21X1 U665 ( .A(rd), .B(n1512), .C(wr), .Y(n1513) );
  NAND3X1 U667 ( .A(n1511), .B(n1029), .C(n1510), .Y(n1512) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1510) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1511) );
  AOI21X1 U670 ( .A(n448), .B(n1508), .C(n1028), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1507), .C(n4), .Y(n1508) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1790), .C(\mem<0><1> ), .D(n1635), .Y(
        n1505) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1810), .C(\mem<2><1> ), .D(n1655), .Y(
        n1506) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1790), .C(\mem<4><1> ), .D(n1635), .Y(
        n1503) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1810), .C(\mem<6><1> ), .D(n1655), .Y(
        n1504) );
  AOI22X1 U678 ( .A(n1595), .B(n892), .C(n1634), .D(n932), .Y(n1509) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1790), .C(\mem<12><1> ), .D(n1635), .Y(
        n1501) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1810), .C(\mem<14><1> ), .D(n1655), .Y(
        n1502) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1790), .C(\mem<8><1> ), .D(n1635), .Y(
        n1499) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1810), .C(\mem<10><1> ), .D(n1655), .Y(
        n1500) );
  AOI21X1 U685 ( .A(n447), .B(n1497), .C(n1028), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1495), .C(n950), .Y(n1497) );
  AOI21X1 U687 ( .A(n1493), .B(n1492), .C(n971), .Y(n1494) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1790), .C(\mem<0><0> ), .D(n1635), .Y(
        n1492) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1810), .C(\mem<2><0> ), .D(n1655), .Y(
        n1493) );
  AOI21X1 U690 ( .A(n1491), .B(n1490), .C(n970), .Y(n1496) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1790), .C(\mem<4><0> ), .D(n1635), .Y(
        n1490) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1810), .C(\mem<6><0> ), .D(n1655), .Y(
        n1491) );
  AOI22X1 U693 ( .A(n1595), .B(n890), .C(n1634), .D(n930), .Y(n1498) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1790), .C(\mem<12><0> ), .D(n1635), .Y(
        n1488) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1810), .C(\mem<14><0> ), .D(n1655), .Y(
        n1489) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1790), .C(\mem<8><0> ), .D(n1635), .Y(
        n1486) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1810), .C(\mem<10><0> ), .D(n1655), .Y(
        n1487) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1485) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1684), .C(\mem<19><7> ), .D(n1703), .Y(
        n1480) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1722), .C(\mem<23><7> ), .D(n1741), .Y(
        n1481) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1760), .C(\mem<27><7> ), .D(n1780), .Y(
        n1483) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1800), .C(\mem<31><7> ), .D(n1821), .Y(
        n1484) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1528), .C(\mem<3><7> ), .D(n1546), .Y(
        n1475) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1566), .C(\mem<7><7> ), .D(n1585), .Y(
        n1476) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1605), .C(\mem<11><7> ), .D(n1624), .Y(
        n1478) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1645), .C(\mem<15><7> ), .D(n1665), .Y(
        n1479) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1474) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1684), .C(\mem<19><6> ), .D(n1703), .Y(
        n1469) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1722), .C(\mem<23><6> ), .D(n1741), .Y(
        n1470) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1760), .C(\mem<27><6> ), .D(n1780), .Y(
        n1472) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1800), .C(\mem<31><6> ), .D(n1821), .Y(
        n1473) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1528), .C(\mem<3><6> ), .D(n1546), .Y(
        n1464) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1566), .C(\mem<7><6> ), .D(n1585), .Y(
        n1465) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1605), .C(\mem<11><6> ), .D(n1624), .Y(
        n1467) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1645), .C(\mem<15><6> ), .D(n1665), .Y(
        n1468) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1463) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1684), .C(\mem<19><5> ), .D(n1703), .Y(
        n1458) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1722), .C(\mem<23><5> ), .D(n1741), .Y(
        n1459) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1760), .C(\mem<27><5> ), .D(n1780), .Y(
        n1461) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1800), .C(\mem<31><5> ), .D(n1821), .Y(
        n1462) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1528), .C(\mem<3><5> ), .D(n1546), .Y(
        n1453) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1566), .C(\mem<7><5> ), .D(n1585), .Y(
        n1454) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1605), .C(\mem<11><5> ), .D(n1624), .Y(
        n1456) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1645), .C(\mem<15><5> ), .D(n1665), .Y(
        n1457) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1452) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1684), .C(\mem<19><4> ), .D(n1703), .Y(
        n1447) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1722), .C(\mem<23><4> ), .D(n1741), .Y(
        n1448) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1760), .C(\mem<27><4> ), .D(n1780), .Y(
        n1450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1800), .C(\mem<31><4> ), .D(n1821), .Y(
        n1451) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1528), .C(\mem<3><4> ), .D(n1546), .Y(
        n1442) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1566), .C(\mem<7><4> ), .D(n1585), .Y(
        n1443) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1605), .C(\mem<11><4> ), .D(n1624), .Y(
        n1445) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1645), .C(\mem<15><4> ), .D(n1665), .Y(
        n1446) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1441) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1684), .C(\mem<19><3> ), .D(n1703), .Y(
        n1436) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1722), .C(\mem<23><3> ), .D(n1741), .Y(
        n1437) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1760), .C(\mem<27><3> ), .D(n1780), .Y(
        n1439) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1800), .C(\mem<31><3> ), .D(n1821), .Y(
        n1440) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1528), .C(\mem<3><3> ), .D(n1546), .Y(
        n1431) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1566), .C(\mem<7><3> ), .D(n1585), .Y(
        n1432) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1605), .C(\mem<11><3> ), .D(n1624), .Y(
        n1434) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1645), .C(\mem<15><3> ), .D(n1665), .Y(
        n1435) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1430) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1684), .C(\mem<19><2> ), .D(n1703), .Y(
        n1425) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1722), .C(\mem<23><2> ), .D(n1741), .Y(
        n1426) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1760), .C(\mem<27><2> ), .D(n1780), .Y(
        n1428) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1800), .C(\mem<31><2> ), .D(n1821), .Y(
        n1429) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1528), .C(\mem<3><2> ), .D(n1546), .Y(
        n1420) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1566), .C(\mem<7><2> ), .D(n1585), .Y(
        n1421) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1605), .C(\mem<11><2> ), .D(n1624), .Y(
        n1423) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1645), .C(\mem<15><2> ), .D(n1665), .Y(
        n1424) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1419) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1684), .C(\mem<19><1> ), .D(n1703), .Y(
        n1414) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1722), .C(\mem<23><1> ), .D(n1741), .Y(
        n1415) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1760), .C(\mem<27><1> ), .D(n1780), .Y(
        n1417) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1800), .C(\mem<31><1> ), .D(n1821), .Y(
        n1418) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1528), .C(\mem<3><1> ), .D(n1546), .Y(
        n1409) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1566), .C(\mem<7><1> ), .D(n1585), .Y(
        n1410) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1605), .C(\mem<11><1> ), .D(n1624), .Y(
        n1412) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1645), .C(\mem<15><1> ), .D(n1665), .Y(
        n1413) );
  AOI21X1 U777 ( .A(n435), .B(n1407), .C(n1028), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1405), .C(n949), .Y(n1407) );
  AOI21X1 U779 ( .A(n1403), .B(n1402), .C(n971), .Y(n1404) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1790), .C(\mem<0><7> ), .D(n1635), .Y(
        n1402) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1810), .C(\mem<2><7> ), .D(n1655), .Y(
        n1403) );
  AOI21X1 U782 ( .A(n1401), .B(n1400), .C(n970), .Y(n1406) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1790), .C(\mem<4><7> ), .D(n1635), .Y(
        n1400) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1810), .C(\mem<6><7> ), .D(n1655), .Y(
        n1401) );
  AOI22X1 U785 ( .A(n1595), .B(n888), .C(n1634), .D(n928), .Y(n1408) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1790), .C(\mem<12><7> ), .D(n1635), .Y(
        n1398) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1810), .C(\mem<14><7> ), .D(n1655), .Y(
        n1399) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1790), .C(\mem<8><7> ), .D(n1635), .Y(
        n1396) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1810), .C(\mem<10><7> ), .D(n1655), .Y(
        n1397) );
  AOI21X1 U792 ( .A(n434), .B(n1394), .C(n1028), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1392), .C(n948), .Y(n1394) );
  AOI21X1 U794 ( .A(n1390), .B(n1389), .C(n971), .Y(n1391) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1790), .C(\mem<0><6> ), .D(n1635), .Y(
        n1389) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1810), .C(\mem<2><6> ), .D(n1655), .Y(
        n1390) );
  AOI21X1 U797 ( .A(n1388), .B(n1387), .C(n970), .Y(n1393) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1790), .C(\mem<4><6> ), .D(n1635), .Y(
        n1387) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1810), .C(\mem<6><6> ), .D(n1655), .Y(
        n1388) );
  AOI22X1 U800 ( .A(n1595), .B(n886), .C(n1634), .D(n926), .Y(n1395) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1790), .C(\mem<12><6> ), .D(n1635), .Y(
        n1385) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1810), .C(\mem<14><6> ), .D(n1655), .Y(
        n1386) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1790), .C(\mem<8><6> ), .D(n1635), .Y(
        n1383) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1810), .C(\mem<10><6> ), .D(n1655), .Y(
        n1384) );
  AOI21X1 U807 ( .A(n422), .B(n1381), .C(n1028), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1379), .C(n947), .Y(n1381) );
  AOI21X1 U809 ( .A(n1377), .B(n1376), .C(n971), .Y(n1378) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1790), .C(\mem<0><5> ), .D(n1635), .Y(
        n1376) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1810), .C(\mem<2><5> ), .D(n1655), .Y(
        n1377) );
  AOI21X1 U812 ( .A(n1375), .B(n1374), .C(n970), .Y(n1380) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1790), .C(\mem<4><5> ), .D(n1635), .Y(
        n1374) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1810), .C(\mem<6><5> ), .D(n1655), .Y(
        n1375) );
  AOI22X1 U815 ( .A(n1595), .B(n884), .C(n1634), .D(n924), .Y(n1382) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1790), .C(\mem<12><5> ), .D(n1635), .Y(
        n1372) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1810), .C(\mem<14><5> ), .D(n1655), .Y(
        n1373) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1790), .C(\mem<8><5> ), .D(n1635), .Y(
        n1370) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1810), .C(\mem<10><5> ), .D(n1655), .Y(
        n1371) );
  AOI21X1 U822 ( .A(n421), .B(n1368), .C(n1028), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1366), .C(n946), .Y(n1368) );
  AOI21X1 U824 ( .A(n1364), .B(n1363), .C(n971), .Y(n1365) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1790), .C(\mem<0><4> ), .D(n1635), .Y(
        n1363) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1810), .C(\mem<2><4> ), .D(n1655), .Y(
        n1364) );
  AOI21X1 U827 ( .A(n1362), .B(n1361), .C(n970), .Y(n1367) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1790), .C(\mem<4><4> ), .D(n1635), .Y(
        n1361) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1810), .C(\mem<6><4> ), .D(n1655), .Y(
        n1362) );
  AOI22X1 U830 ( .A(n1595), .B(n882), .C(n1634), .D(n922), .Y(n1369) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1790), .C(\mem<12><4> ), .D(n1635), .Y(
        n1359) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1810), .C(\mem<14><4> ), .D(n1655), .Y(
        n1360) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1790), .C(\mem<8><4> ), .D(n1635), .Y(
        n1357) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1810), .C(\mem<10><4> ), .D(n1655), .Y(
        n1358) );
  AOI21X1 U837 ( .A(n409), .B(n1355), .C(n1028), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1353), .C(n945), .Y(n1355) );
  AOI21X1 U839 ( .A(n1351), .B(n1350), .C(n971), .Y(n1352) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1790), .C(\mem<0><3> ), .D(n1635), .Y(
        n1350) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1810), .C(\mem<2><3> ), .D(n1655), .Y(
        n1351) );
  AOI21X1 U842 ( .A(n1349), .B(n1348), .C(n970), .Y(n1354) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1790), .C(\mem<4><3> ), .D(n1635), .Y(
        n1348) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1810), .C(\mem<6><3> ), .D(n1655), .Y(
        n1349) );
  AOI22X1 U845 ( .A(n1595), .B(n880), .C(n1634), .D(n920), .Y(n1356) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1790), .C(\mem<12><3> ), .D(n1635), .Y(
        n1346) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1810), .C(\mem<14><3> ), .D(n1655), .Y(
        n1347) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1790), .C(\mem<8><3> ), .D(n1635), .Y(
        n1344) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1810), .C(\mem<10><3> ), .D(n1655), .Y(
        n1345) );
  AOI21X1 U852 ( .A(n408), .B(n1342), .C(n1028), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1340), .C(n944), .Y(n1342) );
  AOI21X1 U854 ( .A(n1338), .B(n1337), .C(n971), .Y(n1339) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1790), .C(\mem<0><2> ), .D(n1635), .Y(
        n1337) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1810), .C(\mem<2><2> ), .D(n1655), .Y(
        n1338) );
  AOI21X1 U857 ( .A(n1336), .B(n1335), .C(n970), .Y(n1341) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1790), .C(\mem<4><2> ), .D(n1635), .Y(
        n1335) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1810), .C(\mem<6><2> ), .D(n1655), .Y(
        n1336) );
  AOI22X1 U860 ( .A(n1595), .B(n878), .C(n1634), .D(n918), .Y(n1343) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1790), .C(\mem<12><2> ), .D(n1635), .Y(
        n1333) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1810), .C(\mem<14><2> ), .D(n1655), .Y(
        n1334) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1790), .C(\mem<8><2> ), .D(n1635), .Y(
        n1331) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1810), .C(\mem<10><2> ), .D(n1655), .Y(
        n1332) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1330) );
  NOR2X1 U868 ( .A(n1033), .B(\addr_1c<4> ), .Y(n1329) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1328) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1684), .C(\mem<19><0> ), .D(n1703), .Y(
        n1323) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1722), .C(\mem<23><0> ), .D(n1741), .Y(
        n1324) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1760), .C(\mem<27><0> ), .D(n1780), .Y(
        n1326) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1800), .C(\mem<31><0> ), .D(n1821), .Y(
        n1327) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1528), .C(\mem<3><0> ), .D(n1546), .Y(
        n1316) );
  NAND2X1 U877 ( .A(n1031), .B(n1032), .Y(n1518) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1566), .C(\mem<7><0> ), .D(n1585), .Y(
        n1317) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1032), .Y(n1556) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1605), .C(\mem<11><0> ), .D(n1624), .Y(
        n1319) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1645), .C(\mem<15><0> ), .D(n1665), .Y(
        n1320) );
  dff_50 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1015) );
  dff_49 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1016) );
  dff_48 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1016)
         );
  dff_47 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1016)
         );
  dff_46 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1016)
         );
  dff_45 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1016)
         );
  dff_44 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1016)
         );
  dff_43 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1016)
         );
  dff_42 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1016)
         );
  dff_41 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1016)
         );
  dff_40 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1015)
         );
  dff_39 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1015)
         );
  dff_38 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1015) );
  dff_37 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1015) );
  dff_36 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1015) );
  dff_35 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1015) );
  dff_34 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1015) );
  dff_33 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1015) );
  dff_32 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1015) );
  dff_31 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1015) );
  dff_30 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1015) );
  dff_29 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1015) );
  dff_28 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1015) );
  dff_27 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1015) );
  dff_26 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1015) );
  dff_25 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1015) );
  dff_24 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1015) );
  dff_23 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1015) );
  dff_22 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1015) );
  dff_21 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1015) );
  dff_20 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1015) );
  dff_19 \reg2[0]  ( .q(\data_out<0> ), .d(n1025), .clk(clk), .rst(n1016) );
  dff_18 \reg2[1]  ( .q(\data_out<1> ), .d(n1024), .clk(clk), .rst(n1016) );
  dff_17 \reg2[2]  ( .q(\data_out<2> ), .d(n1023), .clk(clk), .rst(n1016) );
  dff_16 \reg2[3]  ( .q(\data_out<3> ), .d(n1022), .clk(clk), .rst(n1016) );
  dff_15 \reg2[4]  ( .q(\data_out<4> ), .d(n1021), .clk(clk), .rst(n1016) );
  dff_14 \reg2[5]  ( .q(\data_out<5> ), .d(n1020), .clk(clk), .rst(n1016) );
  dff_13 \reg2[6]  ( .q(\data_out<6> ), .d(n1019), .clk(clk), .rst(n1015) );
  dff_12 \reg2[7]  ( .q(\data_out<7> ), .d(n1018), .clk(clk), .rst(n1015) );
  dff_11 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1015) );
  dff_10 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1015) );
  dff_9 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1015) );
  dff_8 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1015) );
  dff_7 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1015) );
  dff_6 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1015) );
  dff_5 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1015) );
  dff_4 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1015) );
  dff_3 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1015) );
  dff_2 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1015) );
  dff_1 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1015) );
  dff_0 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1016) );
  OR2X1 U2 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1514) );
  AND2X1 U3 ( .A(\addr_1c<4> ), .B(n1528), .Y(n1831) );
  INVX1 U4 ( .A(\addr_1c<3> ), .Y(n1033) );
  INVX1 U5 ( .A(\addr_1c<2> ), .Y(n1032) );
  INVX1 U6 ( .A(wr1), .Y(n1029) );
  OR2X1 U7 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1515) );
  INVX1 U8 ( .A(\addr_1c<0> ), .Y(n1030) );
  AND2X1 U23 ( .A(n1030), .B(n1033), .Y(n1314) );
  AND2X1 U24 ( .A(\addr_1c<0> ), .B(n1033), .Y(n1315) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1322) );
  AND2X1 U26 ( .A(\addr_1c<3> ), .B(n1030), .Y(n1321) );
  INVX1 U27 ( .A(\addr_1c<1> ), .Y(n1031) );
  AND2X1 U28 ( .A(n1595), .B(n1322), .Y(n1780) );
  AND2X1 U29 ( .A(n1595), .B(n1321), .Y(n1760) );
  AND2X1 U35 ( .A(n940), .B(n1322), .Y(n1741) );
  AND2X1 U36 ( .A(n940), .B(n1321), .Y(n1722) );
  AND2X1 U37 ( .A(n1322), .B(n951), .Y(n1703) );
  AND2X1 U38 ( .A(n1321), .B(n951), .Y(n1684) );
  AND2X1 U39 ( .A(n1315), .B(n1595), .Y(n1624) );
  AND2X1 U40 ( .A(n1595), .B(n1314), .Y(n1605) );
  AND2X1 U41 ( .A(n1315), .B(n940), .Y(n1585) );
  AND2X1 U42 ( .A(n940), .B(n1314), .Y(n1566) );
  OR2X1 U43 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U44 ( .A(n1315), .B(n951), .Y(n1546) );
  OR2X1 U46 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U47 ( .A(n1634), .B(n1314), .Y(n1645) );
  AND2X1 U48 ( .A(n1315), .B(n1634), .Y(n1665) );
  AND2X1 U49 ( .A(n1321), .B(n1634), .Y(n1800) );
  AND2X1 U50 ( .A(\addr_1c<2> ), .B(n1031), .Y(n1595) );
  AND2X1 U51 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1634) );
  BUFX2 U52 ( .A(n961), .Y(n1010) );
  BUFX2 U53 ( .A(n961), .Y(n1009) );
  BUFX2 U54 ( .A(n960), .Y(n1007) );
  BUFX2 U55 ( .A(n960), .Y(n1006) );
  BUFX2 U56 ( .A(n959), .Y(n1004) );
  BUFX2 U57 ( .A(n959), .Y(n1003) );
  BUFX2 U58 ( .A(n958), .Y(n1001) );
  BUFX2 U59 ( .A(n958), .Y(n1000) );
  BUFX2 U60 ( .A(n957), .Y(n990) );
  BUFX2 U61 ( .A(n957), .Y(n989) );
  BUFX2 U62 ( .A(n956), .Y(n987) );
  BUFX2 U63 ( .A(n956), .Y(n986) );
  BUFX2 U64 ( .A(n955), .Y(n984) );
  BUFX2 U65 ( .A(n955), .Y(n983) );
  BUFX2 U66 ( .A(n954), .Y(n981) );
  BUFX2 U67 ( .A(n954), .Y(n980) );
  INVX1 U68 ( .A(\data_in_1c<0> ), .Y(n1034) );
  INVX1 U69 ( .A(\data_in_1c<1> ), .Y(n1035) );
  INVX1 U70 ( .A(\data_in_1c<2> ), .Y(n1036) );
  INVX1 U71 ( .A(\data_in_1c<3> ), .Y(n1037) );
  INVX1 U72 ( .A(\data_in_1c<4> ), .Y(n1038) );
  INVX1 U73 ( .A(\data_in_1c<5> ), .Y(n1039) );
  INVX1 U74 ( .A(\data_in_1c<6> ), .Y(n1040) );
  INVX1 U75 ( .A(\data_in_1c<7> ), .Y(n1041) );
  INVX1 U76 ( .A(\data_in_1c<8> ), .Y(n1042) );
  INVX1 U77 ( .A(\data_in_1c<9> ), .Y(n1043) );
  INVX1 U78 ( .A(\data_in_1c<10> ), .Y(n1044) );
  INVX1 U79 ( .A(\data_in_1c<11> ), .Y(n1045) );
  INVX1 U80 ( .A(\data_in_1c<12> ), .Y(n1046) );
  INVX1 U81 ( .A(\data_in_1c<13> ), .Y(n1047) );
  INVX1 U82 ( .A(\data_in_1c<14> ), .Y(n1048) );
  INVX1 U83 ( .A(\data_in_1c<15> ), .Y(n1049) );
  AND2X1 U84 ( .A(n1831), .B(\mem<32><0> ), .Y(n1495) );
  AND2X1 U85 ( .A(n1831), .B(\mem<32><1> ), .Y(n1507) );
  AND2X1 U86 ( .A(n1831), .B(\mem<32><2> ), .Y(n1340) );
  AND2X1 U87 ( .A(n1831), .B(\mem<32><3> ), .Y(n1353) );
  AND2X1 U88 ( .A(n1831), .B(\mem<32><4> ), .Y(n1366) );
  AND2X1 U89 ( .A(n1831), .B(\mem<32><5> ), .Y(n1379) );
  AND2X1 U90 ( .A(n1831), .B(\mem<32><6> ), .Y(n1392) );
  AND2X1 U91 ( .A(n1831), .B(\mem<32><7> ), .Y(n1405) );
  INVX1 U92 ( .A(rd1), .Y(n1028) );
  INVX1 U93 ( .A(n1328), .Y(n1025) );
  INVX1 U129 ( .A(n1419), .Y(n1024) );
  INVX1 U589 ( .A(n1430), .Y(n1023) );
  INVX1 U640 ( .A(n1441), .Y(n1022) );
  INVX1 U659 ( .A(n1452), .Y(n1021) );
  INVX1 U660 ( .A(n1463), .Y(n1020) );
  INVX1 U664 ( .A(n1474), .Y(n1019) );
  INVX1 U666 ( .A(n1485), .Y(n1018) );
  INVX2 U672 ( .A(n1017), .Y(n1015) );
  INVX1 U675 ( .A(n1832), .Y(n1014) );
  AND2X1 U679 ( .A(wr1), .B(n1017), .Y(n1832) );
  INVX1 U682 ( .A(rst), .Y(n1017) );
  AND2X1 U694 ( .A(n1634), .B(n964), .Y(n1811) );
  INVX1 U697 ( .A(n1014), .Y(n1012) );
  AND2X1 U701 ( .A(n1595), .B(n964), .Y(n1770) );
  INVX1 U706 ( .A(n1014), .Y(n1013) );
  AND2X1 U712 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U717 ( .A(n1), .Y(n2) );
  AND2X1 U723 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U728 ( .A(n3), .Y(n4) );
  AND2X1 U734 ( .A(n1821), .B(n189), .Y(n5) );
  INVX1 U739 ( .A(n5), .Y(n6) );
  AND2X1 U745 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U750 ( .A(n7), .Y(n8) );
  OR2X1 U756 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U761 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U767 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U772 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U786 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U789 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U801 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U804 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U816 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U819 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U831 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U834 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U846 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U849 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U861 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U864 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U870 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U875 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U882 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U883 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U884 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U885 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U886 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U887 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U888 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U889 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U890 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U891 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U892 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U893 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U894 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U895 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U896 ( .A(n973), .B(n1832), .Y(n189) );
  AND2X1 U897 ( .A(n1832), .B(n1528), .Y(n289) );
  INVX1 U898 ( .A(n1017), .Y(n1016) );
  AND2X1 U899 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U900 ( .A(n348), .Y(n372) );
  AND2X1 U901 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U902 ( .A(n379), .Y(n381) );
  AND2X1 U903 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U904 ( .A(n386), .Y(n387) );
  AND2X1 U905 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U906 ( .A(n401), .Y(n402) );
  BUFX2 U907 ( .A(n1343), .Y(n408) );
  BUFX2 U908 ( .A(n1356), .Y(n409) );
  BUFX2 U909 ( .A(n1369), .Y(n421) );
  BUFX2 U910 ( .A(n1382), .Y(n422) );
  BUFX2 U911 ( .A(n1395), .Y(n434) );
  BUFX2 U912 ( .A(n1408), .Y(n435) );
  BUFX2 U913 ( .A(n1498), .Y(n447) );
  BUFX2 U914 ( .A(n1509), .Y(n448) );
  AND2X2 U915 ( .A(rd), .B(n1512), .Y(n460) );
  INVX1 U916 ( .A(n460), .Y(n461) );
  INVX1 U917 ( .A(n1318), .Y(n473) );
  INVX1 U918 ( .A(n1319), .Y(n474) );
  INVX1 U919 ( .A(n1320), .Y(n486) );
  INVX1 U920 ( .A(n1411), .Y(n487) );
  INVX1 U921 ( .A(n1412), .Y(n507) );
  INVX1 U922 ( .A(n1413), .Y(n508) );
  INVX1 U923 ( .A(n1422), .Y(n522) );
  INVX1 U924 ( .A(n1423), .Y(n523) );
  INVX1 U925 ( .A(n1424), .Y(n537) );
  INVX1 U926 ( .A(n1433), .Y(n538) );
  INVX1 U927 ( .A(n1434), .Y(n552) );
  INVX1 U928 ( .A(n1435), .Y(n553) );
  INVX1 U929 ( .A(n1444), .Y(n567) );
  INVX1 U930 ( .A(n1445), .Y(n568) );
  INVX1 U931 ( .A(n1446), .Y(n582) );
  INVX1 U932 ( .A(n1455), .Y(n583) );
  INVX1 U933 ( .A(n1456), .Y(n591) );
  INVX1 U934 ( .A(n1457), .Y(n592) );
  INVX1 U935 ( .A(n1466), .Y(n871) );
  INVX1 U936 ( .A(n1467), .Y(n872) );
  INVX1 U937 ( .A(n1468), .Y(n873) );
  INVX1 U938 ( .A(n1477), .Y(n874) );
  INVX1 U939 ( .A(n1478), .Y(n875) );
  INVX1 U940 ( .A(n1479), .Y(n876) );
  AND2X2 U941 ( .A(n1332), .B(n1331), .Y(n877) );
  INVX1 U942 ( .A(n877), .Y(n878) );
  AND2X2 U943 ( .A(n1345), .B(n1344), .Y(n879) );
  INVX1 U944 ( .A(n879), .Y(n880) );
  AND2X2 U945 ( .A(n1358), .B(n1357), .Y(n881) );
  INVX1 U946 ( .A(n881), .Y(n882) );
  AND2X2 U947 ( .A(n1371), .B(n1370), .Y(n883) );
  INVX1 U948 ( .A(n883), .Y(n884) );
  AND2X2 U949 ( .A(n1384), .B(n1383), .Y(n885) );
  INVX1 U950 ( .A(n885), .Y(n886) );
  AND2X2 U951 ( .A(n1397), .B(n1396), .Y(n887) );
  INVX1 U952 ( .A(n887), .Y(n888) );
  AND2X2 U953 ( .A(n1487), .B(n1486), .Y(n889) );
  INVX1 U954 ( .A(n889), .Y(n890) );
  AND2X2 U955 ( .A(n1500), .B(n1499), .Y(n891) );
  INVX1 U956 ( .A(n891), .Y(n892) );
  INVX1 U957 ( .A(n1325), .Y(n893) );
  INVX1 U958 ( .A(n1326), .Y(n894) );
  INVX1 U959 ( .A(n1327), .Y(n895) );
  INVX1 U960 ( .A(n1416), .Y(n896) );
  INVX1 U961 ( .A(n1417), .Y(n897) );
  INVX1 U962 ( .A(n1418), .Y(n898) );
  INVX1 U963 ( .A(n1427), .Y(n899) );
  INVX1 U964 ( .A(n1428), .Y(n900) );
  INVX1 U965 ( .A(n1429), .Y(n901) );
  INVX1 U966 ( .A(n1438), .Y(n902) );
  INVX1 U967 ( .A(n1439), .Y(n903) );
  INVX1 U968 ( .A(n1440), .Y(n904) );
  INVX1 U969 ( .A(n1449), .Y(n905) );
  INVX1 U970 ( .A(n1450), .Y(n906) );
  INVX1 U971 ( .A(n1451), .Y(n907) );
  INVX1 U972 ( .A(n1460), .Y(n908) );
  INVX1 U973 ( .A(n1461), .Y(n909) );
  INVX1 U974 ( .A(n1462), .Y(n910) );
  INVX1 U975 ( .A(n1471), .Y(n911) );
  INVX1 U976 ( .A(n1472), .Y(n912) );
  INVX1 U977 ( .A(n1473), .Y(n913) );
  INVX1 U978 ( .A(n1482), .Y(n914) );
  INVX1 U979 ( .A(n1483), .Y(n915) );
  INVX1 U980 ( .A(n1484), .Y(n916) );
  AND2X2 U981 ( .A(n1334), .B(n1333), .Y(n917) );
  INVX1 U982 ( .A(n917), .Y(n918) );
  AND2X2 U983 ( .A(n1347), .B(n1346), .Y(n919) );
  INVX1 U984 ( .A(n919), .Y(n920) );
  AND2X2 U985 ( .A(n1360), .B(n1359), .Y(n921) );
  INVX1 U986 ( .A(n921), .Y(n922) );
  AND2X2 U987 ( .A(n1373), .B(n1372), .Y(n923) );
  INVX1 U988 ( .A(n923), .Y(n924) );
  AND2X2 U989 ( .A(n1386), .B(n1385), .Y(n925) );
  INVX1 U990 ( .A(n925), .Y(n926) );
  AND2X2 U991 ( .A(n1399), .B(n1398), .Y(n927) );
  INVX1 U992 ( .A(n927), .Y(n928) );
  AND2X2 U993 ( .A(n1489), .B(n1488), .Y(n929) );
  INVX1 U994 ( .A(n929), .Y(n930) );
  AND2X2 U995 ( .A(n1502), .B(n1501), .Y(n931) );
  INVX1 U996 ( .A(n931), .Y(n932) );
  BUFX2 U997 ( .A(n1341), .Y(n933) );
  BUFX2 U998 ( .A(n1354), .Y(n934) );
  BUFX2 U999 ( .A(n1367), .Y(n935) );
  BUFX2 U1000 ( .A(n1380), .Y(n936) );
  BUFX2 U1001 ( .A(n1393), .Y(n937) );
  BUFX2 U1002 ( .A(n1406), .Y(n938) );
  BUFX2 U1003 ( .A(n1496), .Y(n939) );
  INVX1 U1004 ( .A(n970), .Y(n940) );
  INVX1 U1005 ( .A(n1503), .Y(n941) );
  INVX1 U1006 ( .A(n1504), .Y(n942) );
  BUFX2 U1007 ( .A(n1556), .Y(n970) );
  BUFX2 U1008 ( .A(n1842), .Y(err) );
  BUFX2 U1009 ( .A(n1339), .Y(n944) );
  BUFX2 U1010 ( .A(n1352), .Y(n945) );
  BUFX2 U1011 ( .A(n1365), .Y(n946) );
  BUFX2 U1012 ( .A(n1378), .Y(n947) );
  BUFX2 U1013 ( .A(n1391), .Y(n948) );
  BUFX2 U1014 ( .A(n1404), .Y(n949) );
  BUFX2 U1015 ( .A(n1494), .Y(n950) );
  INVX1 U1016 ( .A(n971), .Y(n951) );
  INVX1 U1017 ( .A(n1505), .Y(n952) );
  INVX1 U1018 ( .A(n1506), .Y(n953) );
  BUFX2 U1019 ( .A(n1518), .Y(n971) );
  BUFX2 U1020 ( .A(n1527), .Y(n972) );
  BUFX2 U1021 ( .A(n1545), .Y(n974) );
  BUFX2 U1022 ( .A(n1555), .Y(n975) );
  BUFX2 U1023 ( .A(n1565), .Y(n976) );
  BUFX2 U1024 ( .A(n1575), .Y(n977) );
  BUFX2 U1025 ( .A(n1584), .Y(n978) );
  BUFX2 U1026 ( .A(n1594), .Y(n979) );
  BUFX2 U1027 ( .A(n1614), .Y(n982) );
  BUFX2 U1028 ( .A(n1633), .Y(n985) );
  BUFX2 U1029 ( .A(n1654), .Y(n988) );
  BUFX2 U1030 ( .A(n1674), .Y(n991) );
  BUFX2 U1031 ( .A(n1683), .Y(n992) );
  BUFX2 U1032 ( .A(n1693), .Y(n993) );
  BUFX2 U1033 ( .A(n1702), .Y(n994) );
  BUFX2 U1034 ( .A(n1712), .Y(n995) );
  BUFX2 U1035 ( .A(n1721), .Y(n996) );
  BUFX2 U1036 ( .A(n1731), .Y(n997) );
  BUFX2 U1037 ( .A(n1740), .Y(n998) );
  BUFX2 U1038 ( .A(n1750), .Y(n999) );
  BUFX2 U1039 ( .A(n1769), .Y(n1002) );
  BUFX2 U1040 ( .A(n1789), .Y(n1005) );
  BUFX2 U1041 ( .A(n1809), .Y(n1008) );
  BUFX2 U1042 ( .A(n1822), .Y(n973) );
  AND2X1 U1043 ( .A(n1634), .B(n1322), .Y(n1821) );
  BUFX2 U1044 ( .A(n1841), .Y(n1011) );
  BUFX2 U1045 ( .A(n1604), .Y(n954) );
  BUFX2 U1046 ( .A(n1623), .Y(n955) );
  BUFX2 U1047 ( .A(n1644), .Y(n956) );
  BUFX2 U1048 ( .A(n1664), .Y(n957) );
  BUFX2 U1049 ( .A(n1759), .Y(n958) );
  BUFX2 U1050 ( .A(n1779), .Y(n959) );
  BUFX2 U1051 ( .A(n1799), .Y(n960) );
  BUFX2 U1052 ( .A(n1820), .Y(n961) );
  AND2X1 U1053 ( .A(enable), .B(n1017), .Y(n962) );
  INVX1 U1054 ( .A(n962), .Y(n963) );
  AND2X1 U1055 ( .A(n1517), .B(n1516), .Y(n964) );
  INVX1 U1056 ( .A(n964), .Y(n965) );
  INVX1 U1057 ( .A(n966), .Y(n967) );
  INVX1 U1058 ( .A(n968), .Y(n969) );
  AND2X1 U1059 ( .A(n951), .B(n1314), .Y(n1528) );
  INVX1 U1060 ( .A(rd), .Y(n1026) );
  INVX1 U1061 ( .A(wr), .Y(n1027) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module cache2way_mem_type0 ( enable, clk, rst, createdump, .tag_in({
        \tag_in<4> , \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), 
    .index({\index<7> , \index<6> , \index<5> , \index<4> , \index<3> , 
        \index<2> , \index<1> , \index<0> }), .offset({\offset<2> , 
        \offset<1> , \offset<0> }), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        comp, write, valid_in, invert_victimway, .tag_out({\tag_out<4> , 
        \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> }), .data_out({
        \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> , 
        \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> , 
        \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> , 
        \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> }), hit, 
        dirty, valid, err );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in, invert_victimway;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   \tag_out0<4> , \tag_out0<3> , \tag_out0<2> , \tag_out0<1> ,
         \tag_out0<0> , \data_out0<15> , \data_out0<14> , \data_out0<13> ,
         \data_out0<12> , \data_out0<11> , \data_out0<10> , \data_out0<9> ,
         \data_out0<8> , \data_out0<7> , \data_out0<6> , \data_out0<5> ,
         \data_out0<4> , \data_out0<3> , \data_out0<2> , \data_out0<1> ,
         \data_out0<0> , hit0, dirty0, valid0, err0, \tag_out1<4> ,
         \tag_out1<3> , \tag_out1<2> , \tag_out1<1> , \tag_out1<0> ,
         \data_out1<15> , \data_out1<14> , \data_out1<13> , \data_out1<12> ,
         \data_out1<11> , \data_out1<10> , \data_out1<9> , \data_out1<8> ,
         \data_out1<7> , \data_out1<6> , \data_out1<5> , \data_out1<4> ,
         \data_out1<3> , \data_out1<2> , \data_out1<1> , \data_out1<0> , hit1,
         dirty1, valid1, err1, write1, selectedCache, victimway, victimwayIn,
         selectedCacheIn, n37, net88916, net102974, net103019, net121236,
         net121269, net121268, net121988, net121987, net125797, net126541,
         net126799, net126540, net123323, net123322, n1, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n15, n17, n19, n21, n23, n25, n27, n29, n31,
         n33, n35, n38, n40, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n164;
  assign \data_out<10>  = net126541;

  AOI22X1 U40 ( .A(n157), .B(n164), .C(n123), .D(hit0), .Y(n37) );
  XOR2X1 U41 ( .A(victimway), .B(invert_victimway), .Y(victimwayIn) );
  cache_cache_id0 c0 ( .enable(net121236), .clk(clk), .rst(n133), .createdump(
        createdump), .tag_in({\tag_in<4> , \tag_in<3> , \tag_in<2> , 
        \tag_in<1> , \tag_in<0> }), .index({\index<7> , \index<6> , \index<5> , 
        \index<4> , \index<3> , \index<2> , n135, \index<0> }), .offset({
        \offset<2> , \offset<1> , \offset<0> }), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .comp(n132), .write(net125797), .valid_in(valid_in), 
        .tag_out({\tag_out0<4> , \tag_out0<3> , \tag_out0<2> , \tag_out0<1> , 
        \tag_out0<0> }), .data_out({\data_out0<15> , \data_out0<14> , 
        \data_out0<13> , \data_out0<12> , \data_out0<11> , \data_out0<10> , 
        \data_out0<9> , \data_out0<8> , \data_out0<7> , \data_out0<6> , 
        \data_out0<5> , \data_out0<4> , \data_out0<3> , \data_out0<2> , 
        \data_out0<1> , \data_out0<0> }), .hit(hit0), .dirty(dirty0), .valid(
        valid0), .err(err0) );
  cache_cache_id2 c1 ( .enable(net121269), .clk(clk), .rst(n133), .createdump(
        createdump), .tag_in({\tag_in<4> , \tag_in<3> , \tag_in<2> , 
        \tag_in<1> , \tag_in<0> }), .index({\index<7> , \index<6> , \index<5> , 
        \index<4> , \index<3> , \index<2> , n135, n116}), .offset({\offset<2> , 
        \offset<1> , \offset<0> }), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .comp(n132), .write(write1), .valid_in(valid_in), .tag_out({
        \tag_out1<4> , \tag_out1<3> , \tag_out1<2> , \tag_out1<1> , 
        \tag_out1<0> }), .data_out({\data_out1<15> , \data_out1<14> , 
        \data_out1<13> , \data_out1<12> , \data_out1<11> , \data_out1<10> , 
        \data_out1<9> , \data_out1<8> , \data_out1<7> , \data_out1<6> , 
        \data_out1<5> , \data_out1<4> , \data_out1<3> , \data_out1<2> , 
        \data_out1<1> , \data_out1<0> }), .hit(hit1), .dirty(dirty1), .valid(
        valid1), .err(err1) );
  dff_217 victimway0 ( .q(victimway), .d(victimwayIn), .clk(clk), .rst(n133)
         );
  dff_216 selectedCache0 ( .q(selectedCache), .d(selectedCacheIn), .clk(clk), 
        .rst(n133) );
  BUFX2 U3 ( .A(net121236), .Y(n1) );
  OR2X2 U4 ( .A(n98), .B(n71), .Y(\data_out<9> ) );
  OR2X2 U5 ( .A(n70), .B(n97), .Y(\data_out<8> ) );
  INVX1 U6 ( .A(net102974), .Y(net126799) );
  OR2X1 U7 ( .A(err0), .B(err1), .Y(err) );
  BUFX2 U8 ( .A(enable), .Y(net121236) );
  INVX1 U9 ( .A(n1), .Y(net121268) );
  INVX1 U10 ( .A(n4), .Y(net125797) );
  OR2X2 U11 ( .A(n37), .B(n5), .Y(n4) );
  INVX1 U12 ( .A(write), .Y(n5) );
  INVX1 U13 ( .A(n6), .Y(n7) );
  AND2X2 U14 ( .A(\data_out0<10> ), .B(net102974), .Y(n6) );
  INVX4 U15 ( .A(net88916), .Y(net102974) );
  AND2X2 U16 ( .A(net123323), .B(n7), .Y(net126540) );
  INVX1 U17 ( .A(net126540), .Y(net126541) );
  INVX1 U18 ( .A(net123322), .Y(net123323) );
  AND2X2 U19 ( .A(net121988), .B(\data_out1<10> ), .Y(net123322) );
  INVX1 U20 ( .A(selectedCache), .Y(n164) );
  INVX4 U21 ( .A(n107), .Y(n108) );
  INVX2 U22 ( .A(n144), .Y(selectedCacheIn) );
  INVX1 U23 ( .A(valid0), .Y(n8) );
  INVX1 U24 ( .A(n8), .Y(n9) );
  INVX1 U25 ( .A(n112), .Y(n10) );
  INVX4 U26 ( .A(net102974), .Y(net103019) );
  INVX1 U27 ( .A(n149), .Y(n11) );
  OR2X2 U28 ( .A(n13), .B(net126799), .Y(n12) );
  INVX1 U29 ( .A(\data_out0<13> ), .Y(n13) );
  OR2X2 U30 ( .A(n101), .B(n74), .Y(\data_out<12> ) );
  AND2X2 U31 ( .A(n122), .B(n148), .Y(n15) );
  OR2X2 U32 ( .A(valid1), .B(n9), .Y(valid) );
  AND2X2 U33 ( .A(n55), .B(n82), .Y(n17) );
  INVX1 U34 ( .A(n17), .Y(\data_out<0> ) );
  AND2X2 U35 ( .A(n84), .B(n57), .Y(n19) );
  INVX1 U36 ( .A(n19), .Y(\data_out<1> ) );
  AND2X2 U37 ( .A(n59), .B(n86), .Y(n21) );
  INVX1 U38 ( .A(n21), .Y(\data_out<2> ) );
  AND2X2 U39 ( .A(n61), .B(n88), .Y(n23) );
  INVX1 U42 ( .A(n23), .Y(\data_out<3> ) );
  AND2X2 U43 ( .A(n90), .B(n63), .Y(n25) );
  INVX1 U44 ( .A(n25), .Y(\data_out<4> ) );
  AND2X2 U45 ( .A(n65), .B(n92), .Y(n27) );
  INVX1 U46 ( .A(n27), .Y(\data_out<5> ) );
  AND2X2 U47 ( .A(n67), .B(n94), .Y(n29) );
  INVX1 U48 ( .A(n29), .Y(\data_out<6> ) );
  AND2X2 U49 ( .A(n69), .B(n96), .Y(n31) );
  INVX1 U50 ( .A(n31), .Y(\data_out<7> ) );
  AND2X2 U51 ( .A(n73), .B(n100), .Y(n33) );
  INVX1 U52 ( .A(n33), .Y(\data_out<11> ) );
  AND2X2 U53 ( .A(n76), .B(n12), .Y(n35) );
  INVX1 U54 ( .A(n35), .Y(\data_out<13> ) );
  AND2X2 U55 ( .A(n78), .B(n103), .Y(n38) );
  INVX1 U56 ( .A(n38), .Y(\data_out<14> ) );
  AND2X2 U57 ( .A(n80), .B(n105), .Y(n40) );
  INVX1 U58 ( .A(n40), .Y(\data_out<15> ) );
  AND2X2 U59 ( .A(n111), .B(\tag_out1<0> ), .Y(n42) );
  INVX1 U60 ( .A(n42), .Y(n43) );
  AND2X2 U61 ( .A(n110), .B(\tag_out1<2> ), .Y(n44) );
  AND2X2 U62 ( .A(n111), .B(\tag_out1<3> ), .Y(n45) );
  AND2X2 U63 ( .A(n110), .B(\tag_out1<4> ), .Y(n46) );
  INVX1 U64 ( .A(n46), .Y(n47) );
  AND2X2 U65 ( .A(n144), .B(n151), .Y(n48) );
  INVX1 U66 ( .A(n48), .Y(n49) );
  AND2X2 U67 ( .A(n10), .B(selectedCacheIn), .Y(n50) );
  INVX1 U68 ( .A(n50), .Y(n51) );
  AND2X2 U69 ( .A(n151), .B(n112), .Y(n52) );
  INVX1 U70 ( .A(n52), .Y(n53) );
  AND2X2 U71 ( .A(n108), .B(\data_out1<0> ), .Y(n54) );
  INVX1 U72 ( .A(n54), .Y(n55) );
  AND2X2 U73 ( .A(n108), .B(\data_out1<1> ), .Y(n56) );
  INVX1 U74 ( .A(n56), .Y(n57) );
  AND2X2 U75 ( .A(n108), .B(\data_out1<2> ), .Y(n58) );
  INVX1 U76 ( .A(n58), .Y(n59) );
  AND2X2 U77 ( .A(n108), .B(\data_out1<3> ), .Y(n60) );
  INVX1 U78 ( .A(n60), .Y(n61) );
  AND2X2 U79 ( .A(n108), .B(\data_out1<4> ), .Y(n62) );
  INVX1 U80 ( .A(n62), .Y(n63) );
  AND2X2 U81 ( .A(n108), .B(\data_out1<5> ), .Y(n64) );
  INVX1 U82 ( .A(n64), .Y(n65) );
  AND2X2 U83 ( .A(n108), .B(\data_out1<6> ), .Y(n66) );
  INVX1 U84 ( .A(n66), .Y(n67) );
  AND2X2 U85 ( .A(n108), .B(\data_out1<7> ), .Y(n68) );
  INVX1 U86 ( .A(n68), .Y(n69) );
  AND2X2 U87 ( .A(\data_out0<8> ), .B(net102974), .Y(n70) );
  AND2X2 U88 ( .A(n108), .B(\data_out1<9> ), .Y(n71) );
  AND2X2 U89 ( .A(net121988), .B(\data_out1<11> ), .Y(n72) );
  INVX1 U90 ( .A(n72), .Y(n73) );
  AND2X2 U91 ( .A(n108), .B(\data_out1<12> ), .Y(n74) );
  AND2X2 U92 ( .A(n108), .B(\data_out1<13> ), .Y(n75) );
  INVX1 U93 ( .A(n75), .Y(n76) );
  AND2X2 U94 ( .A(n108), .B(\data_out1<14> ), .Y(n77) );
  INVX1 U95 ( .A(n77), .Y(n78) );
  AND2X2 U96 ( .A(n108), .B(\data_out1<15> ), .Y(n79) );
  INVX1 U97 ( .A(n79), .Y(n80) );
  AND2X2 U98 ( .A(\data_out0<0> ), .B(net102974), .Y(n81) );
  INVX1 U99 ( .A(n81), .Y(n82) );
  AND2X2 U100 ( .A(\data_out0<1> ), .B(net102974), .Y(n83) );
  INVX1 U101 ( .A(n83), .Y(n84) );
  AND2X2 U102 ( .A(\data_out0<2> ), .B(net102974), .Y(n85) );
  INVX1 U103 ( .A(n85), .Y(n86) );
  AND2X2 U104 ( .A(\data_out0<3> ), .B(net102974), .Y(n87) );
  INVX1 U105 ( .A(n87), .Y(n88) );
  AND2X2 U106 ( .A(\data_out0<4> ), .B(net102974), .Y(n89) );
  INVX1 U107 ( .A(n89), .Y(n90) );
  AND2X2 U108 ( .A(\data_out0<5> ), .B(net102974), .Y(n91) );
  INVX1 U109 ( .A(n91), .Y(n92) );
  AND2X2 U110 ( .A(\data_out0<6> ), .B(net102974), .Y(n93) );
  INVX1 U111 ( .A(n93), .Y(n94) );
  AND2X2 U112 ( .A(\data_out0<7> ), .B(net102974), .Y(n95) );
  INVX1 U113 ( .A(n95), .Y(n96) );
  AND2X2 U114 ( .A(net121988), .B(\data_out1<8> ), .Y(n97) );
  AND2X2 U115 ( .A(\data_out0<9> ), .B(net102974), .Y(n98) );
  AND2X2 U116 ( .A(\data_out0<11> ), .B(net102974), .Y(n99) );
  INVX1 U117 ( .A(n99), .Y(n100) );
  AND2X2 U118 ( .A(\data_out0<12> ), .B(net102974), .Y(n101) );
  AND2X2 U119 ( .A(\data_out0<14> ), .B(net102974), .Y(n102) );
  INVX1 U120 ( .A(n102), .Y(n103) );
  AND2X2 U121 ( .A(\data_out0<15> ), .B(net102974), .Y(n104) );
  INVX1 U122 ( .A(n104), .Y(n105) );
  BUFX2 U123 ( .A(n150), .Y(n106) );
  AND2X2 U124 ( .A(n151), .B(n121), .Y(n107) );
  AND2X2 U125 ( .A(n151), .B(n121), .Y(net121987) );
  INVX1 U126 ( .A(net121987), .Y(net121988) );
  AND2X2 U127 ( .A(n151), .B(n51), .Y(n109) );
  INVX1 U128 ( .A(n109), .Y(n110) );
  INVX1 U129 ( .A(n109), .Y(n111) );
  OR2X2 U130 ( .A(n130), .B(n125), .Y(n112) );
  AND2X2 U131 ( .A(n53), .B(n49), .Y(n145) );
  INVX2 U132 ( .A(n125), .Y(n151) );
  AND2X2 U133 ( .A(n140), .B(n139), .Y(n113) );
  INVX1 U134 ( .A(n10), .Y(hit) );
  INVX1 U135 ( .A(net121268), .Y(net121269) );
  INVX1 U136 ( .A(\index<0> ), .Y(n115) );
  INVX1 U137 ( .A(n115), .Y(n116) );
  OR2X2 U138 ( .A(n112), .B(n144), .Y(n121) );
  AND2X2 U139 ( .A(n111), .B(\tag_out1<1> ), .Y(n117) );
  INVX1 U140 ( .A(n117), .Y(n118) );
  INVX1 U141 ( .A(n44), .Y(n119) );
  INVX1 U142 ( .A(n45), .Y(n120) );
  INVX1 U143 ( .A(dirty1), .Y(n146) );
  INVX1 U144 ( .A(dirty0), .Y(n147) );
  INVX1 U145 ( .A(valid0), .Y(n122) );
  OAI21X1 U146 ( .A(valid1), .B(n141), .C(write), .Y(n142) );
  INVX1 U147 ( .A(n143), .Y(n141) );
  INVX1 U148 ( .A(n122), .Y(n123) );
  INVX1 U149 ( .A(n113), .Y(n124) );
  AND2X2 U150 ( .A(valid1), .B(n127), .Y(n125) );
  INVX1 U151 ( .A(\index<1> ), .Y(n136) );
  INVX1 U152 ( .A(n136), .Y(n135) );
  INVX1 U153 ( .A(hit1), .Y(n126) );
  INVX1 U154 ( .A(n126), .Y(n127) );
  INVX1 U155 ( .A(\tag_out0<3> ), .Y(n155) );
  INVX1 U156 ( .A(\tag_out0<4> ), .Y(n156) );
  INVX1 U157 ( .A(\tag_out0<2> ), .Y(n154) );
  INVX1 U158 ( .A(\tag_out0<1> ), .Y(n153) );
  INVX1 U159 ( .A(hit1), .Y(n128) );
  INVX1 U160 ( .A(n126), .Y(n129) );
  INVX1 U161 ( .A(valid1), .Y(n137) );
  AND2X2 U162 ( .A(n11), .B(valid0), .Y(n130) );
  INVX1 U163 ( .A(\tag_out0<0> ), .Y(n152) );
  INVX1 U164 ( .A(hit0), .Y(n149) );
  INVX2 U165 ( .A(comp), .Y(n131) );
  INVX8 U166 ( .A(n131), .Y(n132) );
  INVX1 U167 ( .A(n132), .Y(n157) );
  INVX8 U168 ( .A(n134), .Y(n133) );
  INVX8 U169 ( .A(rst), .Y(n134) );
  OR2X2 U170 ( .A(n127), .B(n157), .Y(n148) );
  OR2X2 U171 ( .A(n132), .B(selectedCache), .Y(n140) );
  NOR3X1 U172 ( .A(victimway), .B(n129), .C(n137), .Y(n138) );
  OAI21X1 U173 ( .A(n11), .B(n138), .C(n132), .Y(n139) );
  OAI21X1 U174 ( .A(n148), .B(n9), .C(n113), .Y(n144) );
  OR2X2 U175 ( .A(n132), .B(n164), .Y(n143) );
  AOI21X1 U176 ( .A(n143), .B(n128), .C(n142), .Y(write1) );
  MUX2X1 U177 ( .B(n147), .A(n146), .S(n145), .Y(dirty) );
  AOI21X1 U178 ( .A(n123), .B(n149), .C(n15), .Y(n150) );
  OAI21X1 U179 ( .A(n124), .B(n106), .C(n151), .Y(net88916) );
  OAI21X1 U180 ( .A(net103019), .B(n152), .C(n43), .Y(\tag_out<0> ) );
  OAI21X1 U181 ( .A(net103019), .B(n153), .C(n118), .Y(\tag_out<1> ) );
  OAI21X1 U182 ( .A(net103019), .B(n154), .C(n119), .Y(\tag_out<2> ) );
  OAI21X1 U183 ( .A(net103019), .B(n155), .C(n120), .Y(\tag_out<3> ) );
  OAI21X1 U184 ( .A(net103019), .B(n156), .C(n47), .Y(\tag_out<4> ) );
endmodule


module four_bank_mem ( clk, rst, createdump, .addr({\addr<15> , \addr<14> , 
        \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> , 
        \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> , 
        \addr<1> , \addr<0> }), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        wr, rd, .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), stall, .busy({\busy<3> , \busy<2> , \busy<1> , 
        \busy<0> }), err );
  input clk, rst, createdump, \addr<15> , \addr<14> , \addr<13> , \addr<12> ,
         \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> ,
         \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> ,
         \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , wr, rd;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , stall,
         \busy<3> , \busy<2> , \busy<1> , \busy<0> , err;
  wire   n121, \en<3> , \en<2> , \en<1> , \en<0> , \data0_out<15> ,
         \data0_out<14> , \data0_out<13> , \data0_out<12> , \data0_out<11> ,
         \data0_out<10> , \data0_out<9> , \data0_out<8> , \data0_out<7> ,
         \data0_out<6> , \data0_out<5> , \data0_out<4> , \data0_out<3> ,
         \data0_out<2> , \data0_out<1> , \data0_out<0> , err0, \data1_out<15> ,
         \data1_out<14> , \data1_out<13> , \data1_out<12> , \data1_out<11> ,
         \data1_out<10> , \data1_out<9> , \data1_out<8> , \data1_out<7> ,
         \data1_out<6> , \data1_out<5> , \data1_out<4> , \data1_out<3> ,
         \data1_out<2> , \data1_out<1> , \data1_out<0> , err1, \data2_out<15> ,
         \data2_out<14> , \data2_out<13> , \data2_out<12> , \data2_out<11> ,
         \data2_out<10> , \data2_out<9> , \data2_out<8> , \data2_out<7> ,
         \data2_out<6> , \data2_out<5> , \data2_out<4> , \data2_out<3> ,
         \data2_out<2> , \data2_out<1> , \data2_out<0> , err2, \data3_out<15> ,
         \data3_out<14> , \data3_out<13> , \data3_out<12> , \data3_out<11> ,
         \data3_out<10> , \data3_out<9> , \data3_out<8> , \data3_out<7> ,
         \data3_out<6> , \data3_out<5> , \data3_out<4> , \data3_out<3> ,
         \data3_out<2> , \data3_out<1> , \data3_out<0> , err3, \bsy0<3> ,
         \bsy0<2> , \bsy0<1> , \bsy0<0> , \bsy1<3> , \bsy1<2> , \bsy1<1> ,
         \bsy1<0> , \bsy2<3> , \bsy2<2> , \bsy2<1> , \bsy2<0> , n9, n10, n11,
         n13, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n1, n2, n3, n4, n5, n6, n7,
         n12, n15, n18, n21, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74,
         n76, n78, n79, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116;

  NOR3X1 U9 ( .A(n97), .B(n98), .C(n2), .Y(stall) );
  OAI21X1 U11 ( .A(\addr<1> ), .B(n11), .C(n6), .Y(n10) );
  OAI21X1 U13 ( .A(\addr<1> ), .B(n13), .C(n4), .Y(n9) );
  AOI21X1 U15 ( .A(n84), .B(n16), .C(n97), .Y(n121) );
  NOR3X1 U16 ( .A(err1), .B(err3), .C(err2), .Y(n16) );
  NOR3X1 U18 ( .A(n92), .B(\busy<3> ), .C(n97), .Y(\en<3> ) );
  NOR3X1 U20 ( .A(n90), .B(n97), .C(n95), .Y(\en<2> ) );
  NOR3X1 U22 ( .A(n88), .B(n97), .C(n116), .Y(\en<1> ) );
  NOR3X1 U24 ( .A(n86), .B(\busy<0> ), .C(n97), .Y(\en<0> ) );
  NOR2X1 U28 ( .A(\data3_out<9> ), .B(\data2_out<9> ), .Y(n23) );
  NOR2X1 U29 ( .A(\data1_out<9> ), .B(\data0_out<9> ), .Y(n22) );
  NOR2X1 U31 ( .A(\data3_out<8> ), .B(\data2_out<8> ), .Y(n25) );
  NOR2X1 U32 ( .A(\data1_out<8> ), .B(\data0_out<8> ), .Y(n24) );
  NOR2X1 U34 ( .A(\data3_out<7> ), .B(\data2_out<7> ), .Y(n27) );
  NOR2X1 U35 ( .A(\data1_out<7> ), .B(\data0_out<7> ), .Y(n26) );
  NOR2X1 U37 ( .A(\data3_out<6> ), .B(\data2_out<6> ), .Y(n29) );
  NOR2X1 U38 ( .A(\data1_out<6> ), .B(\data0_out<6> ), .Y(n28) );
  NOR2X1 U40 ( .A(\data3_out<5> ), .B(\data2_out<5> ), .Y(n31) );
  NOR2X1 U41 ( .A(\data1_out<5> ), .B(\data0_out<5> ), .Y(n30) );
  NOR2X1 U43 ( .A(\data3_out<4> ), .B(\data2_out<4> ), .Y(n33) );
  NOR2X1 U44 ( .A(\data1_out<4> ), .B(\data0_out<4> ), .Y(n32) );
  NOR2X1 U46 ( .A(\data3_out<3> ), .B(\data2_out<3> ), .Y(n35) );
  NOR2X1 U47 ( .A(\data1_out<3> ), .B(\data0_out<3> ), .Y(n34) );
  NOR2X1 U49 ( .A(\data3_out<2> ), .B(\data2_out<2> ), .Y(n37) );
  NOR2X1 U50 ( .A(\data1_out<2> ), .B(\data0_out<2> ), .Y(n36) );
  NOR2X1 U52 ( .A(\data3_out<1> ), .B(\data2_out<1> ), .Y(n39) );
  NOR2X1 U53 ( .A(\data1_out<1> ), .B(\data0_out<1> ), .Y(n38) );
  NOR2X1 U55 ( .A(\data3_out<15> ), .B(\data2_out<15> ), .Y(n41) );
  NOR2X1 U56 ( .A(\data1_out<15> ), .B(\data0_out<15> ), .Y(n40) );
  NOR2X1 U58 ( .A(\data3_out<14> ), .B(\data2_out<14> ), .Y(n43) );
  NOR2X1 U59 ( .A(\data1_out<14> ), .B(\data0_out<14> ), .Y(n42) );
  NOR2X1 U61 ( .A(\data3_out<13> ), .B(\data2_out<13> ), .Y(n45) );
  NOR2X1 U62 ( .A(\data1_out<13> ), .B(\data0_out<13> ), .Y(n44) );
  NOR2X1 U64 ( .A(\data3_out<12> ), .B(\data2_out<12> ), .Y(n47) );
  NOR2X1 U65 ( .A(\data1_out<12> ), .B(\data0_out<12> ), .Y(n46) );
  NOR2X1 U67 ( .A(\data3_out<11> ), .B(\data2_out<11> ), .Y(n49) );
  NOR2X1 U68 ( .A(\data1_out<11> ), .B(\data0_out<11> ), .Y(n48) );
  NOR2X1 U70 ( .A(\data3_out<10> ), .B(\data2_out<10> ), .Y(n51) );
  NOR2X1 U71 ( .A(\data1_out<10> ), .B(\data0_out<10> ), .Y(n50) );
  NOR2X1 U73 ( .A(\data3_out<0> ), .B(\data2_out<0> ), .Y(n53) );
  NOR2X1 U74 ( .A(\data1_out<0> ), .B(\data0_out<0> ), .Y(n52) );
  NOR3X1 U75 ( .A(\bsy0<3> ), .B(\bsy2<3> ), .C(\bsy1<3> ), .Y(n54) );
  NOR3X1 U76 ( .A(\bsy0<2> ), .B(\bsy2<2> ), .C(\bsy1<2> ), .Y(n11) );
  NOR3X1 U77 ( .A(\bsy0<1> ), .B(\bsy2<1> ), .C(\bsy1<1> ), .Y(n20) );
  NOR3X1 U78 ( .A(\bsy0<0> ), .B(\bsy2<0> ), .C(\bsy1<0> ), .Y(n13) );
  final_memory_3 m0 ( .data_out({\data0_out<15> , \data0_out<14> , 
        \data0_out<13> , \data0_out<12> , \data0_out<11> , \data0_out<10> , 
        \data0_out<9> , \data0_out<8> , \data0_out<7> , \data0_out<6> , 
        \data0_out<5> , \data0_out<4> , \data0_out<3> , \data0_out<2> , 
        \data0_out<1> , \data0_out<0> }), .err(err0), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<0> ), .create_dump(createdump), .bank_id({1'b0, 
        1'b0}), .clk(clk), .rst(n98) );
  final_memory_2 m1 ( .data_out({\data1_out<15> , \data1_out<14> , 
        \data1_out<13> , \data1_out<12> , \data1_out<11> , \data1_out<10> , 
        \data1_out<9> , \data1_out<8> , \data1_out<7> , \data1_out<6> , 
        \data1_out<5> , \data1_out<4> , \data1_out<3> , \data1_out<2> , 
        \data1_out<1> , \data1_out<0> }), .err(err1), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<1> ), .create_dump(createdump), .bank_id({1'b0, 
        1'b1}), .clk(clk), .rst(n98) );
  final_memory_1 m2 ( .data_out({\data2_out<15> , \data2_out<14> , 
        \data2_out<13> , \data2_out<12> , \data2_out<11> , \data2_out<10> , 
        \data2_out<9> , \data2_out<8> , \data2_out<7> , \data2_out<6> , 
        \data2_out<5> , \data2_out<4> , \data2_out<3> , \data2_out<2> , 
        \data2_out<1> , \data2_out<0> }), .err(err2), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<2> ), .create_dump(createdump), .bank_id({1'b1, 
        1'b0}), .clk(clk), .rst(n98) );
  final_memory_0 m3 ( .data_out({\data3_out<15> , \data3_out<14> , 
        \data3_out<13> , \data3_out<12> , \data3_out<11> , \data3_out<10> , 
        \data3_out<9> , \data3_out<8> , \data3_out<7> , \data3_out<6> , 
        \data3_out<5> , \data3_out<4> , \data3_out<3> , \data3_out<2> , 
        \data3_out<1> , \data3_out<0> }), .err(err3), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n114, n112, n110, n108, n106, n104, n102, n100}), .wr(wr), 
        .rd(rd), .enable(\en<3> ), .create_dump(createdump), .bank_id({1'b1, 
        1'b1}), .clk(clk), .rst(n98) );
  dff_212 \b0[0]  ( .q(\bsy0<0> ), .d(\en<0> ), .clk(clk), .rst(n98) );
  dff_213 \b0[1]  ( .q(\bsy0<1> ), .d(\en<1> ), .clk(clk), .rst(n98) );
  dff_214 \b0[2]  ( .q(\bsy0<2> ), .d(\en<2> ), .clk(clk), .rst(n98) );
  dff_215 \b0[3]  ( .q(\bsy0<3> ), .d(\en<3> ), .clk(clk), .rst(n98) );
  dff_208 \b1[0]  ( .q(\bsy1<0> ), .d(\bsy0<0> ), .clk(clk), .rst(n98) );
  dff_209 \b1[1]  ( .q(\bsy1<1> ), .d(\bsy0<1> ), .clk(clk), .rst(n98) );
  dff_210 \b1[2]  ( .q(\bsy1<2> ), .d(\bsy0<2> ), .clk(clk), .rst(n98) );
  dff_211 \b1[3]  ( .q(\bsy1<3> ), .d(\bsy0<3> ), .clk(clk), .rst(n98) );
  dff_204 \b2[0]  ( .q(\bsy2<0> ), .d(\bsy1<0> ), .clk(clk), .rst(n98) );
  dff_205 \b2[1]  ( .q(\bsy2<1> ), .d(\bsy1<1> ), .clk(clk), .rst(n98) );
  dff_206 \b2[2]  ( .q(\bsy2<2> ), .d(\bsy1<2> ), .clk(clk), .rst(n98) );
  dff_207 \b2[3]  ( .q(\bsy2<3> ), .d(\bsy1<3> ), .clk(clk), .rst(n98) );
  INVX1 U3 ( .A(n54), .Y(\busy<3> ) );
  INVX1 U4 ( .A(rst), .Y(n99) );
  INVX1 U5 ( .A(n13), .Y(\busy<0> ) );
  AND2X1 U6 ( .A(\addr<2> ), .B(\addr<1> ), .Y(n91) );
  INVX1 U7 ( .A(n101), .Y(n100) );
  INVX1 U8 ( .A(n103), .Y(n102) );
  INVX1 U10 ( .A(n105), .Y(n104) );
  INVX1 U12 ( .A(\addr<5> ), .Y(n105) );
  INVX1 U14 ( .A(n107), .Y(n106) );
  INVX1 U17 ( .A(\addr<6> ), .Y(n107) );
  INVX1 U19 ( .A(n109), .Y(n108) );
  INVX1 U21 ( .A(\addr<7> ), .Y(n109) );
  INVX1 U23 ( .A(n111), .Y(n110) );
  INVX1 U25 ( .A(\addr<8> ), .Y(n111) );
  INVX1 U26 ( .A(n113), .Y(n112) );
  INVX1 U27 ( .A(\addr<9> ), .Y(n113) );
  INVX1 U30 ( .A(n115), .Y(n114) );
  INVX1 U33 ( .A(\addr<10> ), .Y(n115) );
  AND2X1 U36 ( .A(\addr<1> ), .B(\busy<1> ), .Y(n3) );
  INVX1 U39 ( .A(n20), .Y(\busy<1> ) );
  AND2X1 U42 ( .A(\addr<1> ), .B(\busy<3> ), .Y(n5) );
  OR2X1 U45 ( .A(err0), .B(\addr<0> ), .Y(n83) );
  INVX1 U48 ( .A(n11), .Y(\busy<2> ) );
  INVX1 U51 ( .A(n99), .Y(n98) );
  OR2X1 U54 ( .A(n79), .B(n82), .Y(n1) );
  INVX1 U57 ( .A(n1), .Y(n2) );
  INVX1 U60 ( .A(n3), .Y(n4) );
  INVX1 U63 ( .A(n5), .Y(n6) );
  AND2X2 U66 ( .A(n52), .B(n53), .Y(n7) );
  INVX1 U69 ( .A(n7), .Y(\data_out<0> ) );
  AND2X2 U72 ( .A(n50), .B(n51), .Y(n12) );
  INVX1 U79 ( .A(n12), .Y(\data_out<10> ) );
  AND2X2 U80 ( .A(n48), .B(n49), .Y(n15) );
  INVX1 U81 ( .A(n15), .Y(\data_out<11> ) );
  AND2X2 U82 ( .A(n46), .B(n47), .Y(n18) );
  INVX1 U83 ( .A(n18), .Y(\data_out<12> ) );
  AND2X2 U84 ( .A(n44), .B(n45), .Y(n21) );
  INVX1 U85 ( .A(n21), .Y(\data_out<13> ) );
  AND2X2 U86 ( .A(n42), .B(n43), .Y(n56) );
  INVX1 U87 ( .A(n56), .Y(\data_out<14> ) );
  AND2X2 U88 ( .A(n40), .B(n41), .Y(n58) );
  INVX1 U89 ( .A(n58), .Y(\data_out<15> ) );
  AND2X2 U90 ( .A(n38), .B(n39), .Y(n60) );
  INVX1 U91 ( .A(n60), .Y(\data_out<1> ) );
  AND2X2 U92 ( .A(n36), .B(n37), .Y(n62) );
  INVX1 U93 ( .A(n62), .Y(\data_out<2> ) );
  AND2X2 U94 ( .A(n34), .B(n35), .Y(n64) );
  INVX1 U95 ( .A(n64), .Y(\data_out<3> ) );
  AND2X2 U96 ( .A(n32), .B(n33), .Y(n66) );
  INVX1 U97 ( .A(n66), .Y(\data_out<4> ) );
  AND2X2 U98 ( .A(n30), .B(n31), .Y(n68) );
  INVX1 U99 ( .A(n68), .Y(\data_out<5> ) );
  AND2X2 U100 ( .A(n28), .B(n29), .Y(n70) );
  INVX1 U101 ( .A(n70), .Y(\data_out<6> ) );
  AND2X2 U102 ( .A(n26), .B(n27), .Y(n72) );
  INVX1 U103 ( .A(n72), .Y(\data_out<7> ) );
  AND2X2 U104 ( .A(n24), .B(n25), .Y(n74) );
  INVX1 U105 ( .A(n74), .Y(\data_out<8> ) );
  AND2X2 U106 ( .A(n22), .B(n23), .Y(n76) );
  INVX1 U107 ( .A(n76), .Y(\data_out<9> ) );
  OR2X1 U108 ( .A(\addr<2> ), .B(n93), .Y(n78) );
  INVX1 U109 ( .A(n78), .Y(n79) );
  BUFX2 U110 ( .A(n121), .Y(err) );
  OR2X1 U111 ( .A(n94), .B(n95), .Y(n81) );
  INVX1 U112 ( .A(n81), .Y(n82) );
  INVX1 U113 ( .A(n83), .Y(n84) );
  AND2X1 U114 ( .A(n116), .B(n95), .Y(n85) );
  INVX1 U115 ( .A(n85), .Y(n86) );
  AND2X1 U116 ( .A(n20), .B(n95), .Y(n87) );
  INVX1 U117 ( .A(n87), .Y(n88) );
  AND2X1 U118 ( .A(n11), .B(n116), .Y(n89) );
  INVX1 U119 ( .A(n89), .Y(n90) );
  INVX1 U120 ( .A(\addr<1> ), .Y(n116) );
  INVX1 U121 ( .A(n91), .Y(n92) );
  INVX1 U122 ( .A(n9), .Y(n93) );
  INVX1 U123 ( .A(n10), .Y(n94) );
  INVX1 U124 ( .A(\addr<2> ), .Y(n95) );
  OR2X1 U125 ( .A(rd), .B(wr), .Y(n96) );
  INVX1 U126 ( .A(n96), .Y(n97) );
  INVX1 U127 ( .A(\addr<4> ), .Y(n103) );
  INVX1 U128 ( .A(\addr<3> ), .Y(n101) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module mem_system ( .DataOut({\DataOut<15> , \DataOut<14> , \DataOut<13> , 
        \DataOut<12> , \DataOut<11> , \DataOut<10> , \DataOut<9> , 
        \DataOut<8> , \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , 
        \DataOut<3> , \DataOut<2> , \DataOut<1> , \DataOut<0> }), Done, Stall, 
        CacheHit, err, .Addr({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> , \Addr<10> , \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , 
        \Addr<5> , \Addr<4> , \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> }), 
    .DataIn({\DataIn<15> , \DataIn<14> , \DataIn<13> , \DataIn<12> , 
        \DataIn<11> , \DataIn<10> , \DataIn<9> , \DataIn<8> , \DataIn<7> , 
        \DataIn<6> , \DataIn<5> , \DataIn<4> , \DataIn<3> , \DataIn<2> , 
        \DataIn<1> , \DataIn<0> }), Rd, Wr, createdump, clk, rst );
  input \Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , \Addr<11> , \Addr<10> ,
         \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , \Addr<5> , \Addr<4> ,
         \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> , \DataIn<15> ,
         \DataIn<14> , \DataIn<13> , \DataIn<12> , \DataIn<11> , \DataIn<10> ,
         \DataIn<9> , \DataIn<8> , \DataIn<7> , \DataIn<6> , \DataIn<5> ,
         \DataIn<4> , \DataIn<3> , \DataIn<2> , \DataIn<1> , \DataIn<0> , Rd,
         Wr, createdump, clk, rst;
  output \DataOut<15> , \DataOut<14> , \DataOut<13> , \DataOut<12> ,
         \DataOut<11> , \DataOut<10> , \DataOut<9> , \DataOut<8> ,
         \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , \DataOut<3> ,
         \DataOut<2> , \DataOut<1> , \DataOut<0> , Done, Stall, CacheHit, err;
  wire   \cacheTagOut<4> , \cacheTagOut<3> , \cacheTagOut<2> ,
         \cacheTagOut<1> , \cacheTagOut<0> , hit, dirty, valid, cacheErr,
         enable, \cacheAddr<2> , \cacheAddr<1> , cacheWrite, \memDataOut<15> ,
         \memDataOut<14> , \memDataOut<13> , \memDataOut<12> ,
         \memDataOut<11> , \memDataOut<10> , \memDataOut<9> , \memDataOut<8> ,
         \memDataOut<7> , \memDataOut<6> , \memDataOut<5> , \memDataOut<4> ,
         \memDataOut<3> , \memDataOut<2> , \memDataOut<1> , \memDataOut<0> ,
         mem_stall, memErr, memAddr_2, memWrite, memRead, \state<4> ,
         \state<3> , \state<2> , \state<1> , \state<0> , \next_state<4> ,
         \next_state<1> , \next_state<0> , net89031, net89037, net89083,
         net89086, net89097, net89098, net89099, net89119, net89127, net89137,
         net95739, net95788, net95941, net95995, net96034, net102554,
         net102793, net102834, net102842, net102841, net121256, net121261,
         net121272, net121515, net121753, net121828, net121827, net126586,
         net126585, net126592, net126590, net126599, net126598, net126635,
         net126634, net126654, net129873, net129927, net129926, net129930,
         net129949, net130115, net130129, net130138, net95942, net89141,
         net89072, net121245, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472;
  assign CacheHit = net121827;

  cache2way_mem_type0 cache ( .enable(enable), .clk(clk), .rst(n425), 
        .createdump(createdump), .tag_in({\Addr<15> , \Addr<14> , \Addr<13> , 
        \Addr<12> , \Addr<11> }), .index({n438, n436, n434, n432, n430, n428, 
        n422, \Addr<3> }), .offset({\cacheAddr<2> , \cacheAddr<1> , n350}), 
        .data_in({n414, n410, n408, n406, n404, n402, n400, n398, n412, n396, 
        n394, n392, n390, n388, n386, n384}), .comp(net129873), .write(n352), 
        .valid_in(1'b1), .invert_victimway(n348), .tag_out({\cacheTagOut<4> , 
        \cacheTagOut<3> , \cacheTagOut<2> , \cacheTagOut<1> , \cacheTagOut<0> }), .data_out({\DataOut<15> , \DataOut<14> , \DataOut<13> , \DataOut<12> , 
        \DataOut<11> , \DataOut<10> , \DataOut<9> , \DataOut<8> , \DataOut<7> , 
        \DataOut<6> , \DataOut<5> , \DataOut<4> , \DataOut<3> , \DataOut<2> , 
        \DataOut<1> , \DataOut<0> }), .hit(hit), .dirty(dirty), .valid(valid), 
        .err(cacheErr) );
  four_bank_mem mem ( .clk(clk), .rst(n425), .createdump(createdump), .addr({
        n162, n164, n166, n168, n170, n438, n436, n434, n432, n430, n428, n422, 
        n419, n361, n382, 1'b0}), .data_in({n224, n228, \DataOut<13> , 
        \DataOut<12> , n230, net121515, n219, \DataOut<8> , n226, n222, n234, 
        n213, n232, n217, n215, n156}), .wr(memWrite), .rd(memRead), 
        .data_out({\memDataOut<15> , \memDataOut<14> , \memDataOut<13> , 
        \memDataOut<12> , \memDataOut<11> , \memDataOut<10> , \memDataOut<9> , 
        \memDataOut<8> , \memDataOut<7> , \memDataOut<6> , \memDataOut<5> , 
        \memDataOut<4> , \memDataOut<3> , \memDataOut<2> , \memDataOut<1> , 
        \memDataOut<0> }), .stall(mem_stall), .busy(), .err(memErr) );
  dff_218 \SM_Flops[0]  ( .q(\state<0> ), .d(\next_state<0> ), .clk(clk), 
        .rst(n425) );
  dff_219 \SM_Flops[1]  ( .q(\state<1> ), .d(n241), .clk(clk), .rst(n425) );
  dff_220 \SM_Flops[2]  ( .q(\state<2> ), .d(n183), .clk(clk), .rst(n425) );
  dff_221 \SM_Flops[3]  ( .q(\state<3> ), .d(n160), .clk(clk), .rst(n425) );
  dff_222 \SM_Flops[4]  ( .q(\state<4> ), .d(\next_state<4> ), .clk(clk), 
        .rst(n425) );
  INVX1 U159 ( .A(n200), .Y(n140) );
  AND2X2 U160 ( .A(n201), .B(n196), .Y(n326) );
  INVX2 U161 ( .A(n364), .Y(n365) );
  INVX1 U162 ( .A(n206), .Y(n141) );
  INVX1 U163 ( .A(net89141), .Y(n142) );
  INVX1 U164 ( .A(net89099), .Y(n143) );
  AND2X2 U165 ( .A(n145), .B(net126598), .Y(n144) );
  INVX2 U166 ( .A(n165), .Y(n166) );
  INVX2 U167 ( .A(n161), .Y(n162) );
  INVX2 U168 ( .A(n169), .Y(n170) );
  INVX2 U169 ( .A(n167), .Y(n168) );
  AND2X2 U170 ( .A(n453), .B(n177), .Y(n195) );
  AND2X1 U171 ( .A(\memDataOut<1> ), .B(net89037), .Y(n244) );
  AND2X1 U172 ( .A(\memDataOut<3> ), .B(net89037), .Y(n248) );
  AND2X1 U173 ( .A(\memDataOut<4> ), .B(net89037), .Y(n250) );
  AND2X1 U174 ( .A(\memDataOut<0> ), .B(net89037), .Y(n242) );
  AND2X1 U175 ( .A(n257), .B(n291), .Y(n411) );
  AND2X1 U176 ( .A(n259), .B(n293), .Y(n397) );
  INVX1 U177 ( .A(\Addr<0> ), .Y(n463) );
  INVX1 U178 ( .A(n375), .Y(n468) );
  INVX1 U179 ( .A(n163), .Y(n164) );
  INVX1 U180 ( .A(rst), .Y(n426) );
  INVX1 U181 ( .A(\Addr<1> ), .Y(n464) );
  INVX1 U182 ( .A(\Addr<2> ), .Y(n466) );
  AND2X1 U183 ( .A(n245), .B(n279), .Y(n385) );
  AND2X1 U184 ( .A(n247), .B(n281), .Y(n387) );
  AND2X1 U185 ( .A(n249), .B(n283), .Y(n389) );
  AND2X1 U186 ( .A(n251), .B(n285), .Y(n391) );
  AND2X1 U187 ( .A(n253), .B(n287), .Y(n393) );
  AND2X1 U188 ( .A(n255), .B(n289), .Y(n395) );
  AND2X1 U189 ( .A(n261), .B(n295), .Y(n399) );
  AND2X1 U190 ( .A(n263), .B(n297), .Y(n401) );
  AND2X1 U191 ( .A(n265), .B(n299), .Y(n403) );
  AND2X1 U192 ( .A(n267), .B(n301), .Y(n405) );
  AND2X1 U193 ( .A(n269), .B(n303), .Y(n407) );
  AND2X1 U194 ( .A(n271), .B(n305), .Y(n409) );
  AND2X1 U195 ( .A(n375), .B(n171), .Y(n235) );
  AND2X1 U196 ( .A(n273), .B(n307), .Y(n413) );
  OR2X1 U197 ( .A(n420), .B(n330), .Y(n339) );
  INVX1 U198 ( .A(mem_stall), .Y(n452) );
  OR2X1 U199 ( .A(n327), .B(n328), .Y(n337) );
  INVX1 U200 ( .A(\Addr<6> ), .Y(n431) );
  INVX1 U201 ( .A(\Addr<7> ), .Y(n433) );
  INVX1 U202 ( .A(\Addr<8> ), .Y(n435) );
  INVX2 U203 ( .A(n437), .Y(n436) );
  INVX1 U204 ( .A(\Addr<9> ), .Y(n437) );
  INVX1 U205 ( .A(n439), .Y(n438) );
  INVX1 U206 ( .A(\Addr<10> ), .Y(n439) );
  AND2X1 U207 ( .A(n243), .B(n277), .Y(n383) );
  AND2X1 U208 ( .A(n371), .B(n196), .Y(n458) );
  OR2X1 U209 ( .A(cacheErr), .B(memErr), .Y(err) );
  AND2X1 U210 ( .A(n472), .B(n313), .Y(n182) );
  BUFX2 U211 ( .A(\DataOut<10> ), .Y(net121515) );
  NAND3X1 U212 ( .A(net130129), .B(net121272), .C(net121245), .Y(net89072) );
  INVX1 U213 ( .A(n143), .Y(net130129) );
  INVX1 U214 ( .A(\state<1> ), .Y(net121272) );
  INVX1 U215 ( .A(net89141), .Y(net121245) );
  OR2X2 U216 ( .A(\state<0> ), .B(\state<2> ), .Y(net89141) );
  OR2X2 U217 ( .A(net89072), .B(net121261), .Y(net95942) );
  BUFX2 U218 ( .A(net89072), .Y(net95995) );
  INVX1 U219 ( .A(net89141), .Y(net89097) );
  OR2X2 U220 ( .A(net89127), .B(net89141), .Y(net126654) );
  AND2X2 U221 ( .A(net95942), .B(net126654), .Y(n145) );
  INVX1 U222 ( .A(\state<4> ), .Y(net121261) );
  BUFX2 U223 ( .A(net95942), .Y(net121753) );
  NAND3X1 U224 ( .A(net95788), .B(n144), .C(n146), .Y(enable) );
  AND2X2 U225 ( .A(net89083), .B(net95739), .Y(net95788) );
  INVX1 U226 ( .A(net126585), .Y(n146) );
  OR2X2 U227 ( .A(net126635), .B(net126592), .Y(net126585) );
  INVX1 U228 ( .A(net126598), .Y(net126599) );
  AND2X1 U229 ( .A(n275), .B(n465), .Y(n336) );
  AND2X1 U230 ( .A(\cacheTagOut<0> ), .B(memWrite), .Y(n187) );
  AND2X1 U231 ( .A(\cacheTagOut<4> ), .B(memWrite), .Y(n189) );
  INVX1 U232 ( .A(n440), .Y(n147) );
  INVX1 U233 ( .A(n147), .Y(n148) );
  INVX1 U234 ( .A(n195), .Y(n149) );
  INVX1 U235 ( .A(\state<1> ), .Y(net130138) );
  INVX1 U236 ( .A(n179), .Y(n150) );
  INVX1 U237 ( .A(\state<4> ), .Y(net130115) );
  AND2X1 U238 ( .A(\cacheTagOut<2> ), .B(memWrite), .Y(n193) );
  INVX1 U239 ( .A(n152), .Y(n151) );
  AND2X1 U240 ( .A(\cacheTagOut<3> ), .B(memWrite), .Y(n191) );
  INVX1 U241 ( .A(net129926), .Y(net129949) );
  INVX1 U242 ( .A(n462), .Y(n152) );
  INVX1 U243 ( .A(n152), .Y(n153) );
  INVX1 U244 ( .A(net102842), .Y(net129930) );
  INVX1 U245 ( .A(\state<0> ), .Y(net129926) );
  INVX1 U246 ( .A(net129926), .Y(net129927) );
  AND2X2 U247 ( .A(net102841), .B(net129927), .Y(n154) );
  INVX1 U248 ( .A(\DataOut<0> ), .Y(n155) );
  INVX1 U249 ( .A(n155), .Y(n156) );
  INVX1 U250 ( .A(n446), .Y(n157) );
  INVX1 U251 ( .A(n157), .Y(n158) );
  INVX1 U252 ( .A(net126598), .Y(net129873) );
  AND2X1 U253 ( .A(n199), .B(n172), .Y(n465) );
  INVX1 U254 ( .A(n440), .Y(n462) );
  AND2X2 U255 ( .A(n451), .B(n204), .Y(n159) );
  INVX1 U256 ( .A(n159), .Y(n160) );
  AND2X2 U257 ( .A(n317), .B(n190), .Y(n161) );
  AND2X2 U258 ( .A(n319), .B(n192), .Y(n163) );
  AND2X2 U259 ( .A(n321), .B(n194), .Y(n165) );
  AND2X2 U260 ( .A(n323), .B(n315), .Y(n167) );
  AND2X2 U261 ( .A(n325), .B(n188), .Y(n169) );
  AND2X2 U262 ( .A(n380), .B(n236), .Y(n171) );
  OR2X2 U263 ( .A(n442), .B(n148), .Y(n172) );
  AND2X2 U264 ( .A(net129927), .B(net89119), .Y(n173) );
  AND2X2 U265 ( .A(n239), .B(n446), .Y(n174) );
  INVX1 U266 ( .A(n174), .Y(n175) );
  AND2X2 U267 ( .A(n158), .B(net89097), .Y(n176) );
  AND2X2 U268 ( .A(net121256), .B(net121261), .Y(n177) );
  AND2X2 U269 ( .A(n211), .B(net89098), .Y(n178) );
  AND2X2 U270 ( .A(n173), .B(n456), .Y(n179) );
  AND2X2 U271 ( .A(n154), .B(net89098), .Y(n180) );
  INVX1 U272 ( .A(n180), .Y(n181) );
  INVX1 U273 ( .A(n182), .Y(n183) );
  INVX1 U274 ( .A(n237), .Y(n184) );
  OR2X2 U275 ( .A(net126599), .B(net95941), .Y(n185) );
  INVX1 U276 ( .A(n185), .Y(n186) );
  INVX1 U277 ( .A(n187), .Y(n188) );
  INVX1 U278 ( .A(n189), .Y(n190) );
  INVX1 U279 ( .A(n191), .Y(n192) );
  INVX1 U280 ( .A(n193), .Y(n194) );
  AND2X2 U281 ( .A(n141), .B(n172), .Y(net126634) );
  INVX1 U282 ( .A(net126634), .Y(net126635) );
  INVX1 U283 ( .A(n195), .Y(n196) );
  AND2X2 U284 ( .A(n153), .B(n142), .Y(n197) );
  INVX1 U285 ( .A(n197), .Y(n198) );
  INVX1 U286 ( .A(n197), .Y(n199) );
  AND2X2 U287 ( .A(n154), .B(n158), .Y(n200) );
  INVX1 U288 ( .A(n200), .Y(n201) );
  AND2X2 U289 ( .A(n184), .B(n209), .Y(n202) );
  INVX1 U290 ( .A(n202), .Y(n203) );
  INVX1 U291 ( .A(n202), .Y(n204) );
  BUFX2 U292 ( .A(n455), .Y(n205) );
  AND2X2 U293 ( .A(n154), .B(n151), .Y(n206) );
  INVX1 U294 ( .A(n206), .Y(n207) );
  AND2X2 U295 ( .A(n150), .B(n362), .Y(net126598) );
  AND2X2 U296 ( .A(n455), .B(n175), .Y(net126590) );
  INVX1 U297 ( .A(net126590), .Y(net126592) );
  INVX1 U298 ( .A(net126585), .Y(net126586) );
  BUFX2 U299 ( .A(n467), .Y(n208) );
  BUFX2 U300 ( .A(n450), .Y(n209) );
  INVX1 U301 ( .A(n239), .Y(n210) );
  INVX1 U302 ( .A(n210), .Y(n211) );
  INVX1 U303 ( .A(net126654), .Y(net121827) );
  INVX1 U304 ( .A(net121827), .Y(net121828) );
  INVX1 U305 ( .A(\DataOut<4> ), .Y(n212) );
  INVX1 U306 ( .A(n212), .Y(n213) );
  INVX1 U307 ( .A(\DataOut<1> ), .Y(n214) );
  INVX1 U308 ( .A(n214), .Y(n215) );
  INVX1 U309 ( .A(\DataOut<2> ), .Y(n216) );
  INVX1 U310 ( .A(n216), .Y(n217) );
  INVX1 U311 ( .A(\DataOut<9> ), .Y(n218) );
  INVX1 U312 ( .A(n218), .Y(n219) );
  AND2X2 U313 ( .A(n462), .B(n239), .Y(n220) );
  INVX1 U314 ( .A(\state<3> ), .Y(net89099) );
  INVX1 U315 ( .A(\state<4> ), .Y(net89086) );
  INVX1 U316 ( .A(net130138), .Y(net121256) );
  INVX1 U317 ( .A(n444), .Y(n446) );
  INVX1 U318 ( .A(\DataOut<6> ), .Y(n221) );
  INVX1 U319 ( .A(n221), .Y(n222) );
  INVX1 U320 ( .A(\DataOut<15> ), .Y(n223) );
  INVX1 U321 ( .A(n223), .Y(n224) );
  INVX1 U322 ( .A(\DataOut<7> ), .Y(n225) );
  INVX1 U323 ( .A(n225), .Y(n226) );
  INVX1 U324 ( .A(\DataOut<14> ), .Y(n227) );
  INVX1 U325 ( .A(n227), .Y(n228) );
  INVX1 U326 ( .A(\DataOut<11> ), .Y(n229) );
  INVX1 U327 ( .A(n229), .Y(n230) );
  INVX1 U328 ( .A(\DataOut<3> ), .Y(n231) );
  INVX1 U329 ( .A(n231), .Y(n232) );
  INVX1 U330 ( .A(\DataOut<5> ), .Y(n233) );
  INVX1 U331 ( .A(n233), .Y(n234) );
  AND2X2 U332 ( .A(n205), .B(n172), .Y(n236) );
  AND2X2 U333 ( .A(n449), .B(n209), .Y(n237) );
  INVX1 U334 ( .A(n237), .Y(n238) );
  AND2X2 U335 ( .A(\state<0> ), .B(net102842), .Y(n239) );
  INVX1 U336 ( .A(\next_state<1> ), .Y(n240) );
  INVX1 U337 ( .A(n240), .Y(n241) );
  INVX1 U338 ( .A(n242), .Y(n243) );
  INVX1 U339 ( .A(n244), .Y(n245) );
  AND2X1 U340 ( .A(\memDataOut<2> ), .B(net89037), .Y(n246) );
  INVX1 U341 ( .A(n246), .Y(n247) );
  INVX1 U342 ( .A(n248), .Y(n249) );
  INVX1 U343 ( .A(n250), .Y(n251) );
  AND2X1 U344 ( .A(\memDataOut<5> ), .B(net89037), .Y(n252) );
  INVX1 U345 ( .A(n252), .Y(n253) );
  AND2X1 U346 ( .A(\memDataOut<6> ), .B(net89037), .Y(n254) );
  INVX1 U347 ( .A(n254), .Y(n255) );
  AND2X1 U348 ( .A(\memDataOut<7> ), .B(net89037), .Y(n256) );
  INVX1 U349 ( .A(n256), .Y(n257) );
  AND2X1 U350 ( .A(\memDataOut<8> ), .B(net89037), .Y(n258) );
  INVX1 U351 ( .A(n258), .Y(n259) );
  AND2X1 U352 ( .A(\memDataOut<9> ), .B(net89037), .Y(n260) );
  INVX1 U353 ( .A(n260), .Y(n261) );
  AND2X1 U354 ( .A(\memDataOut<10> ), .B(net89037), .Y(n262) );
  INVX1 U355 ( .A(n262), .Y(n263) );
  AND2X1 U356 ( .A(\memDataOut<11> ), .B(net89037), .Y(n264) );
  INVX1 U357 ( .A(n264), .Y(n265) );
  AND2X1 U358 ( .A(\memDataOut<12> ), .B(net89037), .Y(n266) );
  INVX1 U359 ( .A(n266), .Y(n267) );
  AND2X1 U360 ( .A(\memDataOut<13> ), .B(net89037), .Y(n268) );
  INVX1 U361 ( .A(n268), .Y(n269) );
  AND2X1 U362 ( .A(\memDataOut<14> ), .B(net89037), .Y(n270) );
  INVX1 U363 ( .A(n270), .Y(n271) );
  AND2X1 U364 ( .A(\memDataOut<15> ), .B(net89037), .Y(n272) );
  INVX1 U365 ( .A(n272), .Y(n273) );
  OR2X2 U366 ( .A(n200), .B(n366), .Y(n274) );
  INVX1 U367 ( .A(n274), .Y(n275) );
  AND2X1 U368 ( .A(\DataIn<0> ), .B(n416), .Y(n276) );
  INVX1 U369 ( .A(n276), .Y(n277) );
  AND2X1 U370 ( .A(\DataIn<1> ), .B(n416), .Y(n278) );
  INVX1 U371 ( .A(n278), .Y(n279) );
  AND2X1 U372 ( .A(\DataIn<2> ), .B(n416), .Y(n280) );
  INVX1 U373 ( .A(n280), .Y(n281) );
  AND2X1 U374 ( .A(\DataIn<3> ), .B(n416), .Y(n282) );
  INVX1 U375 ( .A(n282), .Y(n283) );
  AND2X1 U376 ( .A(\DataIn<4> ), .B(n416), .Y(n284) );
  INVX1 U377 ( .A(n284), .Y(n285) );
  AND2X1 U378 ( .A(\DataIn<5> ), .B(n416), .Y(n286) );
  INVX1 U379 ( .A(n286), .Y(n287) );
  AND2X1 U380 ( .A(\DataIn<6> ), .B(n416), .Y(n288) );
  INVX1 U381 ( .A(n288), .Y(n289) );
  AND2X1 U382 ( .A(\DataIn<7> ), .B(n416), .Y(n290) );
  INVX1 U383 ( .A(n290), .Y(n291) );
  AND2X1 U384 ( .A(\DataIn<8> ), .B(n416), .Y(n292) );
  INVX1 U385 ( .A(n292), .Y(n293) );
  AND2X1 U386 ( .A(\DataIn<9> ), .B(n416), .Y(n294) );
  INVX1 U387 ( .A(n294), .Y(n295) );
  AND2X1 U388 ( .A(\DataIn<10> ), .B(n416), .Y(n296) );
  INVX1 U389 ( .A(n296), .Y(n297) );
  AND2X1 U390 ( .A(\DataIn<11> ), .B(n416), .Y(n298) );
  INVX1 U391 ( .A(n298), .Y(n299) );
  AND2X1 U392 ( .A(\DataIn<12> ), .B(n416), .Y(n300) );
  INVX1 U393 ( .A(n300), .Y(n301) );
  AND2X1 U394 ( .A(\DataIn<13> ), .B(n416), .Y(n302) );
  INVX1 U395 ( .A(n302), .Y(n303) );
  AND2X1 U396 ( .A(\DataIn<14> ), .B(n416), .Y(n304) );
  INVX1 U397 ( .A(n304), .Y(n305) );
  AND2X1 U398 ( .A(\DataIn<15> ), .B(n416), .Y(n306) );
  INVX1 U399 ( .A(n306), .Y(n307) );
  AND2X2 U400 ( .A(net95995), .B(net121828), .Y(n308) );
  INVX1 U401 ( .A(n308), .Y(n309) );
  OR2X1 U402 ( .A(net89031), .B(n353), .Y(n310) );
  INVX1 U403 ( .A(n310), .Y(n311) );
  OR2X1 U404 ( .A(n471), .B(n470), .Y(n312) );
  INVX1 U405 ( .A(n312), .Y(n313) );
  AND2X1 U406 ( .A(\cacheTagOut<1> ), .B(memWrite), .Y(n314) );
  INVX1 U407 ( .A(n314), .Y(n315) );
  AND2X1 U408 ( .A(\Addr<15> ), .B(n377), .Y(n316) );
  INVX1 U409 ( .A(n316), .Y(n317) );
  AND2X1 U410 ( .A(\Addr<14> ), .B(n377), .Y(n318) );
  INVX1 U411 ( .A(n318), .Y(n319) );
  AND2X1 U412 ( .A(\Addr<13> ), .B(n377), .Y(n320) );
  INVX1 U413 ( .A(n320), .Y(n321) );
  AND2X1 U414 ( .A(\Addr<12> ), .B(n377), .Y(n322) );
  INVX1 U415 ( .A(n322), .Y(n323) );
  AND2X1 U416 ( .A(\Addr<11> ), .B(n377), .Y(n324) );
  INVX1 U417 ( .A(n324), .Y(n325) );
  INVX1 U418 ( .A(n326), .Y(n327) );
  BUFX2 U419 ( .A(n454), .Y(n328) );
  AND2X1 U420 ( .A(n356), .B(n369), .Y(n329) );
  INVX1 U421 ( .A(n329), .Y(n330) );
  AND2X2 U422 ( .A(Stall), .B(n186), .Y(n331) );
  INVX1 U423 ( .A(n331), .Y(n332) );
  AND2X1 U424 ( .A(n452), .B(n366), .Y(n333) );
  INVX1 U425 ( .A(n333), .Y(n334) );
  AND2X1 U426 ( .A(n345), .B(net95995), .Y(Stall) );
  INVX1 U427 ( .A(n337), .Y(n338) );
  INVX1 U428 ( .A(n339), .Y(n340) );
  AND2X1 U429 ( .A(Wr), .B(n420), .Y(n341) );
  INVX1 U430 ( .A(n341), .Y(n342) );
  AND2X1 U431 ( .A(n201), .B(n380), .Y(n343) );
  INVX1 U432 ( .A(n343), .Y(n344) );
  AND2X2 U433 ( .A(net121753), .B(net121828), .Y(n345) );
  INVX1 U434 ( .A(n345), .Y(Done) );
  BUFX2 U435 ( .A(n459), .Y(n347) );
  INVX1 U436 ( .A(n345), .Y(n348) );
  OR2X1 U437 ( .A(n379), .B(n463), .Y(n349) );
  INVX1 U438 ( .A(n349), .Y(n350) );
  INVX1 U439 ( .A(cacheWrite), .Y(n351) );
  INVX1 U440 ( .A(n351), .Y(n352) );
  INVX1 U441 ( .A(n236), .Y(n353) );
  BUFX2 U442 ( .A(n207), .Y(n354) );
  INVX1 U443 ( .A(n354), .Y(n447) );
  AND2X1 U444 ( .A(mem_stall), .B(n358), .Y(n355) );
  INVX1 U445 ( .A(n355), .Y(n356) );
  AND2X2 U446 ( .A(n372), .B(n181), .Y(n357) );
  INVX1 U447 ( .A(n357), .Y(n358) );
  INVX1 U448 ( .A(n172), .Y(n359) );
  INVX1 U449 ( .A(n456), .Y(n360) );
  BUFX2 U450 ( .A(memAddr_2), .Y(n361) );
  INVX1 U451 ( .A(n220), .Y(n362) );
  INVX1 U452 ( .A(n220), .Y(n363) );
  AND2X2 U453 ( .A(n239), .B(n456), .Y(n364) );
  INVX1 U454 ( .A(n175), .Y(n366) );
  INVX1 U455 ( .A(n366), .Y(n367) );
  AND2X1 U456 ( .A(mem_stall), .B(n447), .Y(n368) );
  INVX1 U457 ( .A(n368), .Y(n369) );
  AND2X1 U458 ( .A(Wr), .B(n441), .Y(n370) );
  INVX1 U459 ( .A(n370), .Y(n371) );
  INVX1 U460 ( .A(n196), .Y(n469) );
  INVX1 U461 ( .A(n178), .Y(n372) );
  INVX1 U462 ( .A(n178), .Y(n373) );
  AND2X2 U463 ( .A(n417), .B(n424), .Y(n374) );
  INVX1 U464 ( .A(n374), .Y(n375) );
  AND2X1 U465 ( .A(net102793), .B(n379), .Y(n376) );
  INVX1 U466 ( .A(n376), .Y(n377) );
  OR2X2 U467 ( .A(memRead), .B(n332), .Y(n378) );
  INVX1 U468 ( .A(n378), .Y(n379) );
  INVX1 U469 ( .A(n176), .Y(n380) );
  AND2X1 U470 ( .A(n235), .B(net96034), .Y(n381) );
  INVX1 U471 ( .A(n381), .Y(n382) );
  INVX1 U472 ( .A(n383), .Y(n384) );
  INVX1 U473 ( .A(n385), .Y(n386) );
  INVX1 U474 ( .A(n387), .Y(n388) );
  INVX1 U475 ( .A(n389), .Y(n390) );
  INVX1 U476 ( .A(n391), .Y(n392) );
  INVX1 U477 ( .A(n393), .Y(n394) );
  INVX1 U478 ( .A(n395), .Y(n396) );
  INVX1 U479 ( .A(n397), .Y(n398) );
  INVX1 U480 ( .A(n399), .Y(n400) );
  INVX1 U481 ( .A(n401), .Y(n402) );
  INVX1 U482 ( .A(n403), .Y(n404) );
  INVX1 U483 ( .A(n405), .Y(n406) );
  INVX1 U484 ( .A(n407), .Y(n408) );
  INVX1 U485 ( .A(n409), .Y(n410) );
  INVX1 U486 ( .A(n411), .Y(n412) );
  INVX1 U487 ( .A(n413), .Y(n414) );
  AND2X2 U488 ( .A(net126586), .B(n379), .Y(n415) );
  INVX1 U489 ( .A(n415), .Y(n416) );
  AND2X2 U490 ( .A(net102834), .B(net89137), .Y(n417) );
  INVX1 U491 ( .A(\state<0> ), .Y(net89137) );
  NAND3X1 U492 ( .A(net121261), .B(net121272), .C(net89099), .Y(n418) );
  INVX1 U493 ( .A(n418), .Y(n456) );
  INVX2 U494 ( .A(\Addr<5> ), .Y(n429) );
  BUFX2 U495 ( .A(\Addr<3> ), .Y(n419) );
  INVX1 U496 ( .A(\state<2> ), .Y(net102841) );
  INVX1 U497 ( .A(net102841), .Y(net102842) );
  INVX1 U498 ( .A(net89119), .Y(net102834) );
  INVX1 U499 ( .A(n150), .Y(n420) );
  INVX1 U500 ( .A(n420), .Y(n421) );
  INVX1 U501 ( .A(net89127), .Y(net89098) );
  INVX1 U502 ( .A(\state<2> ), .Y(net89119) );
  BUFX2 U503 ( .A(net95788), .Y(net102793) );
  INVX1 U504 ( .A(n199), .Y(n441) );
  INVX1 U505 ( .A(n427), .Y(n422) );
  INVX1 U506 ( .A(dirty), .Y(n449) );
  NOR3X1 U507 ( .A(n176), .B(n358), .C(n374), .Y(n423) );
  INVX8 U508 ( .A(n423), .Y(memRead) );
  INVX1 U509 ( .A(net130129), .Y(net102554) );
  INVX1 U510 ( .A(n360), .Y(n424) );
  INVX1 U511 ( .A(net89031), .Y(net96034) );
  INVX1 U512 ( .A(net130115), .Y(net95941) );
  INVX1 U513 ( .A(\Addr<4> ), .Y(n427) );
  INVX1 U514 ( .A(net102793), .Y(net89037) );
  AND2X2 U515 ( .A(n365), .B(n140), .Y(net89083) );
  INVX1 U516 ( .A(n365), .Y(n470) );
  INVX1 U517 ( .A(net126586), .Y(memWrite) );
  AND2X2 U518 ( .A(n149), .B(n198), .Y(net95739) );
  INVX1 U519 ( .A(net95739), .Y(net89031) );
  INVX8 U520 ( .A(n426), .Y(n425) );
  INVX8 U521 ( .A(n429), .Y(n428) );
  INVX8 U522 ( .A(n431), .Y(n430) );
  INVX8 U523 ( .A(n433), .Y(n432) );
  INVX8 U524 ( .A(n435), .Y(n434) );
  NAND3X1 U525 ( .A(\state<1> ), .B(\state<3> ), .C(net89086), .Y(n440) );
  NAND2X1 U526 ( .A(net102834), .B(net89137), .Y(n442) );
  MUX2X1 U527 ( .B(n447), .A(n359), .S(mem_stall), .Y(n445) );
  NOR2X1 U528 ( .A(net121256), .B(net95941), .Y(n443) );
  NAND3X1 U529 ( .A(net102554), .B(n417), .C(n443), .Y(n455) );
  NAND3X1 U530 ( .A(\state<3> ), .B(net130138), .C(net130115), .Y(n444) );
  NAND3X1 U531 ( .A(n371), .B(n445), .C(net126590), .Y(n467) );
  NAND2X1 U532 ( .A(net130129), .B(n177), .Y(net89127) );
  OAI21X1 U533 ( .A(n372), .B(mem_stall), .C(n369), .Y(n448) );
  NOR3X1 U534 ( .A(n208), .B(n344), .C(n448), .Y(n451) );
  AOI21X1 U535 ( .A(hit), .B(valid), .C(n421), .Y(n450) );
  NOR3X1 U536 ( .A(\state<3> ), .B(net129930), .C(net129949), .Y(n453) );
  NAND3X1 U537 ( .A(n172), .B(n365), .C(n371), .Y(n454) );
  NAND3X1 U538 ( .A(n334), .B(n338), .C(n340), .Y(\next_state<1> ) );
  MUX2X1 U539 ( .B(n235), .A(n367), .S(mem_stall), .Y(n460) );
  OAI21X1 U540 ( .A(Wr), .B(Rd), .C(n309), .Y(n457) );
  NAND3X1 U541 ( .A(n458), .B(n457), .C(n356), .Y(n459) );
  NOR3X1 U542 ( .A(n368), .B(n460), .C(n347), .Y(n461) );
  NAND3X1 U543 ( .A(n461), .B(n203), .C(n238), .Y(\next_state<0> ) );
  NAND3X1 U544 ( .A(n363), .B(net102793), .C(n342), .Y(cacheWrite) );
  OAI21X1 U545 ( .A(n379), .B(n464), .C(n311), .Y(\cacheAddr<1> ) );
  OAI21X1 U546 ( .A(n379), .B(n466), .C(n336), .Y(\cacheAddr<2> ) );
  OAI21X1 U547 ( .A(n199), .B(Wr), .C(n363), .Y(\next_state<4> ) );
  NOR3X1 U548 ( .A(n208), .B(n468), .C(n469), .Y(n472) );
  MUX2X1 U549 ( .B(n181), .A(n373), .S(mem_stall), .Y(n471) );
  NAND3X1 U550 ( .A(n380), .B(n336), .C(n373), .Y(memAddr_2) );
endmodule

