
module fulladder_1_15 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2, n3, n4, n5, n7, n8, n9;

  AND2X2 U1 ( .A(n7), .B(B), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  AND2X2 U3 ( .A(A), .B(n8), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  AND2X2 U5 ( .A(n4), .B(n2), .Y(n5) );
  INVX1 U6 ( .A(n5), .Y(p) );
  INVX1 U7 ( .A(A), .Y(n7) );
  INVX1 U8 ( .A(B), .Y(n8) );
  INVX1 U9 ( .A(p), .Y(n9) );
  XNOR2X1 U10 ( .A(Cin), .B(n9), .Y(S) );
  AND2X2 U11 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_14 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n3, n4, n5, n7, n8, n9;

  INVX1 U1 ( .A(B), .Y(n9) );
  INVX1 U2 ( .A(n9), .Y(n1) );
  AND2X2 U3 ( .A(n1), .B(A), .Y(g) );
  INVX1 U4 ( .A(g), .Y(n3) );
  AND2X2 U5 ( .A(n9), .B(n8), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(n5) );
  AND2X2 U7 ( .A(n3), .B(n5), .Y(p) );
  INVX1 U8 ( .A(p), .Y(n7) );
  INVX1 U9 ( .A(A), .Y(n8) );
  XNOR2X1 U10 ( .A(Cin), .B(n7), .Y(S) );
endmodule


module fulladder_1_13 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2;

  INVX2 U1 ( .A(n2), .Y(p) );
  XOR2X1 U2 ( .A(Cin), .B(p), .Y(S) );
  XOR2X1 U3 ( .A(n1), .B(B), .Y(n2) );
  INVX1 U4 ( .A(A), .Y(n1) );
  AND2X2 U5 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_12 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n1), .Y(p) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_3 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40;

  INVX1 U1 ( .A(\g<0> ), .Y(n35) );
  INVX1 U2 ( .A(\g<1> ), .Y(n36) );
  AND2X1 U3 ( .A(\p<1> ), .B(\g<0> ), .Y(n11) );
  AND2X1 U4 ( .A(n22), .B(n25), .Y(n15) );
  INVX1 U5 ( .A(\g<3> ), .Y(n38) );
  AND2X2 U6 ( .A(Cin), .B(n24), .Y(n17) );
  OR2X2 U7 ( .A(n28), .B(n39), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(pg) );
  OR2X2 U9 ( .A(\g<2> ), .B(\g<1> ), .Y(n3) );
  INVX1 U10 ( .A(n3), .Y(n4) );
  AND2X2 U11 ( .A(n33), .B(n19), .Y(n5) );
  INVX1 U12 ( .A(n5), .Y(n6) );
  AND2X2 U13 ( .A(n4), .B(n12), .Y(n7) );
  INVX1 U14 ( .A(n7), .Y(n8) );
  AND2X2 U15 ( .A(n29), .B(n30), .Y(n9) );
  INVX1 U16 ( .A(n9), .Y(n10) );
  INVX1 U17 ( .A(n11), .Y(n12) );
  AND2X2 U18 ( .A(n8), .B(n10), .Y(n13) );
  INVX1 U19 ( .A(n13), .Y(n14) );
  INVX1 U20 ( .A(n15), .Y(n16) );
  INVX1 U21 ( .A(n17), .Y(n18) );
  INVX1 U22 ( .A(n17), .Y(n19) );
  AND2X2 U23 ( .A(n35), .B(n18), .Y(n20) );
  INVX1 U24 ( .A(n20), .Y(\c<0> ) );
  INVX1 U25 ( .A(n20), .Y(n22) );
  BUFX2 U26 ( .A(\c<2> ), .Y(n23) );
  BUFX2 U27 ( .A(\p<0> ), .Y(n24) );
  BUFX2 U28 ( .A(\p<1> ), .Y(n25) );
  BUFX2 U29 ( .A(n37), .Y(n26) );
  INVX1 U30 ( .A(n34), .Y(n27) );
  INVX1 U31 ( .A(n27), .Y(n28) );
  OAI21X1 U32 ( .A(n30), .B(n16), .C(n26), .Y(\c<2> ) );
  INVX1 U33 ( .A(\g<2> ), .Y(n29) );
  INVX1 U34 ( .A(\p<2> ), .Y(n30) );
  INVX1 U35 ( .A(\p<3> ), .Y(n39) );
  INVX1 U36 ( .A(n23), .Y(n40) );
  AND2X2 U37 ( .A(n6), .B(n31), .Y(\c<1> ) );
  OR2X2 U38 ( .A(n32), .B(n25), .Y(n31) );
  INVX1 U39 ( .A(n36), .Y(n32) );
  AND2X2 U40 ( .A(n35), .B(n36), .Y(n33) );
  OAI21X1 U41 ( .A(n39), .B(n14), .C(n38), .Y(gg) );
  NAND3X1 U42 ( .A(\p<1> ), .B(\p<0> ), .C(\p<2> ), .Y(n34) );
  AOI21X1 U43 ( .A(\g<1> ), .B(\p<2> ), .C(\g<2> ), .Y(n37) );
  OAI21X1 U44 ( .A(n39), .B(n40), .C(n38), .Y(\c<3> ) );
endmodule


module fulladder_1_11 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n2;

  XNOR2X1 U1 ( .A(B), .B(A), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(B), .B(A), .Y(g) );
endmodule


module fulladder_1_10 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n3;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  BUFX2 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(p) );
  XNOR2X1 U4 ( .A(B), .B(A), .Y(n3) );
  AND2X2 U5 ( .A(B), .B(A), .Y(g) );
endmodule


module fulladder_1_9 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2, n3, n5, n6, n7;

  INVX1 U1 ( .A(B), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  BUFX2 U3 ( .A(n7), .Y(n3) );
  INVX1 U4 ( .A(n6), .Y(n5) );
  XNOR2X1 U5 ( .A(Cin), .B(n3), .Y(S) );
  INVX1 U6 ( .A(n7), .Y(p) );
  XNOR2X1 U7 ( .A(n2), .B(n5), .Y(n7) );
  INVX2 U8 ( .A(A), .Y(n6) );
  AND2X2 U9 ( .A(B), .B(A), .Y(g) );
endmodule


module fulladder_1_8 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2, n3, n4, n6;

  INVX1 U1 ( .A(n6), .Y(p) );
  INVX1 U2 ( .A(B), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  BUFX2 U4 ( .A(Cin), .Y(n3) );
  BUFX2 U5 ( .A(p), .Y(n4) );
  XNOR2X1 U6 ( .A(n2), .B(A), .Y(n6) );
  XOR2X1 U7 ( .A(n3), .B(n4), .Y(S) );
  AND2X2 U8 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_2 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n2, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47;

  AND2X1 U1 ( .A(n11), .B(\p<1> ), .Y(n19) );
  INVX1 U2 ( .A(\g<0> ), .Y(n43) );
  INVX1 U3 ( .A(\g<1> ), .Y(n44) );
  INVX1 U4 ( .A(n45), .Y(n1) );
  INVX1 U5 ( .A(\g<3> ), .Y(n45) );
  OR2X2 U6 ( .A(n14), .B(n41), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(gg) );
  INVX1 U8 ( .A(n10), .Y(\c<0> ) );
  OR2X2 U9 ( .A(n1), .B(n32), .Y(n5) );
  OR2X2 U10 ( .A(n16), .B(n18), .Y(n6) );
  INVX1 U11 ( .A(n6), .Y(pg) );
  AND2X2 U12 ( .A(n36), .B(n24), .Y(n8) );
  INVX1 U13 ( .A(n8), .Y(n9) );
  AND2X2 U14 ( .A(n43), .B(n12), .Y(n10) );
  INVX1 U15 ( .A(n10), .Y(n11) );
  INVX1 U16 ( .A(n23), .Y(n12) );
  OR2X2 U17 ( .A(n33), .B(n21), .Y(n13) );
  INVX1 U18 ( .A(n13), .Y(n14) );
  AND2X2 U19 ( .A(\p<0> ), .B(\p<1> ), .Y(n15) );
  INVX1 U20 ( .A(n15), .Y(n16) );
  AND2X2 U21 ( .A(\p<2> ), .B(\p<3> ), .Y(n17) );
  INVX1 U22 ( .A(n17), .Y(n18) );
  INVX1 U23 ( .A(n19), .Y(n20) );
  OR2X2 U24 ( .A(\g<2> ), .B(\g<3> ), .Y(n21) );
  INVX1 U25 ( .A(n21), .Y(n22) );
  AND2X2 U26 ( .A(Cin), .B(n30), .Y(n23) );
  INVX1 U27 ( .A(n23), .Y(n24) );
  OR2X2 U28 ( .A(n39), .B(\g<2> ), .Y(n25) );
  INVX1 U29 ( .A(n25), .Y(n26) );
  OR2X2 U30 ( .A(\g<2> ), .B(\g<1> ), .Y(n27) );
  INVX1 U31 ( .A(n27), .Y(n28) );
  BUFX2 U32 ( .A(n47), .Y(n29) );
  BUFX2 U33 ( .A(\p<0> ), .Y(n30) );
  INVX1 U34 ( .A(\p<3> ), .Y(n31) );
  INVX1 U35 ( .A(n31), .Y(n32) );
  INVX1 U36 ( .A(n42), .Y(n33) );
  AND2X2 U37 ( .A(n9), .B(n34), .Y(\c<1> ) );
  OR2X2 U38 ( .A(n35), .B(\p<1> ), .Y(n34) );
  INVX1 U39 ( .A(n44), .Y(n35) );
  AND2X2 U40 ( .A(n43), .B(n44), .Y(n36) );
  BUFX2 U41 ( .A(\c<1> ), .Y(n37) );
  INVX1 U42 ( .A(\p<2> ), .Y(n38) );
  INVX1 U43 ( .A(n38), .Y(n39) );
  INVX1 U44 ( .A(n22), .Y(n40) );
  INVX1 U45 ( .A(n32), .Y(n46) );
  AOI21X1 U46 ( .A(\g<0> ), .B(\p<1> ), .C(\g<1> ), .Y(n42) );
  OAI21X1 U47 ( .A(n39), .B(n40), .C(n5), .Y(n41) );
  AOI21X1 U48 ( .A(n28), .B(n20), .C(n26), .Y(\c<2> ) );
  AOI21X1 U49 ( .A(n39), .B(n37), .C(\g<2> ), .Y(n47) );
  OAI21X1 U50 ( .A(n29), .B(n46), .C(n45), .Y(\c<3> ) );
endmodule


module fulladder_1_7 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  INVX2 U1 ( .A(n1), .Y(p) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_6 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2;

  BUFX2 U1 ( .A(n2), .Y(n1) );
  XNOR2X1 U2 ( .A(Cin), .B(n1), .Y(S) );
  INVX1 U3 ( .A(n2), .Y(p) );
  XNOR2X1 U4 ( .A(B), .B(A), .Y(n2) );
  AND2X2 U5 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_5 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(Cin), .B(n1), .Y(S) );
  XNOR2X1 U2 ( .A(B), .B(A), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(p) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_4 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2, n3;

  INVX1 U1 ( .A(n3), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(p) );
  XNOR2X1 U4 ( .A(Cin), .B(n2), .Y(S) );
  XNOR2X1 U5 ( .A(B), .B(A), .Y(n3) );
  AND2X2 U6 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_1 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26;

  INVX1 U1 ( .A(\g<0> ), .Y(n20) );
  OR2X2 U2 ( .A(n9), .B(n11), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(pg) );
  OR2X2 U4 ( .A(\g<1> ), .B(\g<2> ), .Y(n3) );
  AND2X2 U5 ( .A(Cin), .B(\p<0> ), .Y(n4) );
  INVX1 U6 ( .A(n4), .Y(n5) );
  AND2X2 U7 ( .A(\p<2> ), .B(\c<1> ), .Y(n6) );
  INVX1 U8 ( .A(n6), .Y(n7) );
  AND2X2 U9 ( .A(\p<0> ), .B(\p<1> ), .Y(n8) );
  INVX1 U10 ( .A(n8), .Y(n9) );
  AND2X2 U11 ( .A(\p<3> ), .B(\p<2> ), .Y(n10) );
  INVX1 U12 ( .A(n10), .Y(n11) );
  AND2X2 U13 ( .A(\p<1> ), .B(\g<0> ), .Y(n12) );
  INVX1 U14 ( .A(n12), .Y(n13) );
  OR2X2 U15 ( .A(\g<3> ), .B(n3), .Y(n14) );
  INVX1 U16 ( .A(n14), .Y(n15) );
  AND2X2 U17 ( .A(n23), .B(n7), .Y(n16) );
  INVX1 U18 ( .A(n16), .Y(\c<2> ) );
  INVX1 U19 ( .A(\g<3> ), .Y(n24) );
  INVX1 U20 ( .A(\g<1> ), .Y(n21) );
  INVX1 U21 ( .A(\p<3> ), .Y(n25) );
  INVX1 U22 ( .A(\p<1> ), .Y(n22) );
  INVX1 U23 ( .A(\g<2> ), .Y(n23) );
  AND2X2 U24 ( .A(n20), .B(n5), .Y(n18) );
  INVX1 U25 ( .A(n18), .Y(\c<0> ) );
  INVX1 U26 ( .A(\c<2> ), .Y(n26) );
  OAI21X1 U27 ( .A(\g<2> ), .B(\p<2> ), .C(\p<3> ), .Y(n19) );
  AOI22X1 U28 ( .A(n15), .B(n13), .C(n24), .D(n19), .Y(gg) );
  OAI21X1 U29 ( .A(n18), .B(n22), .C(n21), .Y(\c<1> ) );
  OAI21X1 U30 ( .A(n26), .B(n25), .C(n24), .Y(\c<3> ) );
endmodule


module fulladder_1_3 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2;

  INVX1 U1 ( .A(Cin), .Y(n2) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(p) );
  XNOR2X1 U4 ( .A(p), .B(n2), .Y(S) );
  AND2X2 U5 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_2 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n3, n4, n5, n6, n7, n8;

  INVX1 U1 ( .A(B), .Y(n1) );
  AND2X2 U2 ( .A(n5), .B(n4), .Y(p) );
  AND2X2 U3 ( .A(n6), .B(n1), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n4) );
  INVX1 U5 ( .A(g), .Y(n5) );
  INVX1 U6 ( .A(A), .Y(n6) );
  INVX1 U7 ( .A(n1), .Y(n7) );
  BUFX2 U8 ( .A(p), .Y(n8) );
  XOR2X1 U9 ( .A(Cin), .B(n8), .Y(S) );
  AND2X2 U10 ( .A(A), .B(n7), .Y(g) );
endmodule


module fulladder_1_1 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_0 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  INVX4 U1 ( .A(n1), .Y(p) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_0 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33;

  INVX1 U1 ( .A(\g<2> ), .Y(n30) );
  AND2X2 U2 ( .A(n12), .B(n5), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(gg) );
  OR2X2 U4 ( .A(n14), .B(n16), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(pg) );
  AND2X2 U6 ( .A(n31), .B(n11), .Y(n5) );
  AND2X2 U7 ( .A(\g<0> ), .B(\p<1> ), .Y(n6) );
  INVX1 U8 ( .A(n6), .Y(n7) );
  AND2X2 U9 ( .A(\p<2> ), .B(\c<1> ), .Y(n8) );
  INVX1 U10 ( .A(n8), .Y(n9) );
  AND2X2 U11 ( .A(\p<3> ), .B(\g<2> ), .Y(n10) );
  INVX1 U12 ( .A(n10), .Y(n11) );
  BUFX2 U13 ( .A(n26), .Y(n12) );
  AND2X2 U14 ( .A(\p<0> ), .B(n25), .Y(n13) );
  INVX1 U15 ( .A(n13), .Y(n14) );
  AND2X2 U16 ( .A(\p<2> ), .B(\p<3> ), .Y(n15) );
  INVX1 U17 ( .A(n15), .Y(n16) );
  AND2X2 U18 ( .A(n7), .B(n28), .Y(n17) );
  INVX1 U19 ( .A(n17), .Y(n18) );
  AND2X2 U20 ( .A(n30), .B(n9), .Y(n19) );
  INVX1 U21 ( .A(n19), .Y(\c<2> ) );
  INVX1 U22 ( .A(n19), .Y(n21) );
  INVX1 U23 ( .A(n24), .Y(\c<1> ) );
  INVX1 U24 ( .A(n21), .Y(n33) );
  OAI21X1 U25 ( .A(n22), .B(n23), .C(n27), .Y(\c<0> ) );
  INVX1 U26 ( .A(Cin), .Y(n22) );
  INVX1 U27 ( .A(\p<0> ), .Y(n23) );
  INVX1 U28 ( .A(\g<0> ), .Y(n27) );
  AOI21X1 U29 ( .A(\c<0> ), .B(n25), .C(\g<1> ), .Y(n24) );
  INVX1 U30 ( .A(\g<1> ), .Y(n28) );
  INVX1 U31 ( .A(n29), .Y(n25) );
  INVX1 U32 ( .A(\p<3> ), .Y(n32) );
  INVX1 U33 ( .A(\p<1> ), .Y(n29) );
  INVX1 U34 ( .A(\g<3> ), .Y(n31) );
  NAND3X1 U35 ( .A(\p<3> ), .B(\p<2> ), .C(n18), .Y(n26) );
  OAI21X1 U36 ( .A(n33), .B(n32), .C(n31), .Y(\c<3> ) );
endmodule


module fulladder_1_47 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(g) );
  INVX1 U2 ( .A(n1), .Y(p) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(p), .Y(S) );
endmodule


module fulladder_1_46 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;


  AND2X1 U1 ( .A(A), .B(B), .Y(g) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
endmodule


module fulladder_1_45 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;


  AND2X1 U1 ( .A(A), .B(B), .Y(g) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
endmodule


module fulladder_1_44 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;


  AND2X1 U1 ( .A(A), .B(B), .Y(g) );
  XOR2X1 U2 ( .A(A), .B(B), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
endmodule


module groupcla_12 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n2, n3, n4, n5, n7, n8, n10, n11, n12, n13, n14, n15, n16, n18,
         n19, n20, n21, n22, n24, n25, n26, n27;

  NOR3X1 U8 ( .A(n16), .B(n24), .C(n26), .Y(pg) );
  OAI21X1 U10 ( .A(n14), .B(n26), .C(n25), .Y(gg) );
  AOI21X1 U11 ( .A(\p<2> ), .B(n13), .C(\g<2> ), .Y(n27) );
  INVX1 U1 ( .A(\g<0> ), .Y(n18) );
  INVX1 U2 ( .A(\p<1> ), .Y(n19) );
  INVX1 U3 ( .A(\g<1> ), .Y(n22) );
  INVX1 U4 ( .A(\g<2> ), .Y(n20) );
  AND2X1 U5 ( .A(n22), .B(n11), .Y(n12) );
  INVX1 U6 ( .A(\p<2> ), .Y(n24) );
  INVX1 U7 ( .A(\g<3> ), .Y(n25) );
  INVX1 U9 ( .A(\p<3> ), .Y(n26) );
  AND2X2 U12 ( .A(\p<0> ), .B(Cin), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  AND2X2 U14 ( .A(\p<2> ), .B(\c<1> ), .Y(n3) );
  INVX1 U15 ( .A(n3), .Y(n4) );
  AND2X2 U16 ( .A(n20), .B(n4), .Y(n5) );
  INVX1 U17 ( .A(n5), .Y(\c<2> ) );
  INVX1 U18 ( .A(n5), .Y(n7) );
  AND2X2 U19 ( .A(n18), .B(n2), .Y(n8) );
  AND2X1 U20 ( .A(\p<1> ), .B(\g<0> ), .Y(n10) );
  INVX1 U21 ( .A(n10), .Y(n11) );
  INVX1 U22 ( .A(n12), .Y(n13) );
  BUFX2 U23 ( .A(n27), .Y(n14) );
  AND2X1 U24 ( .A(\p<1> ), .B(\p<0> ), .Y(n15) );
  INVX1 U25 ( .A(n15), .Y(n16) );
  INVX1 U26 ( .A(n8), .Y(\c<0> ) );
  INVX1 U27 ( .A(n7), .Y(n21) );
  OAI21X1 U28 ( .A(n8), .B(n19), .C(n22), .Y(\c<1> ) );
  OAI21X1 U29 ( .A(n21), .B(n26), .C(n25), .Y(\c<3> ) );
endmodule


module fulladder_1_43 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(g) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(p) );
  XOR2X1 U4 ( .A(Cin), .B(p), .Y(S) );
endmodule


module fulladder_1_42 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(g) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(p) );
  XOR2X1 U4 ( .A(Cin), .B(p), .Y(S) );
endmodule


module fulladder_1_41 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(g) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(p) );
  XOR2X1 U4 ( .A(Cin), .B(p), .Y(S) );
endmodule


module fulladder_1_40 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(g) );
  INVX1 U2 ( .A(n1), .Y(p) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XOR2X1 U4 ( .A(Cin), .B(p), .Y(S) );
endmodule


module groupcla_11 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n13, n14, n16, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33;

  NOR3X1 U8 ( .A(n25), .B(n30), .C(n32), .Y(pg) );
  OAI21X1 U10 ( .A(n23), .B(n32), .C(n31), .Y(gg) );
  AOI21X1 U11 ( .A(\p<2> ), .B(n20), .C(\g<2> ), .Y(n33) );
  INVX1 U1 ( .A(\g<2> ), .Y(n27) );
  INVX1 U2 ( .A(\p<3> ), .Y(n32) );
  INVX1 U3 ( .A(\g<1> ), .Y(n29) );
  INVX1 U4 ( .A(\g<0> ), .Y(n26) );
  INVX1 U5 ( .A(\p<2> ), .Y(n30) );
  INVX1 U6 ( .A(n32), .Y(n28) );
  INVX1 U7 ( .A(\g<3> ), .Y(n31) );
  AND2X2 U9 ( .A(\p<0> ), .B(Cin), .Y(n1) );
  INVX1 U12 ( .A(n1), .Y(n2) );
  AND2X2 U13 ( .A(\p<1> ), .B(n11), .Y(n3) );
  INVX1 U14 ( .A(n3), .Y(n4) );
  AND2X2 U15 ( .A(\p<2> ), .B(n14), .Y(n5) );
  INVX1 U16 ( .A(n5), .Y(n6) );
  AND2X2 U17 ( .A(\p<1> ), .B(\g<0> ), .Y(n7) );
  INVX1 U18 ( .A(n7), .Y(n8) );
  AND2X2 U19 ( .A(n26), .B(n2), .Y(n10) );
  INVX1 U20 ( .A(n10), .Y(n11) );
  INVX1 U21 ( .A(n10), .Y(\c<0> ) );
  AND2X2 U22 ( .A(n29), .B(n4), .Y(n13) );
  INVX1 U23 ( .A(n13), .Y(n14) );
  INVX1 U24 ( .A(n13), .Y(\c<1> ) );
  AND2X2 U25 ( .A(n27), .B(n6), .Y(n16) );
  INVX1 U26 ( .A(n16), .Y(\c<2> ) );
  INVX1 U27 ( .A(n16), .Y(n18) );
  AND2X2 U28 ( .A(n29), .B(n8), .Y(n19) );
  INVX1 U29 ( .A(n19), .Y(n20) );
  AND2X1 U30 ( .A(n28), .B(n18), .Y(n21) );
  INVX1 U31 ( .A(n21), .Y(n22) );
  BUFX2 U32 ( .A(n33), .Y(n23) );
  AND2X1 U33 ( .A(\p<1> ), .B(\p<0> ), .Y(n24) );
  INVX1 U34 ( .A(n24), .Y(n25) );
  NAND2X1 U35 ( .A(n31), .B(n22), .Y(\c<3> ) );
endmodule


module fulladder_1_39 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_38 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_37 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  AND2X1 U1 ( .A(A), .B(B), .Y(g) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(p) );
  XOR2X1 U4 ( .A(Cin), .B(p), .Y(S) );
endmodule


module fulladder_1_36 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_10 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  INVX1 U1 ( .A(\g<1> ), .Y(n25) );
  INVX1 U2 ( .A(\p<1> ), .Y(n26) );
  INVX1 U3 ( .A(\g<2> ), .Y(n27) );
  INVX1 U4 ( .A(\g<3> ), .Y(n28) );
  INVX1 U5 ( .A(\p<2> ), .Y(n21) );
  INVX1 U6 ( .A(\g<0> ), .Y(n24) );
  INVX1 U7 ( .A(\p<3> ), .Y(n29) );
  AND2X2 U8 ( .A(n28), .B(n10), .Y(n1) );
  INVX1 U9 ( .A(n1), .Y(gg) );
  OR2X2 U10 ( .A(n12), .B(n20), .Y(n3) );
  INVX1 U11 ( .A(n3), .Y(pg) );
  AND2X2 U12 ( .A(Cin), .B(\p<0> ), .Y(n5) );
  INVX1 U13 ( .A(n5), .Y(n6) );
  AND2X2 U14 ( .A(\p<2> ), .B(\c<1> ), .Y(n7) );
  INVX1 U15 ( .A(n7), .Y(n8) );
  AND2X2 U16 ( .A(\p<3> ), .B(n23), .Y(n9) );
  INVX1 U17 ( .A(n9), .Y(n10) );
  AND2X2 U18 ( .A(\p<0> ), .B(\p<1> ), .Y(n11) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  BUFX2 U20 ( .A(n22), .Y(n13) );
  AND2X2 U21 ( .A(n27), .B(n8), .Y(n14) );
  INVX1 U22 ( .A(n14), .Y(\c<2> ) );
  INVX1 U23 ( .A(n14), .Y(n16) );
  AND2X2 U24 ( .A(n24), .B(n6), .Y(n17) );
  INVX1 U25 ( .A(n17), .Y(\c<0> ) );
  AND2X2 U26 ( .A(\p<3> ), .B(\p<2> ), .Y(n19) );
  INVX1 U27 ( .A(n19), .Y(n20) );
  INVX1 U28 ( .A(n16), .Y(n30) );
  AOI21X1 U29 ( .A(\p<1> ), .B(\g<0> ), .C(\g<1> ), .Y(n22) );
  OAI21X1 U30 ( .A(n13), .B(n21), .C(n27), .Y(n23) );
  OAI21X1 U31 ( .A(n17), .B(n26), .C(n25), .Y(\c<1> ) );
  OAI21X1 U32 ( .A(n30), .B(n29), .C(n28), .Y(\c<3> ) );
endmodule


module fulladder_1_35 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2;

  INVX1 U1 ( .A(Cin), .Y(n2) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(p) );
  XNOR2X1 U4 ( .A(p), .B(n2), .Y(S) );
  AND2X2 U5 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_34 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_33 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_32 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_9 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  INVX1 U1 ( .A(\g<1> ), .Y(n23) );
  INVX1 U2 ( .A(\p<1> ), .Y(n24) );
  INVX1 U3 ( .A(\p<2> ), .Y(n18) );
  INVX1 U4 ( .A(\g<0> ), .Y(n22) );
  INVX1 U5 ( .A(\p<0> ), .Y(n21) );
  INVX1 U6 ( .A(\g<3> ), .Y(n26) );
  INVX1 U7 ( .A(\p<3> ), .Y(n27) );
  INVX1 U8 ( .A(\g<2> ), .Y(n25) );
  AND2X2 U9 ( .A(n26), .B(n8), .Y(n1) );
  INVX1 U10 ( .A(n1), .Y(gg) );
  AND2X2 U11 ( .A(Cin), .B(\p<0> ), .Y(n3) );
  INVX1 U12 ( .A(n3), .Y(n4) );
  AND2X2 U13 ( .A(\p<2> ), .B(\c<1> ), .Y(n5) );
  INVX1 U14 ( .A(n5), .Y(n6) );
  AND2X2 U15 ( .A(\p<3> ), .B(n20), .Y(n7) );
  INVX1 U16 ( .A(n7), .Y(n8) );
  AND2X2 U17 ( .A(\p<3> ), .B(\p<2> ), .Y(n9) );
  INVX1 U18 ( .A(n9), .Y(n10) );
  AND2X2 U19 ( .A(n25), .B(n6), .Y(n11) );
  INVX1 U20 ( .A(n11), .Y(\c<2> ) );
  INVX1 U21 ( .A(n11), .Y(n13) );
  AND2X2 U22 ( .A(n22), .B(n4), .Y(n14) );
  INVX1 U23 ( .A(n14), .Y(\c<0> ) );
  INVX1 U24 ( .A(n19), .Y(n16) );
  INVX1 U25 ( .A(n16), .Y(n17) );
  INVX1 U26 ( .A(n13), .Y(n28) );
  AOI21X1 U27 ( .A(\p<1> ), .B(\g<0> ), .C(\g<1> ), .Y(n19) );
  OAI21X1 U28 ( .A(n17), .B(n18), .C(n25), .Y(n20) );
  NOR3X1 U29 ( .A(n10), .B(n24), .C(n21), .Y(pg) );
  OAI21X1 U30 ( .A(n14), .B(n24), .C(n23), .Y(\c<1> ) );
  OAI21X1 U31 ( .A(n28), .B(n27), .C(n26), .Y(\c<3> ) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(n1), .B(rst), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U3 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n1) );
  NOR2X1 U4 ( .A(n1), .B(rst), .Y(N3) );
endmodule


module shifter_1 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), .op({\op<2> , \op<1> , \op<0> }), 
        sh, .out({\out<15> , \out<14> , \out<13> , \out<12> , \out<11> , 
        \out<10> , \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , 
        \out<3> , \out<2> , \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , \op<2> , \op<1> , \op<0> , sh;
  output \out<15> , \out<14> , \out<13> , \out<12> , \out<11> , \out<10> ,
         \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> ,
         \out<2> , \out<1> , \out<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142;

  INVX1 U2 ( .A(\op<2> ), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n100), .Y(n3) );
  NOR3X1 U5 ( .A(n131), .B(n141), .C(n127), .Y(n4) );
  INVX2 U6 ( .A(n4), .Y(n128) );
  INVX4 U7 ( .A(sh), .Y(n131) );
  INVX2 U8 ( .A(\in<15> ), .Y(n141) );
  INVX1 U9 ( .A(n122), .Y(n5) );
  OR2X2 U10 ( .A(n35), .B(n36), .Y(n6) );
  INVX1 U11 ( .A(n122), .Y(n7) );
  INVX1 U12 ( .A(n100), .Y(n8) );
  INVX1 U13 ( .A(n99), .Y(n140) );
  INVX1 U14 ( .A(n124), .Y(n9) );
  INVX1 U15 ( .A(n123), .Y(n10) );
  INVX1 U16 ( .A(n136), .Y(n11) );
  INVX1 U17 ( .A(n11), .Y(n12) );
  AND2X2 U18 ( .A(n109), .B(n34), .Y(n13) );
  INVX1 U19 ( .A(n13), .Y(\out<0> ) );
  OR2X2 U20 ( .A(n128), .B(\op<1> ), .Y(n15) );
  INVX1 U21 ( .A(n15), .Y(n16) );
  AND2X2 U22 ( .A(\in<4> ), .B(n132), .Y(n17) );
  AND2X2 U23 ( .A(\in<3> ), .B(n133), .Y(n18) );
  INVX1 U24 ( .A(n18), .Y(n19) );
  AND2X2 U25 ( .A(\in<5> ), .B(n130), .Y(n20) );
  INVX1 U26 ( .A(n20), .Y(n21) );
  AND2X2 U27 ( .A(\in<6> ), .B(n133), .Y(n22) );
  INVX1 U28 ( .A(n22), .Y(n23) );
  AND2X2 U29 ( .A(\in<7> ), .B(n133), .Y(n24) );
  INVX1 U30 ( .A(n24), .Y(n25) );
  AND2X2 U31 ( .A(\in<8> ), .B(n133), .Y(n26) );
  INVX1 U32 ( .A(n26), .Y(n27) );
  AND2X2 U33 ( .A(\in<10> ), .B(n135), .Y(n28) );
  INVX1 U34 ( .A(n28), .Y(n29) );
  AND2X2 U35 ( .A(\in<12> ), .B(n137), .Y(n30) );
  INVX1 U36 ( .A(n30), .Y(n31) );
  AND2X2 U37 ( .A(\in<13> ), .B(n135), .Y(n32) );
  INVX1 U38 ( .A(n32), .Y(n33) );
  BUFX2 U39 ( .A(n129), .Y(n34) );
  AND2X2 U40 ( .A(n126), .B(\op<0> ), .Y(n35) );
  AND2X2 U41 ( .A(n122), .B(\op<2> ), .Y(n36) );
  AND2X2 U42 ( .A(\in<2> ), .B(n120), .Y(n37) );
  INVX1 U43 ( .A(n37), .Y(n38) );
  AND2X2 U44 ( .A(\in<3> ), .B(n140), .Y(n39) );
  INVX1 U45 ( .A(n39), .Y(n40) );
  AND2X2 U46 ( .A(\in<5> ), .B(n140), .Y(n41) );
  INVX1 U47 ( .A(n41), .Y(n42) );
  AND2X2 U48 ( .A(\in<6> ), .B(n140), .Y(n43) );
  INVX1 U49 ( .A(n43), .Y(n44) );
  AND2X2 U50 ( .A(\in<7> ), .B(n120), .Y(n45) );
  INVX1 U51 ( .A(n45), .Y(n46) );
  AND2X2 U52 ( .A(\in<8> ), .B(n8), .Y(n47) );
  INVX1 U53 ( .A(n47), .Y(n48) );
  AND2X2 U54 ( .A(\in<10> ), .B(n8), .Y(n49) );
  INVX1 U55 ( .A(n49), .Y(n50) );
  AND2X2 U56 ( .A(\in<11> ), .B(n120), .Y(n51) );
  INVX1 U57 ( .A(n51), .Y(n52) );
  AND2X2 U58 ( .A(\in<12> ), .B(n8), .Y(n53) );
  INVX1 U59 ( .A(n53), .Y(n54) );
  AND2X2 U60 ( .A(n136), .B(n103), .Y(n55) );
  INVX1 U61 ( .A(n55), .Y(n56) );
  AND2X2 U62 ( .A(\in<0> ), .B(sh), .Y(n57) );
  INVX1 U63 ( .A(n57), .Y(n58) );
  AND2X2 U64 ( .A(n134), .B(\in<2> ), .Y(n59) );
  INVX1 U65 ( .A(n59), .Y(n60) );
  AND2X2 U66 ( .A(\in<1> ), .B(n3), .Y(n61) );
  INVX1 U67 ( .A(n61), .Y(n62) );
  AND2X2 U68 ( .A(\in<6> ), .B(n139), .Y(n63) );
  INVX1 U69 ( .A(n63), .Y(n64) );
  AND2X2 U70 ( .A(\in<8> ), .B(n134), .Y(n65) );
  INVX1 U71 ( .A(n65), .Y(n66) );
  AND2X2 U72 ( .A(\in<9> ), .B(n3), .Y(n67) );
  INVX1 U73 ( .A(n67), .Y(n68) );
  AND2X2 U74 ( .A(\in<12> ), .B(n138), .Y(n69) );
  INVX1 U75 ( .A(n69), .Y(n70) );
  AND2X2 U76 ( .A(\in<14> ), .B(n138), .Y(n71) );
  INVX1 U77 ( .A(n71), .Y(n72) );
  AND2X2 U78 ( .A(\in<13> ), .B(n120), .Y(n73) );
  INVX1 U79 ( .A(n73), .Y(n74) );
  AND2X2 U80 ( .A(\in<14> ), .B(n140), .Y(n75) );
  INVX1 U81 ( .A(n75), .Y(n76) );
  AND2X2 U82 ( .A(n142), .B(n7), .Y(n77) );
  INVX1 U83 ( .A(n77), .Y(n78) );
  AND2X2 U84 ( .A(\in<0> ), .B(n140), .Y(n79) );
  INVX1 U85 ( .A(n79), .Y(n80) );
  AND2X2 U86 ( .A(n136), .B(\in<3> ), .Y(n81) );
  INVX1 U87 ( .A(n81), .Y(n82) );
  AND2X2 U88 ( .A(\in<5> ), .B(n139), .Y(n83) );
  INVX1 U89 ( .A(n83), .Y(n84) );
  AND2X2 U90 ( .A(\in<4> ), .B(n3), .Y(n85) );
  INVX1 U91 ( .A(n85), .Y(n86) );
  AND2X2 U92 ( .A(\in<7> ), .B(n10), .Y(n87) );
  INVX1 U93 ( .A(n87), .Y(n88) );
  AND2X2 U94 ( .A(\in<9> ), .B(n10), .Y(n89) );
  INVX1 U95 ( .A(n89), .Y(n90) );
  AND2X2 U96 ( .A(\in<10> ), .B(n9), .Y(n91) );
  INVX1 U97 ( .A(n91), .Y(n92) );
  AND2X2 U98 ( .A(\in<11> ), .B(n10), .Y(n93) );
  INVX1 U99 ( .A(n93), .Y(n94) );
  AND2X2 U100 ( .A(n132), .B(\in<13> ), .Y(n95) );
  INVX1 U101 ( .A(n95), .Y(n96) );
  AND2X2 U102 ( .A(sh), .B(n6), .Y(n97) );
  AND2X2 U103 ( .A(sh), .B(n121), .Y(n98) );
  INVX1 U104 ( .A(n98), .Y(n99) );
  INVX1 U105 ( .A(n98), .Y(n100) );
  AND2X2 U106 ( .A(\in<2> ), .B(n130), .Y(n101) );
  INVX1 U107 ( .A(n101), .Y(n102) );
  INVX1 U108 ( .A(\op<1> ), .Y(n104) );
  INVX1 U109 ( .A(n141), .Y(n103) );
  MUX2X1 U110 ( .B(n141), .A(n58), .S(n104), .Y(n142) );
  AND2X2 U111 ( .A(\in<4> ), .B(n131), .Y(n105) );
  INVX1 U112 ( .A(n105), .Y(n106) );
  INVX1 U113 ( .A(n17), .Y(n107) );
  AND2X2 U114 ( .A(n131), .B(\in<0> ), .Y(n108) );
  INVX1 U115 ( .A(n108), .Y(n109) );
  AND2X2 U116 ( .A(\in<1> ), .B(n137), .Y(n110) );
  INVX1 U117 ( .A(n110), .Y(n111) );
  AND2X2 U118 ( .A(n137), .B(\in<14> ), .Y(n112) );
  INVX1 U119 ( .A(n112), .Y(n113) );
  AND2X2 U120 ( .A(n103), .B(n131), .Y(n114) );
  INVX1 U121 ( .A(n114), .Y(n115) );
  AND2X2 U122 ( .A(\in<9> ), .B(n135), .Y(n116) );
  INVX1 U123 ( .A(n116), .Y(n117) );
  AND2X2 U124 ( .A(\in<11> ), .B(n130), .Y(n118) );
  INVX1 U125 ( .A(n118), .Y(n119) );
  NAND3X1 U126 ( .A(n21), .B(n64), .C(n86), .Y(\out<5> ) );
  NAND3X1 U127 ( .A(n111), .B(n80), .C(n60), .Y(\out<1> ) );
  INVX1 U128 ( .A(n100), .Y(n120) );
  INVX1 U129 ( .A(n127), .Y(n121) );
  INVX1 U130 ( .A(\op<0> ), .Y(n122) );
  INVX1 U131 ( .A(\op<2> ), .Y(n126) );
  INVX1 U132 ( .A(n97), .Y(n123) );
  INVX1 U133 ( .A(n97), .Y(n124) );
  INVX1 U134 ( .A(n97), .Y(n125) );
  INVX1 U135 ( .A(sh), .Y(n133) );
  INVX1 U136 ( .A(sh), .Y(n130) );
  INVX1 U137 ( .A(sh), .Y(n135) );
  INVX1 U138 ( .A(sh), .Y(n137) );
  OR2X2 U139 ( .A(n2), .B(n5), .Y(n127) );
  INVX1 U140 ( .A(n125), .Y(n134) );
  INVX1 U141 ( .A(n125), .Y(n138) );
  INVX1 U142 ( .A(n124), .Y(n139) );
  INVX1 U143 ( .A(n123), .Y(n136) );
  INVX1 U144 ( .A(n123), .Y(n132) );
  AOI21X1 U145 ( .A(\in<1> ), .B(n12), .C(n16), .Y(n129) );
  NAND3X1 U146 ( .A(n102), .B(n62), .C(n82), .Y(\out<2> ) );
  NAND3X1 U147 ( .A(n38), .B(n107), .C(n19), .Y(\out<3> ) );
  NAND3X1 U148 ( .A(n40), .B(n106), .C(n84), .Y(\out<4> ) );
  NAND3X1 U149 ( .A(n42), .B(n23), .C(n88), .Y(\out<6> ) );
  NAND3X1 U150 ( .A(n44), .B(n25), .C(n66), .Y(\out<7> ) );
  NAND3X1 U151 ( .A(n46), .B(n27), .C(n90), .Y(\out<8> ) );
  NAND3X1 U152 ( .A(n48), .B(n117), .C(n92), .Y(\out<9> ) );
  NAND3X1 U153 ( .A(n29), .B(n68), .C(n94), .Y(\out<10> ) );
  NAND3X1 U154 ( .A(n50), .B(n119), .C(n70), .Y(\out<11> ) );
  NAND3X1 U155 ( .A(n52), .B(n31), .C(n96), .Y(\out<12> ) );
  NAND3X1 U156 ( .A(n54), .B(n33), .C(n72), .Y(\out<13> ) );
  NAND3X1 U157 ( .A(n113), .B(n74), .C(n56), .Y(\out<14> ) );
  NAND3X1 U158 ( .A(n115), .B(n76), .C(n78), .Y(\out<15> ) );
endmodule


module shifter_2 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), .op({\op<2> , \op<1> , \op<0> }), 
        sh, .out({\out<15> , \out<14> , \out<13> , \out<12> , \out<11> , 
        \out<10> , \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , 
        \out<3> , \out<2> , \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , \op<2> , \op<1> , \op<0> , sh;
  output \out<15> , \out<14> , \out<13> , \out<12> , \out<11> , \out<10> ,
         \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> ,
         \out<2> , \out<1> , \out<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148;

  INVX1 U2 ( .A(n114), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n121), .Y(n3) );
  INVX1 U5 ( .A(n3), .Y(n4) );
  INVX1 U6 ( .A(n116), .Y(n5) );
  INVX1 U7 ( .A(n5), .Y(n6) );
  BUFX2 U8 ( .A(n121), .Y(n7) );
  INVX1 U9 ( .A(n117), .Y(n8) );
  INVX1 U10 ( .A(n8), .Y(n9) );
  AND2X2 U11 ( .A(n115), .B(n21), .Y(n62) );
  INVX1 U12 ( .A(n119), .Y(n10) );
  INVX1 U13 ( .A(n10), .Y(n11) );
  INVX1 U14 ( .A(n106), .Y(n12) );
  INVX1 U15 ( .A(n12), .Y(n13) );
  INVX1 U16 ( .A(n106), .Y(n14) );
  BUFX2 U17 ( .A(\in<0> ), .Y(n15) );
  INVX1 U18 ( .A(n17), .Y(\out<2> ) );
  AND2X2 U19 ( .A(n112), .B(n136), .Y(n40) );
  AND2X2 U20 ( .A(n35), .B(n36), .Y(n16) );
  AND2X2 U21 ( .A(n25), .B(n16), .Y(n17) );
  AND2X2 U22 ( .A(n31), .B(n34), .Y(n19) );
  INVX1 U23 ( .A(n19), .Y(\out<10> ) );
  AND2X2 U24 ( .A(n144), .B(n123), .Y(n21) );
  OR2X2 U25 ( .A(n109), .B(\op<1> ), .Y(n22) );
  INVX1 U26 ( .A(n22), .Y(n23) );
  AND2X2 U27 ( .A(n145), .B(n125), .Y(n24) );
  INVX1 U28 ( .A(n24), .Y(n25) );
  AND2X2 U29 ( .A(n113), .B(n136), .Y(n26) );
  INVX1 U30 ( .A(n26), .Y(n27) );
  AND2X2 U31 ( .A(n118), .B(n145), .Y(n28) );
  INVX1 U32 ( .A(n28), .Y(n29) );
  AND2X2 U33 ( .A(n120), .B(n145), .Y(n30) );
  INVX1 U34 ( .A(n30), .Y(n31) );
  AND2X2 U35 ( .A(n117), .B(n145), .Y(n32) );
  BUFX2 U36 ( .A(n142), .Y(n33) );
  BUFX2 U37 ( .A(n141), .Y(n34) );
  OR2X2 U38 ( .A(n128), .B(n127), .Y(n35) );
  OR2X2 U39 ( .A(n126), .B(n14), .Y(n36) );
  BUFX2 U40 ( .A(n140), .Y(n37) );
  AND2X2 U41 ( .A(\in<0> ), .B(n145), .Y(n38) );
  INVX1 U42 ( .A(n38), .Y(n39) );
  INVX1 U43 ( .A(n40), .Y(n41) );
  AND2X2 U44 ( .A(n13), .B(n145), .Y(n42) );
  INVX1 U45 ( .A(n42), .Y(n43) );
  AND2X2 U46 ( .A(n147), .B(n110), .Y(n44) );
  INVX1 U47 ( .A(n44), .Y(n45) );
  AND2X2 U48 ( .A(n106), .B(n147), .Y(n46) );
  INVX1 U49 ( .A(n46), .Y(n47) );
  AND2X2 U50 ( .A(n7), .B(n145), .Y(n48) );
  INVX1 U51 ( .A(n48), .Y(n49) );
  AND2X2 U52 ( .A(n147), .B(n118), .Y(n50) );
  INVX1 U53 ( .A(n50), .Y(n51) );
  AND2X2 U54 ( .A(n147), .B(n121), .Y(n52) );
  INVX1 U55 ( .A(n52), .Y(n53) );
  AND2X2 U56 ( .A(n9), .B(n136), .Y(n54) );
  INVX1 U57 ( .A(n54), .Y(n55) );
  AND2X2 U58 ( .A(n145), .B(n107), .Y(n56) );
  INVX1 U59 ( .A(n56), .Y(n57) );
  AND2X2 U60 ( .A(n147), .B(n117), .Y(n58) );
  INVX1 U61 ( .A(n58), .Y(n59) );
  AND2X2 U62 ( .A(n137), .B(sh), .Y(n60) );
  INVX1 U63 ( .A(n60), .Y(n61) );
  INVX1 U64 ( .A(n62), .Y(n63) );
  AND2X2 U65 ( .A(n111), .B(n136), .Y(n64) );
  INVX1 U66 ( .A(n64), .Y(n65) );
  AND2X2 U67 ( .A(n110), .B(n132), .Y(n66) );
  INVX1 U68 ( .A(n66), .Y(n67) );
  AND2X2 U69 ( .A(n115), .B(n147), .Y(n68) );
  INVX1 U70 ( .A(n68), .Y(n69) );
  AND2X2 U71 ( .A(n147), .B(n111), .Y(n70) );
  INVX1 U72 ( .A(n70), .Y(n71) );
  AND2X2 U73 ( .A(n4), .B(n132), .Y(n72) );
  INVX1 U74 ( .A(n72), .Y(n73) );
  AND2X2 U75 ( .A(n11), .B(n132), .Y(n74) );
  INVX1 U76 ( .A(n74), .Y(n75) );
  AND2X2 U77 ( .A(n145), .B(n113), .Y(n76) );
  INVX1 U78 ( .A(n76), .Y(n77) );
  AND2X2 U79 ( .A(n136), .B(n116), .Y(n78) );
  INVX1 U80 ( .A(n78), .Y(n79) );
  AND2X2 U81 ( .A(n6), .B(n145), .Y(n80) );
  INVX1 U82 ( .A(n80), .Y(n81) );
  AND2X2 U83 ( .A(n147), .B(n120), .Y(n82) );
  INVX1 U84 ( .A(n82), .Y(n83) );
  AND2X2 U85 ( .A(n116), .B(n147), .Y(n84) );
  INVX1 U86 ( .A(n84), .Y(n85) );
  AND2X2 U87 ( .A(n145), .B(n112), .Y(n86) );
  INVX1 U88 ( .A(n86), .Y(n87) );
  AND2X2 U89 ( .A(n23), .B(n108), .Y(n88) );
  INVX1 U90 ( .A(n88), .Y(n89) );
  AND2X2 U91 ( .A(n145), .B(n110), .Y(n90) );
  INVX1 U92 ( .A(n90), .Y(n91) );
  AND2X2 U93 ( .A(n118), .B(n136), .Y(n92) );
  INVX1 U94 ( .A(n92), .Y(n93) );
  AND2X2 U95 ( .A(n112), .B(n147), .Y(n94) );
  INVX1 U96 ( .A(n94), .Y(n95) );
  AND2X2 U97 ( .A(n136), .B(n120), .Y(n96) );
  INVX1 U98 ( .A(n96), .Y(n97) );
  AND2X2 U99 ( .A(n145), .B(n119), .Y(n98) );
  INVX1 U100 ( .A(n98), .Y(n99) );
  AND2X2 U101 ( .A(n11), .B(n147), .Y(n100) );
  INVX1 U102 ( .A(n100), .Y(n101) );
  AND2X2 U103 ( .A(n136), .B(n108), .Y(n102) );
  INVX1 U104 ( .A(n102), .Y(n103) );
  AND2X2 U105 ( .A(n114), .B(n132), .Y(n104) );
  INVX1 U106 ( .A(n104), .Y(n105) );
  BUFX2 U107 ( .A(\in<4> ), .Y(n106) );
  BUFX2 U108 ( .A(\in<12> ), .Y(n107) );
  BUFX2 U109 ( .A(\in<14> ), .Y(n108) );
  BUFX2 U110 ( .A(n138), .Y(n109) );
  BUFX2 U111 ( .A(\in<3> ), .Y(n110) );
  BUFX2 U112 ( .A(\in<2> ), .Y(n111) );
  BUFX2 U113 ( .A(\in<5> ), .Y(n112) );
  BUFX2 U114 ( .A(\in<8> ), .Y(n113) );
  BUFX2 U115 ( .A(\in<15> ), .Y(n114) );
  BUFX2 U116 ( .A(\in<1> ), .Y(n115) );
  BUFX2 U117 ( .A(\in<11> ), .Y(n116) );
  BUFX2 U118 ( .A(\in<13> ), .Y(n117) );
  BUFX2 U119 ( .A(\in<6> ), .Y(n118) );
  BUFX2 U120 ( .A(\in<9> ), .Y(n119) );
  BUFX2 U121 ( .A(\in<10> ), .Y(n120) );
  BUFX2 U122 ( .A(\in<7> ), .Y(n121) );
  INVX1 U123 ( .A(n32), .Y(n122) );
  AND2X2 U124 ( .A(\op<0> ), .B(sh), .Y(n123) );
  MUX2X1 U125 ( .B(n61), .A(n130), .S(n133), .Y(n131) );
  INVX1 U126 ( .A(n111), .Y(n124) );
  INVX1 U127 ( .A(n124), .Y(n125) );
  INVX2 U128 ( .A(sh), .Y(n145) );
  INVX1 U129 ( .A(n132), .Y(n126) );
  INVX1 U130 ( .A(n147), .Y(n127) );
  INVX1 U131 ( .A(\in<0> ), .Y(n128) );
  BUFX4 U132 ( .A(n131), .Y(n132) );
  NAND3X1 U133 ( .A(n122), .B(n85), .C(n105), .Y(\out<13> ) );
  AND2X2 U134 ( .A(n145), .B(n115), .Y(n129) );
  INVX1 U135 ( .A(n129), .Y(n139) );
  NAND3X1 U136 ( .A(n49), .B(n75), .C(n95), .Y(\out<7> ) );
  INVX1 U137 ( .A(n123), .Y(n130) );
  MUX2X1 U138 ( .B(n2), .A(n15), .S(n144), .Y(n143) );
  INVX1 U139 ( .A(\op<1> ), .Y(n144) );
  INVX1 U140 ( .A(\op<2> ), .Y(n133) );
  INVX1 U141 ( .A(n107), .Y(n134) );
  INVX1 U142 ( .A(n134), .Y(n135) );
  INVX1 U143 ( .A(\op<0> ), .Y(n137) );
  BUFX4 U144 ( .A(n131), .Y(n136) );
  INVX4 U145 ( .A(n109), .Y(n147) );
  NAND3X1 U146 ( .A(n137), .B(sh), .C(n133), .Y(n138) );
  NAND3X1 U147 ( .A(n39), .B(n65), .C(n89), .Y(\out<0> ) );
  NAND3X1 U148 ( .A(n114), .B(n147), .C(n144), .Y(n140) );
  NAND3X1 U149 ( .A(n37), .B(n67), .C(n139), .Y(\out<1> ) );
  NAND3X1 U150 ( .A(n41), .B(n69), .C(n91), .Y(\out<3> ) );
  NAND3X1 U151 ( .A(n71), .B(n93), .C(n43), .Y(\out<4> ) );
  NAND3X1 U152 ( .A(n45), .B(n73), .C(n87), .Y(\out<5> ) );
  NAND3X1 U153 ( .A(n47), .B(n27), .C(n29), .Y(\out<6> ) );
  NAND3X1 U154 ( .A(n51), .B(n77), .C(n97), .Y(\out<8> ) );
  NAND3X1 U155 ( .A(n99), .B(n53), .C(n79), .Y(\out<9> ) );
  AOI22X1 U156 ( .A(n132), .B(n107), .C(n113), .D(n147), .Y(n141) );
  NAND3X1 U157 ( .A(n55), .B(n81), .C(n101), .Y(\out<11> ) );
  NAND3X1 U158 ( .A(n57), .B(n83), .C(n103), .Y(\out<12> ) );
  AOI22X1 U159 ( .A(n145), .B(n108), .C(n135), .D(n147), .Y(n142) );
  OAI21X1 U160 ( .A(n130), .B(n143), .C(n33), .Y(\out<14> ) );
  AND2X2 U161 ( .A(\op<1> ), .B(\op<0> ), .Y(n146) );
  OAI21X1 U162 ( .A(n146), .B(n145), .C(n2), .Y(n148) );
  NAND3X1 U163 ( .A(n59), .B(n63), .C(n148), .Y(\out<15> ) );
endmodule


module shifter_4 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), .op({\op<2> , \op<1> , \op<0> }), 
        sh, .out({\out<15> , \out<14> , \out<13> , \out<12> , \out<11> , 
        \out<10> , \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , 
        \out<3> , \out<2> , \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , \op<2> , \op<1> , \op<0> , sh;
  output \out<15> , \out<14> , \out<13> , \out<12> , \out<11> , \out<10> ,
         \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> ,
         \out<2> , \out<1> , \out<0> ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n10, n11, n13, n15, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144;

  INVX1 U2 ( .A(n108), .Y(n1) );
  INVX1 U3 ( .A(n1), .Y(n2) );
  INVX1 U4 ( .A(n118), .Y(n3) );
  INVX2 U5 ( .A(n133), .Y(n136) );
  AND2X1 U6 ( .A(n101), .B(n142), .Y(n32) );
  AND2X1 U7 ( .A(n100), .B(n142), .Y(n68) );
  INVX1 U8 ( .A(n96), .Y(n4) );
  INVX1 U9 ( .A(n129), .Y(n5) );
  INVX1 U10 ( .A(n7), .Y(n6) );
  INVX1 U11 ( .A(\in<2> ), .Y(n7) );
  INVX1 U12 ( .A(n7), .Y(n8) );
  AND2X2 U13 ( .A(n100), .B(n112), .Y(n124) );
  OR2X2 U14 ( .A(n10), .B(n21), .Y(\out<5> ) );
  INVX1 U15 ( .A(n139), .Y(n10) );
  AND2X2 U16 ( .A(n104), .B(n142), .Y(n21) );
  AND2X2 U17 ( .A(n96), .B(n142), .Y(n39) );
  AND2X2 U18 ( .A(n40), .B(n36), .Y(n11) );
  INVX1 U19 ( .A(n11), .Y(\out<1> ) );
  AND2X2 U20 ( .A(n42), .B(n37), .Y(n13) );
  INVX1 U21 ( .A(n13), .Y(\out<3> ) );
  AND2X2 U22 ( .A(n44), .B(n38), .Y(n15) );
  INVX1 U23 ( .A(n15), .Y(\out<15> ) );
  AND2X2 U24 ( .A(\op<1> ), .B(n109), .Y(n17) );
  AND2X2 U25 ( .A(sh), .B(n134), .Y(n18) );
  AND2X2 U26 ( .A(n100), .B(n18), .Y(n19) );
  INVX1 U27 ( .A(n19), .Y(n20) );
  AND2X2 U28 ( .A(n112), .B(n6), .Y(n22) );
  INVX1 U29 ( .A(n22), .Y(n23) );
  AND2X2 U30 ( .A(n18), .B(\in<10> ), .Y(n24) );
  INVX1 U31 ( .A(n24), .Y(n25) );
  AND2X2 U32 ( .A(n101), .B(n18), .Y(n26) );
  INVX1 U33 ( .A(n26), .Y(n27) );
  AND2X2 U34 ( .A(n3), .B(n142), .Y(n28) );
  INVX1 U35 ( .A(n28), .Y(n29) );
  AND2X2 U36 ( .A(n142), .B(\in<10> ), .Y(n30) );
  INVX1 U37 ( .A(n30), .Y(n31) );
  INVX1 U38 ( .A(n32), .Y(n33) );
  AND2X2 U39 ( .A(n122), .B(n110), .Y(n34) );
  INVX1 U40 ( .A(n34), .Y(n35) );
  BUFX2 U41 ( .A(n135), .Y(n36) );
  BUFX2 U42 ( .A(n137), .Y(n37) );
  BUFX2 U43 ( .A(n144), .Y(n38) );
  INVX1 U44 ( .A(n39), .Y(n40) );
  AND2X1 U45 ( .A(n128), .B(n142), .Y(n41) );
  INVX1 U46 ( .A(n41), .Y(n42) );
  AND2X1 U47 ( .A(n101), .B(n112), .Y(n43) );
  INVX1 U48 ( .A(n43), .Y(n44) );
  AND2X2 U49 ( .A(n136), .B(n94), .Y(n45) );
  INVX1 U50 ( .A(n45), .Y(n46) );
  AND2X1 U51 ( .A(\in<2> ), .B(n142), .Y(n47) );
  INVX1 U52 ( .A(n47), .Y(n48) );
  AND2X2 U53 ( .A(n122), .B(n112), .Y(n49) );
  INVX1 U54 ( .A(n49), .Y(n50) );
  AND2X2 U55 ( .A(n128), .B(n112), .Y(n51) );
  INVX1 U56 ( .A(n51), .Y(n52) );
  AND2X2 U57 ( .A(n112), .B(n98), .Y(n53) );
  INVX1 U58 ( .A(n53), .Y(n54) );
  AND2X2 U59 ( .A(n112), .B(n104), .Y(n55) );
  INVX1 U60 ( .A(n55), .Y(n56) );
  AND2X2 U61 ( .A(n18), .B(\in<14> ), .Y(n57) );
  INVX1 U62 ( .A(n57), .Y(n58) );
  AND2X2 U63 ( .A(n102), .B(n112), .Y(n59) );
  INVX1 U64 ( .A(n59), .Y(n60) );
  AND2X2 U65 ( .A(n142), .B(n126), .Y(n61) );
  INVX1 U66 ( .A(n61), .Y(n62) );
  BUFX2 U67 ( .A(n141), .Y(n63) );
  AND2X1 U68 ( .A(n95), .B(n142), .Y(n64) );
  INVX1 U69 ( .A(n64), .Y(n65) );
  AND2X2 U70 ( .A(\in<14> ), .B(n136), .Y(n66) );
  INVX1 U71 ( .A(n66), .Y(n67) );
  INVX1 U72 ( .A(n68), .Y(n69) );
  AND2X2 U73 ( .A(n99), .B(n112), .Y(n70) );
  INVX1 U74 ( .A(n70), .Y(n71) );
  AND2X2 U75 ( .A(n130), .B(n18), .Y(n72) );
  INVX1 U76 ( .A(n72), .Y(n73) );
  BUFX2 U77 ( .A(n143), .Y(n74) );
  OR2X2 U78 ( .A(n124), .B(n123), .Y(n75) );
  INVX1 U79 ( .A(n75), .Y(n76) );
  AND2X2 U80 ( .A(n18), .B(n98), .Y(n77) );
  INVX1 U81 ( .A(n77), .Y(n78) );
  AND2X2 U82 ( .A(n18), .B(n99), .Y(n79) );
  INVX1 U83 ( .A(n79), .Y(n80) );
  AND2X2 U84 ( .A(n142), .B(n98), .Y(n81) );
  INVX1 U85 ( .A(n81), .Y(n82) );
  AND2X1 U86 ( .A(n120), .B(n142), .Y(n83) );
  INVX1 U87 ( .A(n83), .Y(n84) );
  AND2X1 U88 ( .A(n102), .B(n142), .Y(n85) );
  INVX1 U89 ( .A(n85), .Y(n86) );
  AND2X2 U90 ( .A(n18), .B(n94), .Y(n87) );
  INVX1 U91 ( .A(n87), .Y(n88) );
  AND2X2 U92 ( .A(n108), .B(n18), .Y(n89) );
  INVX1 U93 ( .A(n89), .Y(n90) );
  AND2X2 U94 ( .A(n96), .B(n110), .Y(n91) );
  INVX1 U95 ( .A(n91), .Y(n92) );
  BUFX2 U96 ( .A(\in<15> ), .Y(n93) );
  BUFX2 U97 ( .A(\in<12> ), .Y(n94) );
  BUFX2 U98 ( .A(\in<0> ), .Y(n95) );
  BUFX2 U99 ( .A(\in<1> ), .Y(n96) );
  BUFX2 U100 ( .A(\in<3> ), .Y(n97) );
  BUFX2 U101 ( .A(\in<4> ), .Y(n98) );
  BUFX2 U102 ( .A(\in<6> ), .Y(n99) );
  BUFX2 U103 ( .A(\in<8> ), .Y(n100) );
  BUFX2 U104 ( .A(\in<11> ), .Y(n101) );
  BUFX2 U105 ( .A(\in<7> ), .Y(n102) );
  BUFX2 U106 ( .A(\in<9> ), .Y(n103) );
  BUFX2 U107 ( .A(\in<5> ), .Y(n104) );
  AND2X2 U108 ( .A(n17), .B(n93), .Y(n105) );
  INVX1 U109 ( .A(n105), .Y(n106) );
  INVX1 U110 ( .A(n105), .Y(n107) );
  BUFX2 U111 ( .A(\in<13> ), .Y(n108) );
  AND2X2 U112 ( .A(sh), .B(\op<0> ), .Y(n109) );
  AND2X2 U113 ( .A(n140), .B(n109), .Y(n110) );
  BUFX2 U114 ( .A(n138), .Y(n111) );
  INVX1 U115 ( .A(n111), .Y(n112) );
  BUFX2 U116 ( .A(n107), .Y(n113) );
  INVX1 U117 ( .A(\op<1> ), .Y(n140) );
  AND2X2 U118 ( .A(\op<1> ), .B(\op<0> ), .Y(n114) );
  INVX1 U119 ( .A(n114), .Y(n115) );
  AND2X2 U120 ( .A(n115), .B(sh), .Y(n116) );
  INVX1 U121 ( .A(n116), .Y(n117) );
  INVX1 U122 ( .A(n103), .Y(n118) );
  INVX1 U123 ( .A(n118), .Y(n119) );
  BUFX2 U124 ( .A(n99), .Y(n120) );
  INVX1 U125 ( .A(n95), .Y(n121) );
  INVX1 U126 ( .A(n121), .Y(n122) );
  AND2X2 U127 ( .A(n142), .B(n94), .Y(n123) );
  INVX1 U128 ( .A(n4), .Y(n125) );
  BUFX2 U129 ( .A(\in<14> ), .Y(n126) );
  INVX1 U130 ( .A(sh), .Y(n142) );
  INVX1 U131 ( .A(\op<2> ), .Y(n131) );
  INVX1 U132 ( .A(\op<0> ), .Y(n132) );
  INVX1 U133 ( .A(n97), .Y(n127) );
  INVX1 U134 ( .A(n127), .Y(n128) );
  INVX1 U135 ( .A(n93), .Y(n129) );
  INVX1 U136 ( .A(n129), .Y(n130) );
  NAND3X1 U137 ( .A(sh), .B(n132), .C(n131), .Y(n138) );
  OR2X2 U138 ( .A(n111), .B(\op<1> ), .Y(n133) );
  XOR2X1 U139 ( .A(\op<2> ), .B(\op<0> ), .Y(n134) );
  NAND3X1 U140 ( .A(n65), .B(n46), .C(n78), .Y(\out<0> ) );
  AOI22X1 U141 ( .A(n18), .B(n104), .C(n2), .D(n136), .Y(n135) );
  NAND3X1 U142 ( .A(n67), .B(n48), .C(n80), .Y(\out<2> ) );
  AOI22X1 U143 ( .A(n18), .B(n102), .C(n5), .D(n136), .Y(n137) );
  NAND3X1 U144 ( .A(n50), .B(n20), .C(n82), .Y(\out<4> ) );
  AOI22X1 U145 ( .A(n119), .B(n18), .C(n125), .D(n112), .Y(n139) );
  NAND3X1 U146 ( .A(n23), .B(n25), .C(n84), .Y(\out<6> ) );
  NAND3X1 U147 ( .A(n52), .B(n27), .C(n86), .Y(\out<7> ) );
  NAND3X1 U148 ( .A(n88), .B(n69), .C(n54), .Y(\out<8> ) );
  NAND3X1 U149 ( .A(n56), .B(n29), .C(n90), .Y(\out<9> ) );
  NAND3X1 U150 ( .A(n58), .B(n71), .C(n31), .Y(\out<10> ) );
  NAND3X1 U151 ( .A(n60), .B(n73), .C(n33), .Y(\out<11> ) );
  NAND3X1 U152 ( .A(n35), .B(n107), .C(n76), .Y(\out<12> ) );
  AOI22X1 U153 ( .A(n112), .B(n103), .C(n142), .D(n108), .Y(n141) );
  NAND3X1 U154 ( .A(n106), .B(n92), .C(n63), .Y(\out<13> ) );
  AOI22X1 U155 ( .A(n112), .B(\in<10> ), .C(n110), .D(n8), .Y(n143) );
  NAND3X1 U156 ( .A(n62), .B(n113), .C(n74), .Y(\out<14> ) );
  AOI22X1 U157 ( .A(n110), .B(n97), .C(n93), .D(n117), .Y(n144) );
endmodule


module shifter_8 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), .op({\op<2> , \op<1> , \op<0> }), 
        sh, .out({\out<15> , \out<14> , \out<13> , \out<12> , \out<11> , 
        \out<10> , \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , 
        \out<3> , \out<2> , \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , \op<2> , \op<1> , \op<0> , sh;
  output \out<15> , \out<14> , \out<13> , \out<12> , \out<11> , \out<10> ,
         \out<9> , \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> ,
         \out<2> , \out<1> , \out<0> ;
  wire   n1, n2, n3, n4, n6, n8, n10, n12, n14, n16, n18, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  AND2X1 U2 ( .A(n33), .B(n35), .Y(n101) );
  AND2X1 U3 ( .A(n91), .B(n120), .Y(n64) );
  AND2X1 U4 ( .A(n93), .B(n120), .Y(n68) );
  AND2X1 U5 ( .A(n94), .B(n120), .Y(n21) );
  BUFX2 U6 ( .A(n98), .Y(n1) );
  INVX1 U7 ( .A(n88), .Y(n2) );
  INVX1 U8 ( .A(n2), .Y(n3) );
  AND2X2 U9 ( .A(\in<15> ), .B(n20), .Y(n86) );
  AND2X1 U10 ( .A(\in<1> ), .B(n120), .Y(n52) );
  INVX1 U11 ( .A(n86), .Y(n113) );
  AND2X2 U12 ( .A(n37), .B(n51), .Y(n4) );
  INVX1 U13 ( .A(n4), .Y(\out<0> ) );
  AND2X2 U14 ( .A(n53), .B(n39), .Y(n6) );
  INVX1 U15 ( .A(n6), .Y(\out<1> ) );
  AND2X2 U16 ( .A(n41), .B(n55), .Y(n8) );
  INVX1 U17 ( .A(n8), .Y(\out<2> ) );
  AND2X2 U18 ( .A(n57), .B(n43), .Y(n10) );
  INVX1 U19 ( .A(n10), .Y(\out<3> ) );
  AND2X2 U20 ( .A(n22), .B(n45), .Y(n12) );
  INVX1 U21 ( .A(n12), .Y(\out<4> ) );
  AND2X2 U22 ( .A(n59), .B(n47), .Y(n14) );
  INVX1 U23 ( .A(n14), .Y(\out<5> ) );
  AND2X2 U24 ( .A(n61), .B(n49), .Y(n16) );
  INVX1 U25 ( .A(n16), .Y(\out<6> ) );
  AND2X2 U26 ( .A(n63), .B(n31), .Y(n18) );
  INVX1 U27 ( .A(n18), .Y(\out<15> ) );
  AND2X2 U28 ( .A(\op<1> ), .B(n118), .Y(n20) );
  INVX1 U29 ( .A(n21), .Y(n22) );
  AND2X2 U30 ( .A(sh), .B(n100), .Y(n23) );
  AND2X2 U31 ( .A(n119), .B(n23), .Y(n24) );
  AND2X2 U32 ( .A(n3), .B(n120), .Y(n25) );
  AND2X2 U33 ( .A(n92), .B(n120), .Y(n26) );
  INVX1 U34 ( .A(n26), .Y(n27) );
  AND2X2 U35 ( .A(\in<3> ), .B(n24), .Y(n28) );
  INVX1 U36 ( .A(n28), .Y(n29) );
  AND2X2 U37 ( .A(n104), .B(n107), .Y(n30) );
  INVX1 U38 ( .A(n30), .Y(n31) );
  AND2X1 U39 ( .A(n96), .B(n120), .Y(n32) );
  INVX1 U40 ( .A(n32), .Y(n33) );
  AND2X2 U41 ( .A(n117), .B(n107), .Y(n34) );
  INVX1 U42 ( .A(n34), .Y(n35) );
  AND2X2 U43 ( .A(n117), .B(n88), .Y(n36) );
  INVX1 U44 ( .A(n36), .Y(n37) );
  AND2X2 U45 ( .A(n117), .B(n91), .Y(n38) );
  INVX1 U46 ( .A(n38), .Y(n39) );
  AND2X2 U47 ( .A(n117), .B(n92), .Y(n40) );
  INVX1 U48 ( .A(n40), .Y(n41) );
  AND2X2 U49 ( .A(n97), .B(n117), .Y(n42) );
  INVX1 U50 ( .A(n42), .Y(n43) );
  AND2X2 U51 ( .A(n117), .B(n90), .Y(n44) );
  INVX1 U52 ( .A(n44), .Y(n45) );
  AND2X2 U53 ( .A(n1), .B(n117), .Y(n46) );
  INVX1 U54 ( .A(n46), .Y(n47) );
  AND2X2 U55 ( .A(n93), .B(n117), .Y(n48) );
  INVX1 U56 ( .A(n48), .Y(n49) );
  AND2X1 U57 ( .A(n105), .B(n120), .Y(n50) );
  INVX1 U58 ( .A(n50), .Y(n51) );
  INVX1 U59 ( .A(n52), .Y(n53) );
  AND2X1 U60 ( .A(n89), .B(n120), .Y(n54) );
  INVX1 U61 ( .A(n54), .Y(n55) );
  AND2X2 U62 ( .A(n120), .B(\in<3> ), .Y(n56) );
  INVX1 U63 ( .A(n56), .Y(n57) );
  AND2X2 U64 ( .A(n120), .B(\in<5> ), .Y(n58) );
  INVX1 U65 ( .A(n58), .Y(n59) );
  AND2X1 U66 ( .A(n95), .B(n120), .Y(n60) );
  INVX1 U67 ( .A(n60), .Y(n61) );
  AND2X2 U68 ( .A(n96), .B(n24), .Y(n62) );
  INVX1 U69 ( .A(n62), .Y(n63) );
  INVX1 U70 ( .A(n64), .Y(n65) );
  AND2X1 U71 ( .A(n97), .B(n120), .Y(n66) );
  INVX1 U72 ( .A(n66), .Y(n67) );
  INVX1 U73 ( .A(n68), .Y(n69) );
  AND2X2 U74 ( .A(n111), .B(n24), .Y(n70) );
  INVX1 U75 ( .A(n70), .Y(n71) );
  AND2X2 U76 ( .A(\in<1> ), .B(n24), .Y(n72) );
  INVX1 U77 ( .A(n72), .Y(n73) );
  AND2X2 U78 ( .A(n24), .B(n109), .Y(n74) );
  INVX1 U79 ( .A(n74), .Y(n75) );
  AND2X2 U80 ( .A(n94), .B(n24), .Y(n76) );
  INVX1 U81 ( .A(n76), .Y(n77) );
  AND2X1 U82 ( .A(n98), .B(n120), .Y(n78) );
  INVX1 U83 ( .A(n78), .Y(n79) );
  AND2X2 U84 ( .A(n95), .B(n24), .Y(n80) );
  INVX1 U85 ( .A(n80), .Y(n81) );
  AND2X2 U86 ( .A(n90), .B(n120), .Y(n82) );
  INVX1 U87 ( .A(n82), .Y(n83) );
  AND2X2 U88 ( .A(\in<5> ), .B(n24), .Y(n84) );
  INVX1 U89 ( .A(n84), .Y(n85) );
  INVX1 U90 ( .A(n86), .Y(n87) );
  BUFX2 U91 ( .A(\in<8> ), .Y(n88) );
  BUFX2 U92 ( .A(\in<2> ), .Y(n89) );
  BUFX2 U93 ( .A(\in<12> ), .Y(n90) );
  BUFX2 U94 ( .A(\in<9> ), .Y(n91) );
  BUFX2 U95 ( .A(\in<10> ), .Y(n92) );
  BUFX2 U96 ( .A(\in<14> ), .Y(n93) );
  BUFX2 U97 ( .A(\in<4> ), .Y(n94) );
  BUFX2 U98 ( .A(\in<6> ), .Y(n95) );
  BUFX2 U99 ( .A(\in<7> ), .Y(n96) );
  BUFX2 U100 ( .A(\in<11> ), .Y(n97) );
  BUFX2 U101 ( .A(\in<13> ), .Y(n98) );
  INVX1 U102 ( .A(\op<1> ), .Y(n115) );
  INVX1 U103 ( .A(sh), .Y(n120) );
  AND2X2 U104 ( .A(\op<1> ), .B(\op<0> ), .Y(n99) );
  INVX1 U105 ( .A(n99), .Y(n100) );
  INVX1 U106 ( .A(n101), .Y(\out<7> ) );
  INVX1 U107 ( .A(n25), .Y(n103) );
  INVX1 U108 ( .A(n23), .Y(n104) );
  BUFX2 U109 ( .A(\in<0> ), .Y(n105) );
  INVX1 U110 ( .A(\in<15> ), .Y(n106) );
  INVX1 U111 ( .A(n106), .Y(n107) );
  INVX1 U112 ( .A(n89), .Y(n108) );
  INVX1 U113 ( .A(n108), .Y(n109) );
  INVX1 U114 ( .A(n105), .Y(n110) );
  INVX1 U115 ( .A(n110), .Y(n111) );
  INVX1 U116 ( .A(\op<2> ), .Y(n119) );
  INVX1 U117 ( .A(n87), .Y(n112) );
  INVX1 U118 ( .A(n112), .Y(n114) );
  OAI21X1 U119 ( .A(\op<0> ), .B(n115), .C(sh), .Y(n116) );
  INVX2 U120 ( .A(n116), .Y(n117) );
  AND2X2 U121 ( .A(\op<0> ), .B(sh), .Y(n118) );
  NAND3X1 U122 ( .A(n113), .B(n71), .C(n103), .Y(\out<8> ) );
  NAND3X1 U123 ( .A(n65), .B(n73), .C(n87), .Y(\out<9> ) );
  NAND3X1 U124 ( .A(n113), .B(n75), .C(n27), .Y(\out<10> ) );
  NAND3X1 U125 ( .A(n67), .B(n29), .C(n114), .Y(\out<11> ) );
  NAND3X1 U126 ( .A(n114), .B(n77), .C(n83), .Y(\out<12> ) );
  NAND3X1 U127 ( .A(n85), .B(n113), .C(n79), .Y(\out<13> ) );
  NAND3X1 U128 ( .A(n114), .B(n81), .C(n69), .Y(\out<14> ) );
endmodule


module cla_4_3 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3, n1, n2;

  fulladder_1_15 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(n2), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_14 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_13 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_12 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_3 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
  INVX1 U1 ( .A(Cin), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
endmodule


module cla_4_2 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3, n1;

  fulladder_1_11 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(n1), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_10 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_9 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_8 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_2 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
  BUFX2 U1 ( .A(Cin), .Y(n1) );
endmodule


module cla_4_1 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3, n1, n2;

  fulladder_1_7 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(n2), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_6 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_5 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_4 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_1 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
  INVX1 U1 ( .A(Cin), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
endmodule


module cla_4_0 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3;

  fulladder_1_3 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_2 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_1 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_0 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_0 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
endmodule


module groupcla_8 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37;

  AND2X1 U1 ( .A(n25), .B(n12), .Y(n13) );
  INVX2 U2 ( .A(n35), .Y(n34) );
  INVX1 U3 ( .A(n31), .Y(n1) );
  BUFX2 U4 ( .A(n36), .Y(n2) );
  AND2X2 U5 ( .A(\p<1> ), .B(n26), .Y(n3) );
  INVX1 U6 ( .A(n3), .Y(n4) );
  INVX1 U7 ( .A(n3), .Y(n5) );
  OR2X2 U8 ( .A(n23), .B(\g<0> ), .Y(n6) );
  INVX1 U9 ( .A(n6), .Y(n7) );
  INVX1 U10 ( .A(n6), .Y(n8) );
  INVX1 U11 ( .A(\p<3> ), .Y(n9) );
  INVX1 U12 ( .A(n9), .Y(n10) );
  INVX1 U13 ( .A(\g<1> ), .Y(n33) );
  AND2X2 U14 ( .A(n20), .B(n21), .Y(n11) );
  INVX1 U15 ( .A(n11), .Y(n12) );
  INVX1 U16 ( .A(n13), .Y(n14) );
  BUFX2 U17 ( .A(n29), .Y(n15) );
  AND2X1 U18 ( .A(n20), .B(n22), .Y(n16) );
  INVX1 U19 ( .A(n16), .Y(n17) );
  INVX1 U20 ( .A(n6), .Y(n18) );
  OAI21X1 U21 ( .A(n30), .B(n8), .C(n33), .Y(\c<1> ) );
  BUFX2 U22 ( .A(\g<3> ), .Y(n19) );
  INVX1 U23 ( .A(n30), .Y(n20) );
  BUFX2 U24 ( .A(\g<0> ), .Y(n21) );
  BUFX2 U25 ( .A(\p<0> ), .Y(n22) );
  INVX1 U26 ( .A(\p<1> ), .Y(n30) );
  INVX1 U27 ( .A(n7), .Y(\c<0> ) );
  AND2X2 U28 ( .A(\p<0> ), .B(Cin), .Y(n23) );
  INVX1 U29 ( .A(n26), .Y(n24) );
  INVX1 U30 ( .A(\p<2> ), .Y(n32) );
  BUFX2 U31 ( .A(n33), .Y(n25) );
  INVX1 U32 ( .A(n19), .Y(n28) );
  INVX1 U33 ( .A(n32), .Y(n26) );
  INVX1 U34 ( .A(n24), .Y(n27) );
  INVX1 U35 ( .A(\g<2> ), .Y(n31) );
  AOI21X1 U36 ( .A(n27), .B(n14), .C(n1), .Y(n29) );
  OAI21X1 U37 ( .A(n15), .B(n9), .C(n28), .Y(gg) );
  NOR3X1 U38 ( .A(n17), .B(n9), .C(n24), .Y(pg) );
  OAI21X1 U39 ( .A(n33), .B(n32), .C(n31), .Y(n35) );
  OAI21X1 U40 ( .A(n4), .B(n18), .C(n34), .Y(\c<2> ) );
  OAI21X1 U41 ( .A(n23), .B(n21), .C(\p<3> ), .Y(n37) );
  AOI21X1 U42 ( .A(n10), .B(n35), .C(\g<3> ), .Y(n36) );
  OAI21X1 U43 ( .A(n5), .B(n37), .C(n2), .Y(\c<3> ) );
endmodule


module fulladder_1_31 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_30 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;


  XOR2X1 U1 ( .A(A), .B(B), .Y(p) );
  XOR2X1 U2 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U3 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_29 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_28 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  AND2X2 U1 ( .A(A), .B(B), .Y(g) );
  XNOR2X1 U2 ( .A(A), .B(B), .Y(n1) );
  INVX2 U3 ( .A(n1), .Y(p) );
  XOR2X1 U4 ( .A(Cin), .B(p), .Y(S) );
endmodule


module groupcla_7 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n2, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n23, n24, n25;

  NOR3X1 U8 ( .A(n15), .B(n23), .C(n25), .Y(pg) );
  INVX1 U1 ( .A(\g<1> ), .Y(n18) );
  INVX1 U2 ( .A(\g<0> ), .Y(n17) );
  INVX1 U3 ( .A(\p<1> ), .Y(n19) );
  INVX1 U4 ( .A(\g<2> ), .Y(n20) );
  INVX1 U5 ( .A(\p<2> ), .Y(n23) );
  INVX1 U6 ( .A(\g<3> ), .Y(n24) );
  INVX1 U7 ( .A(\p<3> ), .Y(n25) );
  AND2X2 U9 ( .A(\p<0> ), .B(Cin), .Y(n1) );
  INVX1 U10 ( .A(n1), .Y(n2) );
  AND2X2 U11 ( .A(\p<2> ), .B(\c<1> ), .Y(n3) );
  INVX1 U12 ( .A(n3), .Y(n4) );
  AND2X2 U13 ( .A(n20), .B(n4), .Y(n5) );
  INVX1 U14 ( .A(n5), .Y(\c<2> ) );
  AND2X2 U15 ( .A(n17), .B(n2), .Y(n7) );
  INVX1 U16 ( .A(n7), .Y(\c<0> ) );
  AND2X2 U17 ( .A(\p<1> ), .B(\g<0> ), .Y(n9) );
  INVX1 U18 ( .A(n9), .Y(n10) );
  AND2X2 U19 ( .A(n18), .B(n10), .Y(n11) );
  INVX1 U20 ( .A(n11), .Y(n12) );
  BUFX2 U21 ( .A(n16), .Y(n13) );
  AND2X2 U22 ( .A(\p<1> ), .B(\p<0> ), .Y(n14) );
  INVX1 U23 ( .A(n14), .Y(n15) );
  INVX1 U24 ( .A(\c<2> ), .Y(n21) );
  AOI21X1 U25 ( .A(\p<2> ), .B(n12), .C(\g<2> ), .Y(n16) );
  OAI21X1 U26 ( .A(n13), .B(n25), .C(n24), .Y(gg) );
  OAI21X1 U27 ( .A(n7), .B(n19), .C(n18), .Y(\c<1> ) );
  OAI21X1 U28 ( .A(n21), .B(n25), .C(n24), .Y(\c<3> ) );
endmodule


module fulladder_1_27 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_26 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_25 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_24 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_6 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28;

  INVX1 U1 ( .A(\g<1> ), .Y(n23) );
  INVX1 U2 ( .A(\g<0> ), .Y(n22) );
  INVX1 U3 ( .A(\p<1> ), .Y(n24) );
  AND2X1 U4 ( .A(\p<1> ), .B(\g<0> ), .Y(n10) );
  INVX1 U5 ( .A(\g<2> ), .Y(n25) );
  INVX1 U6 ( .A(\g<3> ), .Y(n26) );
  INVX1 U7 ( .A(\p<3> ), .Y(n27) );
  AND2X2 U8 ( .A(n26), .B(n19), .Y(n1) );
  INVX1 U9 ( .A(n1), .Y(gg) );
  OR2X2 U10 ( .A(n21), .B(n14), .Y(n3) );
  INVX1 U11 ( .A(n3), .Y(pg) );
  AND2X2 U12 ( .A(n22), .B(n13), .Y(n5) );
  AND2X2 U13 ( .A(n23), .B(n11), .Y(n6) );
  INVX1 U14 ( .A(n6), .Y(n7) );
  AND2X2 U15 ( .A(\p<2> ), .B(\c<1> ), .Y(n8) );
  INVX1 U16 ( .A(n8), .Y(n9) );
  INVX1 U17 ( .A(n10), .Y(n11) );
  AND2X2 U18 ( .A(Cin), .B(\p<0> ), .Y(n12) );
  INVX1 U19 ( .A(n12), .Y(n13) );
  BUFX2 U20 ( .A(n20), .Y(n14) );
  AND2X2 U21 ( .A(n25), .B(n9), .Y(n15) );
  INVX1 U22 ( .A(n15), .Y(\c<2> ) );
  INVX1 U23 ( .A(n5), .Y(\c<0> ) );
  INVX1 U24 ( .A(\c<2> ), .Y(n28) );
  AND2X2 U25 ( .A(\p<2> ), .B(n7), .Y(n18) );
  OAI21X1 U26 ( .A(n18), .B(\g<2> ), .C(\p<3> ), .Y(n19) );
  INVX2 U27 ( .A(\p<2> ), .Y(n21) );
  NAND3X1 U28 ( .A(\p<0> ), .B(\p<1> ), .C(\p<3> ), .Y(n20) );
  OAI21X1 U29 ( .A(n5), .B(n24), .C(n23), .Y(\c<1> ) );
  OAI21X1 U30 ( .A(n28), .B(n27), .C(n26), .Y(\c<3> ) );
endmodule


module fulladder_1_23 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_22 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_21 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_20 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;


  XOR2X1 U1 ( .A(A), .B(B), .Y(p) );
  XOR2X1 U2 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U3 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_5 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n15, n16, n17, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  INVX1 U1 ( .A(\p<2> ), .Y(n19) );
  INVX1 U2 ( .A(\g<0> ), .Y(n23) );
  INVX1 U3 ( .A(\g<2> ), .Y(n26) );
  INVX1 U4 ( .A(\g<1> ), .Y(n24) );
  INVX1 U5 ( .A(\p<1> ), .Y(n25) );
  INVX1 U6 ( .A(\g<3> ), .Y(n27) );
  AND2X2 U7 ( .A(n27), .B(n8), .Y(n1) );
  INVX1 U8 ( .A(n1), .Y(gg) );
  AND2X2 U9 ( .A(Cin), .B(\p<0> ), .Y(n3) );
  INVX1 U10 ( .A(n3), .Y(n4) );
  AND2X2 U11 ( .A(\p<2> ), .B(\c<1> ), .Y(n5) );
  INVX1 U12 ( .A(n5), .Y(n6) );
  AND2X2 U13 ( .A(\p<3> ), .B(n21), .Y(n7) );
  INVX1 U14 ( .A(n7), .Y(n8) );
  BUFX2 U15 ( .A(n20), .Y(n9) );
  AND2X2 U16 ( .A(n26), .B(n6), .Y(n10) );
  INVX1 U17 ( .A(n10), .Y(\c<2> ) );
  INVX1 U18 ( .A(n10), .Y(n12) );
  AND2X2 U19 ( .A(n23), .B(n4), .Y(n13) );
  INVX1 U20 ( .A(n13), .Y(\c<0> ) );
  INVX1 U21 ( .A(n22), .Y(n15) );
  INVX1 U22 ( .A(n15), .Y(n16) );
  INVX1 U23 ( .A(n12), .Y(n29) );
  OR2X2 U24 ( .A(n28), .B(n16), .Y(n17) );
  INVX1 U25 ( .A(n17), .Y(pg) );
  AOI21X1 U26 ( .A(\p<1> ), .B(\g<0> ), .C(\g<1> ), .Y(n20) );
  OAI21X1 U27 ( .A(n9), .B(n19), .C(n26), .Y(n21) );
  INVX2 U28 ( .A(\p<3> ), .Y(n28) );
  NAND3X1 U29 ( .A(\p<0> ), .B(\p<1> ), .C(\p<2> ), .Y(n22) );
  OAI21X1 U30 ( .A(n13), .B(n25), .C(n24), .Y(\c<1> ) );
  OAI21X1 U31 ( .A(n29), .B(n28), .C(n27), .Y(\c<3> ) );
endmodule


module fulladder_1_19 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1, n2;

  INVX1 U1 ( .A(Cin), .Y(n2) );
  INVX1 U2 ( .A(n1), .Y(p) );
  XNOR2X1 U3 ( .A(A), .B(B), .Y(n1) );
  XNOR2X1 U4 ( .A(p), .B(n2), .Y(S) );
  AND2X2 U5 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_18 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_17 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module fulladder_1_16 ( A, B, Cin, p, g, S );
  input A, B, Cin;
  output p, g, S;
  wire   n1;

  XNOR2X1 U1 ( .A(A), .B(B), .Y(n1) );
  INVX2 U2 ( .A(n1), .Y(p) );
  XOR2X1 U3 ( .A(Cin), .B(p), .Y(S) );
  AND2X2 U4 ( .A(A), .B(B), .Y(g) );
endmodule


module groupcla_4 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n22, n23, n24, n25;

  INVX1 U1 ( .A(\g<0> ), .Y(n20) );
  INVX1 U2 ( .A(\p<2> ), .Y(n19) );
  INVX1 U3 ( .A(\g<2> ), .Y(n23) );
  INVX1 U4 ( .A(\g<1> ), .Y(n21) );
  INVX1 U5 ( .A(\p<1> ), .Y(n22) );
  INVX1 U6 ( .A(\g<3> ), .Y(n24) );
  INVX1 U7 ( .A(\p<3> ), .Y(n25) );
  AND2X2 U8 ( .A(n24), .B(n12), .Y(n1) );
  INVX1 U9 ( .A(n1), .Y(gg) );
  AND2X2 U10 ( .A(\p<0> ), .B(\p<1> ), .Y(n3) );
  INVX1 U11 ( .A(n3), .Y(n4) );
  AND2X2 U12 ( .A(Cin), .B(\p<0> ), .Y(n5) );
  INVX1 U13 ( .A(n5), .Y(n6) );
  AND2X2 U14 ( .A(\p<2> ), .B(\c<1> ), .Y(n7) );
  INVX1 U15 ( .A(n7), .Y(n8) );
  AND2X2 U16 ( .A(n23), .B(n8), .Y(n9) );
  INVX1 U17 ( .A(n9), .Y(\c<2> ) );
  AND2X2 U18 ( .A(\p<3> ), .B(n18), .Y(n11) );
  INVX1 U19 ( .A(n11), .Y(n12) );
  AND2X2 U20 ( .A(n20), .B(n6), .Y(n13) );
  INVX1 U21 ( .A(n17), .Y(n14) );
  INVX1 U22 ( .A(n14), .Y(n15) );
  INVX1 U23 ( .A(n13), .Y(\c<0> ) );
  AOI21X1 U24 ( .A(\p<1> ), .B(\g<0> ), .C(\g<1> ), .Y(n17) );
  OAI21X1 U25 ( .A(n15), .B(n19), .C(n23), .Y(n18) );
  NOR3X1 U26 ( .A(n4), .B(n19), .C(n25), .Y(pg) );
  OAI21X1 U27 ( .A(n13), .B(n22), .C(n21), .Y(\c<1> ) );
  OAI21X1 U28 ( .A(n9), .B(n25), .C(n24), .Y(\c<3> ) );
endmodule


module cla_4_11 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3, n1, n2, n3;

  fulladder_1_47 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(n3), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_46 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_45 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_44 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_12 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(n1), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
  BUFX2 U1 ( .A(Cin), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
endmodule


module cla_4_10 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3;

  fulladder_1_43 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_42 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_41 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_40 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_11 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c(
        {Cout, c3, c2, c1}), .pg(p), .gg(g) );
endmodule


module cla_4_9 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3;

  fulladder_1_39 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_38 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_37 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_36 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_10 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c(
        {Cout, c3, c2, c1}), .pg(p), .gg(g) );
endmodule


module cla_4_8 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3;

  fulladder_1_35 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_34 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_33 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_32 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_9 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
endmodule


module groupcla_14 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28;

  NOR3X1 U8 ( .A(n19), .B(n26), .C(n28), .Y(pg) );
  AND2X2 U1 ( .A(n24), .B(n3), .Y(n8) );
  INVX1 U2 ( .A(\c<0> ), .Y(n23) );
  INVX1 U3 ( .A(\g<3> ), .Y(n27) );
  INVX1 U4 ( .A(\p<2> ), .Y(n26) );
  INVX1 U5 ( .A(\p<3> ), .Y(n28) );
  INVX1 U6 ( .A(n8), .Y(\c<2> ) );
  AND2X2 U7 ( .A(\p<2> ), .B(\c<1> ), .Y(n2) );
  INVX1 U9 ( .A(n2), .Y(n3) );
  INVX1 U10 ( .A(n22), .Y(n4) );
  INVX1 U11 ( .A(n17), .Y(n5) );
  INVX1 U12 ( .A(\g<1> ), .Y(n22) );
  AND2X1 U13 ( .A(n14), .B(n10), .Y(n6) );
  INVX1 U14 ( .A(n6), .Y(n7) );
  AND2X1 U15 ( .A(n15), .B(n17), .Y(n9) );
  INVX1 U16 ( .A(n9), .Y(n10) );
  AND2X1 U17 ( .A(\p<3> ), .B(n20), .Y(n11) );
  INVX1 U18 ( .A(n11), .Y(n12) );
  AND2X1 U19 ( .A(n15), .B(n16), .Y(n13) );
  INVX1 U20 ( .A(n13), .Y(n14) );
  INVX1 U21 ( .A(n21), .Y(\c<0> ) );
  INVX1 U22 ( .A(n4), .Y(n15) );
  INVX1 U23 ( .A(\g<0> ), .Y(n16) );
  INVX1 U24 ( .A(\p<1> ), .Y(n17) );
  AND2X2 U25 ( .A(n5), .B(\p<0> ), .Y(n18) );
  INVX1 U26 ( .A(n18), .Y(n19) );
  INVX2 U27 ( .A(\g<2> ), .Y(n24) );
  OAI21X1 U28 ( .A(n7), .B(n26), .C(n24), .Y(n20) );
  NAND2X1 U29 ( .A(n27), .B(n12), .Y(gg) );
  AOI21X1 U30 ( .A(\p<0> ), .B(Cin), .C(\g<0> ), .Y(n21) );
  OAI21X1 U31 ( .A(n23), .B(n17), .C(n22), .Y(\c<1> ) );
  OAI21X1 U32 ( .A(n8), .B(n28), .C(n27), .Y(\c<3> ) );
endmodule


module register_7 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_112 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(n1) );
  dff_113 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(n1) );
  dff_114 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(rst) );
  dff_115 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(rst) );
  dff_116 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_117 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_118 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_119 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_120 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_121 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_122 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_123 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_124 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_125 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_126 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_127 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module register_6 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_111 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(n1) );
  dff_110 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(rst) );
  dff_109 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(rst) );
  dff_108 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(rst) );
  dff_107 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_106 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_105 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_104 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_103 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_102 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_101 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_100 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_99 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_98 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_97 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_96 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module register_5 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_95 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(rst) );
  dff_94 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(n1) );
  dff_93 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(rst) );
  dff_92 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(rst) );
  dff_91 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_90 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_89 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_88 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_87 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_86 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_85 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_84 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_83 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_82 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_81 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_80 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module register_4 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_79 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(n1) );
  dff_78 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(n1) );
  dff_77 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(rst) );
  dff_76 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(rst) );
  dff_75 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_74 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_73 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_72 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_71 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_70 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_69 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_68 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_67 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_66 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_65 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_64 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module register_3 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_63 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(n1) );
  dff_62 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(n1) );
  dff_61 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(rst) );
  dff_60 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(rst) );
  dff_59 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_58 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_57 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_56 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_55 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_54 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_53 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_52 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_51 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_50 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_49 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_48 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module register_2 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_47 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(rst) );
  dff_46 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(rst) );
  dff_45 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(rst) );
  dff_44 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(n1) );
  dff_43 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_42 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_41 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_40 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_39 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_38 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_37 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_36 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_35 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_34 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_33 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_32 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module register_1 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_31 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(rst) );
  dff_30 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(rst) );
  dff_29 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(n1) );
  dff_28 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(n1) );
  dff_27 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_26 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_25 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_24 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_23 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_22 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_21 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_20 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_19 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_18 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_17 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_16 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module register_0 ( .in({\in<15> , \in<14> , \in<13> , \in<12> , \in<11> , 
        \in<10> , \in<9> , \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , 
        \in<3> , \in<2> , \in<1> , \in<0> }), clk, rst, .out({\out<15> , 
        \out<14> , \out<13> , \out<12> , \out<11> , \out<10> , \out<9> , 
        \out<8> , \out<7> , \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , 
        \out<1> , \out<0> }) );
  input \in<15> , \in<14> , \in<13> , \in<12> , \in<11> , \in<10> , \in<9> ,
         \in<8> , \in<7> , \in<6> , \in<5> , \in<4> , \in<3> , \in<2> ,
         \in<1> , \in<0> , clk, rst, \out<15> , \out<14> , \out<13> ,
         \out<12> , \out<11> , \out<10> , \out<9> , \out<8> , \out<7> ,
         \out<6> , \out<5> , \out<4> , \out<3> , \out<2> , \out<1> , \out<0> ;
  wire   n1, n2;

  dff_15 \val[0]  ( .q(), .d(\in<0> ), .clk(clk), .rst(rst) );
  dff_14 \val[1]  ( .q(), .d(\in<1> ), .clk(clk), .rst(n1) );
  dff_13 \val[2]  ( .q(), .d(\in<2> ), .clk(clk), .rst(rst) );
  dff_12 \val[3]  ( .q(), .d(\in<3> ), .clk(clk), .rst(rst) );
  dff_11 \val[4]  ( .q(), .d(\in<4> ), .clk(clk), .rst(n1) );
  dff_10 \val[5]  ( .q(), .d(\in<5> ), .clk(clk), .rst(n1) );
  dff_9 \val[6]  ( .q(), .d(\in<6> ), .clk(clk), .rst(n1) );
  dff_8 \val[7]  ( .q(), .d(\in<7> ), .clk(clk), .rst(n1) );
  dff_7 \val[8]  ( .q(), .d(\in<8> ), .clk(clk), .rst(n1) );
  dff_6 \val[9]  ( .q(), .d(\in<9> ), .clk(clk), .rst(n1) );
  dff_5 \val[10]  ( .q(), .d(\in<10> ), .clk(clk), .rst(n1) );
  dff_4 \val[11]  ( .q(), .d(\in<11> ), .clk(clk), .rst(n1) );
  dff_3 \val[12]  ( .q(), .d(\in<12> ), .clk(clk), .rst(n1) );
  dff_2 \val[13]  ( .q(), .d(\in<13> ), .clk(clk), .rst(n1) );
  dff_1 \val[14]  ( .q(), .d(\in<14> ), .clk(clk), .rst(n1) );
  dff_0 \val[15]  ( .q(), .d(\in<15> ), .clk(clk), .rst(n1) );
  INVX1 U1 ( .A(rst), .Y(n2) );
  INVX1 U2 ( .A(n2), .Y(n1) );
endmodule


module shifter ( .In({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .Cnt({\Cnt<3> , \Cnt<2> , 
        \Cnt<1> , \Cnt<0> }), .Op({\Op<2> , \Op<1> , \Op<0> }), .Out({
        \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> , 
        \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> , 
        \Out<2> , \Out<1> , \Out<0> }) );
  input \In<15> , \In<14> , \In<13> , \In<12> , \In<11> , \In<10> , \In<9> ,
         \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , \In<3> , \In<2> ,
         \In<1> , \In<0> , \Cnt<3> , \Cnt<2> , \Cnt<1> , \Cnt<0> , \Op<2> ,
         \Op<1> , \Op<0> ;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> ;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, \sh1<15> ,
         \sh1<14> , \sh1<13> , \sh1<12> , \sh1<11> , \sh1<10> , \sh1<9> ,
         \sh1<8> , \sh1<7> , \sh1<6> , \sh1<5> , \sh1<4> , \sh1<3> , \sh1<2> ,
         \sh1<1> , \sh1<0> , \sh2<15> , \sh2<14> , \sh2<13> , \sh2<12> ,
         \sh2<11> , \sh2<10> , \sh2<9> , \sh2<8> , \sh2<7> , \sh2<6> ,
         \sh2<5> , \sh2<4> , \sh2<3> , \sh2<2> , \sh2<1> , \sh2<0> , \sh3<15> ,
         \sh3<14> , \sh3<13> , \sh3<12> , \sh3<11> , \sh3<10> , \sh3<9> ,
         \sh3<8> , \sh3<7> , \sh3<6> , \sh3<5> , \sh3<4> , \sh3<3> , \sh3<2> ,
         \sh3<1> , \sh3<0> , n1, n2, n13, n14;

  shifter_1 sh_1 ( .in({\In<15> , \In<14> , \In<13> , \In<12> , \In<11> , 
        \In<10> , \In<9> , \In<8> , \In<7> , \In<6> , \In<5> , \In<4> , 
        \In<3> , \In<2> , \In<1> , \In<0> }), .op({\Op<2> , \Op<1> , \Op<0> }), 
        .sh(\Cnt<0> ), .out({\sh1<15> , \sh1<14> , \sh1<13> , \sh1<12> , 
        \sh1<11> , \sh1<10> , \sh1<9> , \sh1<8> , \sh1<7> , \sh1<6> , \sh1<5> , 
        \sh1<4> , \sh1<3> , \sh1<2> , \sh1<1> , \sh1<0> }) );
  shifter_2 sh_2 ( .in({\sh1<15> , \sh1<14> , \sh1<13> , \sh1<12> , \sh1<11> , 
        \sh1<10> , \sh1<9> , \sh1<8> , \sh1<7> , \sh1<6> , \sh1<5> , \sh1<4> , 
        \sh1<3> , \sh1<2> , \sh1<1> , \sh1<0> }), .op({n1, \Op<1> , n2}), .sh(
        \Cnt<1> ), .out({\sh2<15> , \sh2<14> , \sh2<13> , \sh2<12> , \sh2<11> , 
        \sh2<10> , \sh2<9> , \sh2<8> , \sh2<7> , \sh2<6> , \sh2<5> , \sh2<4> , 
        \sh2<3> , \sh2<2> , \sh2<1> , \sh2<0> }) );
  shifter_4 sh_4 ( .in({\sh2<15> , \sh2<14> , \sh2<13> , \sh2<12> , \sh2<11> , 
        \sh2<10> , \sh2<9> , \sh2<8> , \sh2<7> , \sh2<6> , \sh2<5> , \sh2<4> , 
        \sh2<3> , \sh2<2> , \sh2<1> , \sh2<0> }), .op({n14, \Op<1> , n2}), 
        .sh(\Cnt<2> ), .out({\sh3<15> , \sh3<14> , \sh3<13> , \sh3<12> , 
        \sh3<11> , \sh3<10> , \sh3<9> , \sh3<8> , \sh3<7> , \sh3<6> , \sh3<5> , 
        \sh3<4> , \sh3<3> , \sh3<2> , \sh3<1> , \sh3<0> }) );
  shifter_8 sh_8 ( .in({\sh3<15> , \sh3<14> , \sh3<13> , \sh3<12> , \sh3<11> , 
        \sh3<10> , \sh3<9> , \sh3<8> , \sh3<7> , \sh3<6> , \sh3<5> , \sh3<4> , 
        \sh3<3> , \sh3<2> , \sh3<1> , \sh3<0> }), .op({n14, \Op<1> , n2}), 
        .sh(\Cnt<3> ), .out({n15, n16, n17, n18, n19, n20, n21, n22, \Out<7> , 
        \Out<6> , n23, \Out<4> , n24, \Out<2> , \Out<1> , \Out<0> }) );
  INVX1 U1 ( .A(n13), .Y(n1) );
  BUFX2 U2 ( .A(\Op<0> ), .Y(n2) );
  BUFX2 U3 ( .A(n23), .Y(\Out<5> ) );
  BUFX2 U4 ( .A(n17), .Y(\Out<13> ) );
  BUFX2 U5 ( .A(n24), .Y(\Out<3> ) );
  BUFX2 U6 ( .A(n21), .Y(\Out<9> ) );
  BUFX2 U7 ( .A(n20), .Y(\Out<10> ) );
  BUFX2 U8 ( .A(n16), .Y(\Out<14> ) );
  BUFX2 U9 ( .A(n15), .Y(\Out<15> ) );
  BUFX2 U10 ( .A(n22), .Y(\Out<8> ) );
  BUFX2 U11 ( .A(n19), .Y(\Out<11> ) );
  BUFX2 U12 ( .A(n18), .Y(\Out<12> ) );
  INVX1 U13 ( .A(\Op<2> ), .Y(n13) );
  INVX1 U14 ( .A(n13), .Y(n14) );
endmodule


module adder_0 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Overflow, Cout, .Sum({\Sum<15> , \Sum<14> , \Sum<13> , 
        \Sum<12> , \Sum<11> , \Sum<10> , \Sum<9> , \Sum<8> , \Sum<7> , 
        \Sum<6> , \Sum<5> , \Sum<4> , \Sum<3> , \Sum<2> , \Sum<1> , \Sum<0> })
 );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Overflow, Cout, \Sum<15> , \Sum<14> , \Sum<13> , \Sum<12> , \Sum<11> ,
         \Sum<10> , \Sum<9> , \Sum<8> , \Sum<7> , \Sum<6> , \Sum<5> , \Sum<4> ,
         \Sum<3> , \Sum<2> , \Sum<1> , \Sum<0> ;
  wire   c12, p12, g12, c8, p8, g8, c4, p4, g4, p0, g0, n2, n3, n4, n5;

  FAX1 U1 ( .A(n2), .B(\A<15> ), .C(n5), .YC(), .YS(Overflow) );
  XOR2X1 U2 ( .A(n3), .B(n4), .Y(n5) );
  cla_4_3 add1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(c12), .p(p12), .g(g12), .S({
        \Sum<15> , \Sum<14> , \Sum<13> , \Sum<12> }), .Cout() );
  cla_4_2 add2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(c8), .p(p8), .g(g8), .S({\Sum<11> , \Sum<10> , 
        \Sum<9> , \Sum<8> }), .Cout() );
  cla_4_1 add3 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(c4), .p(p4), .g(g4), .S({\Sum<7> , \Sum<6> , 
        \Sum<5> , \Sum<4> }), .Cout() );
  cla_4_0 add4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .p(p0), .g(g0), .S({\Sum<3> , \Sum<2> , 
        \Sum<1> , \Sum<0> }), .Cout() );
  groupcla_8 cla ( .p({p12, p8, p4, p0}), .g({g12, g8, g4, g0}), .Cin(Cin), 
        .c({Cout, c12, c8, c4}), .pg(), .gg() );
  BUFX2 U3 ( .A(\B<15> ), .Y(n2) );
  BUFX2 U4 ( .A(\Sum<15> ), .Y(n3) );
  BUFX2 U5 ( .A(Cout), .Y(n4) );
endmodule


module cla_4_7 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3, n1, n2, n3;

  fulladder_1_31 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(n3), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_30 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_29 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_28 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_7 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(n1), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
  BUFX2 U1 ( .A(Cin), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(n2) );
  INVX1 U3 ( .A(n2), .Y(n3) );
endmodule


module cla_4_6 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3;

  fulladder_1_27 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_26 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_25 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_24 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_6 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
endmodule


module cla_4_5 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3;

  fulladder_1_23 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_22 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_21 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_20 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_5 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
endmodule


module cla_4_4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), Cin, p, g, .S({\S<3> , \S<2> , \S<1> , \S<0> }), 
        Cout );
  input \A<3> , \A<2> , \A<1> , \A<0> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output p, g, \S<3> , \S<2> , \S<1> , \S<0> , Cout;
  wire   p0, g0, c1, p1, g1, c2, p2, g2, c3, p3, g3;

  fulladder_1_19 fa1 ( .A(\A<0> ), .B(\B<0> ), .Cin(Cin), .p(p0), .g(g0), .S(
        \S<0> ) );
  fulladder_1_18 fa2 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .p(p1), .g(g1), .S(
        \S<1> ) );
  fulladder_1_17 fa3 ( .A(\A<2> ), .B(\B<2> ), .Cin(c2), .p(p2), .g(g2), .S(
        \S<2> ) );
  fulladder_1_16 fa4 ( .A(\A<3> ), .B(\B<3> ), .Cin(c3), .p(p3), .g(g3), .S(
        \S<3> ) );
  groupcla_4 cla ( .p({p3, p2, p1, p0}), .g({g3, g2, g1, g0}), .Cin(Cin), .c({
        Cout, c3, c2, c1}), .pg(p), .gg(g) );
endmodule


module groupcla_13 ( .p({\p<3> , \p<2> , \p<1> , \p<0> }), .g({\g<3> , \g<2> , 
        \g<1> , \g<0> }), Cin, .c({\c<3> , \c<2> , \c<1> , \c<0> }), pg, gg );
  input \p<3> , \p<2> , \p<1> , \p<0> , \g<3> , \g<2> , \g<1> , \g<0> , Cin;
  output \c<3> , \c<2> , \c<1> , \c<0> , pg, gg;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n24;

  NOR3X1 U8 ( .A(n14), .B(n12), .C(n24), .Y(pg) );
  INVX1 U1 ( .A(\g<3> ), .Y(n23) );
  INVX1 U2 ( .A(\p<3> ), .Y(n24) );
  AND2X2 U3 ( .A(n21), .B(n16), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(\c<2> ) );
  BUFX2 U5 ( .A(n21), .Y(n3) );
  INVX1 U6 ( .A(\g<2> ), .Y(n21) );
  BUFX2 U7 ( .A(\g<0> ), .Y(n4) );
  AND2X1 U9 ( .A(n10), .B(n8), .Y(n5) );
  INVX1 U10 ( .A(n5), .Y(n6) );
  AND2X1 U11 ( .A(n3), .B(n12), .Y(n7) );
  INVX1 U12 ( .A(n7), .Y(n8) );
  AND2X1 U13 ( .A(n3), .B(n11), .Y(n9) );
  INVX1 U14 ( .A(n9), .Y(n10) );
  INVX1 U15 ( .A(n19), .Y(\c<0> ) );
  INVX1 U16 ( .A(n20), .Y(\c<1> ) );
  INVX1 U17 ( .A(n18), .Y(n11) );
  INVX1 U18 ( .A(\p<2> ), .Y(n12) );
  INVX1 U19 ( .A(n17), .Y(n18) );
  AND2X2 U20 ( .A(\p<1> ), .B(\p<0> ), .Y(n13) );
  INVX1 U21 ( .A(n13), .Y(n14) );
  AND2X2 U22 ( .A(\p<2> ), .B(\c<1> ), .Y(n15) );
  INVX1 U23 ( .A(n15), .Y(n16) );
  AOI21X1 U24 ( .A(\p<1> ), .B(n4), .C(\g<1> ), .Y(n17) );
  OAI21X1 U25 ( .A(n6), .B(n24), .C(n23), .Y(gg) );
  AOI21X1 U26 ( .A(\p<0> ), .B(Cin), .C(\g<0> ), .Y(n19) );
  AOI21X1 U27 ( .A(\p<1> ), .B(\c<0> ), .C(\g<1> ), .Y(n20) );
  OAI21X1 U28 ( .A(n1), .B(n24), .C(n23), .Y(\c<3> ) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module memory2c_1 ( .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), .addr({
        \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , 
        \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), enable, wr, createdump, 
        clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<15> , \addr<14> ,
         \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> ,
         \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , enable, wr, createdump, clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N177, N178, N179, N180, N181, N182, \mem<0><7> , \mem<0><6> ,
         \mem<0><5> , \mem<0><4> , \mem<0><3> , \mem<0><2> , \mem<0><1> ,
         \mem<0><0> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><7> ,
         \mem<2><6> , \mem<2><5> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><7> , \mem<3><6> , \mem<3><5> ,
         \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> , \mem<3><0> ,
         \mem<4><7> , \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> ,
         \mem<4><2> , \mem<4><1> , \mem<4><0> , \mem<5><7> , \mem<5><6> ,
         \mem<5><5> , \mem<5><4> , \mem<5><3> , \mem<5><2> , \mem<5><1> ,
         \mem<5><0> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><7> ,
         \mem<7><6> , \mem<7><5> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><7> , \mem<8><6> , \mem<8><5> ,
         \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> , \mem<8><0> ,
         \mem<9><7> , \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> ,
         \mem<9><2> , \mem<9><1> , \mem<9><0> , \mem<10><7> , \mem<10><6> ,
         \mem<10><5> , \mem<10><4> , \mem<10><3> , \mem<10><2> , \mem<10><1> ,
         \mem<10><0> , \mem<11><7> , \mem<11><6> , \mem<11><5> , \mem<11><4> ,
         \mem<11><3> , \mem<11><2> , \mem<11><1> , \mem<11><0> , \mem<12><7> ,
         \mem<12><6> , \mem<12><5> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><7> , \mem<13><6> , \mem<13><5> ,
         \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> , \mem<13><0> ,
         \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> , \mem<14><3> ,
         \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><7> ,
         \mem<17><6> , \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><7> , \mem<18><6> , \mem<18><5> ,
         \mem<18><4> , \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> ,
         \mem<19><7> , \mem<19><6> , \mem<19><5> , \mem<19><4> , \mem<19><3> ,
         \mem<19><2> , \mem<19><1> , \mem<19><0> , \mem<20><7> , \mem<20><6> ,
         \mem<20><5> , \mem<20><4> , \mem<20><3> , \mem<20><2> , \mem<20><1> ,
         \mem<20><0> , \mem<21><7> , \mem<21><6> , \mem<21><5> , \mem<21><4> ,
         \mem<21><3> , \mem<21><2> , \mem<21><1> , \mem<21><0> , \mem<22><7> ,
         \mem<22><6> , \mem<22><5> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><7> , \mem<23><6> , \mem<23><5> ,
         \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> , \mem<23><0> ,
         \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> , \mem<24><3> ,
         \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><7> ,
         \mem<27><6> , \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><7> , \mem<28><6> , \mem<28><5> ,
         \mem<28><4> , \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> ,
         \mem<29><7> , \mem<29><6> , \mem<29><5> , \mem<29><4> , \mem<29><3> ,
         \mem<29><2> , \mem<29><1> , \mem<29><0> , \mem<30><7> , \mem<30><6> ,
         \mem<30><5> , \mem<30><4> , \mem<30><3> , \mem<30><2> , \mem<30><1> ,
         \mem<30><0> , \mem<31><7> , \mem<31><6> , \mem<31><5> , \mem<31><4> ,
         \mem<31><3> , \mem<31><2> , \mem<31><1> , \mem<31><0> , \mem<32><7> ,
         \mem<32><6> , \mem<32><5> , \mem<32><4> , \mem<32><3> , \mem<32><2> ,
         \mem<32><1> , \mem<32><0> , \mem<33><7> , \mem<33><6> , \mem<33><5> ,
         \mem<33><4> , \mem<33><3> , \mem<33><2> , \mem<33><1> , \mem<33><0> ,
         \mem<34><7> , \mem<34><6> , \mem<34><5> , \mem<34><4> , \mem<34><3> ,
         \mem<34><2> , \mem<34><1> , \mem<34><0> , \mem<35><7> , \mem<35><6> ,
         \mem<35><5> , \mem<35><4> , \mem<35><3> , \mem<35><2> , \mem<35><1> ,
         \mem<35><0> , \mem<36><7> , \mem<36><6> , \mem<36><5> , \mem<36><4> ,
         \mem<36><3> , \mem<36><2> , \mem<36><1> , \mem<36><0> , \mem<37><7> ,
         \mem<37><6> , \mem<37><5> , \mem<37><4> , \mem<37><3> , \mem<37><2> ,
         \mem<37><1> , \mem<37><0> , \mem<38><7> , \mem<38><6> , \mem<38><5> ,
         \mem<38><4> , \mem<38><3> , \mem<38><2> , \mem<38><1> , \mem<38><0> ,
         \mem<39><7> , \mem<39><6> , \mem<39><5> , \mem<39><4> , \mem<39><3> ,
         \mem<39><2> , \mem<39><1> , \mem<39><0> , \mem<40><7> , \mem<40><6> ,
         \mem<40><5> , \mem<40><4> , \mem<40><3> , \mem<40><2> , \mem<40><1> ,
         \mem<40><0> , \mem<41><7> , \mem<41><6> , \mem<41><5> , \mem<41><4> ,
         \mem<41><3> , \mem<41><2> , \mem<41><1> , \mem<41><0> , \mem<42><7> ,
         \mem<42><6> , \mem<42><5> , \mem<42><4> , \mem<42><3> , \mem<42><2> ,
         \mem<42><1> , \mem<42><0> , \mem<43><7> , \mem<43><6> , \mem<43><5> ,
         \mem<43><4> , \mem<43><3> , \mem<43><2> , \mem<43><1> , \mem<43><0> ,
         \mem<44><7> , \mem<44><6> , \mem<44><5> , \mem<44><4> , \mem<44><3> ,
         \mem<44><2> , \mem<44><1> , \mem<44><0> , \mem<45><7> , \mem<45><6> ,
         \mem<45><5> , \mem<45><4> , \mem<45><3> , \mem<45><2> , \mem<45><1> ,
         \mem<45><0> , \mem<46><7> , \mem<46><6> , \mem<46><5> , \mem<46><4> ,
         \mem<46><3> , \mem<46><2> , \mem<46><1> , \mem<46><0> , \mem<47><7> ,
         \mem<47><6> , \mem<47><5> , \mem<47><4> , \mem<47><3> , \mem<47><2> ,
         \mem<47><1> , \mem<47><0> , \mem<48><7> , \mem<48><6> , \mem<48><5> ,
         \mem<48><4> , \mem<48><3> , \mem<48><2> , \mem<48><1> , \mem<48><0> ,
         \mem<49><7> , \mem<49><6> , \mem<49><5> , \mem<49><4> , \mem<49><3> ,
         \mem<49><2> , \mem<49><1> , \mem<49><0> , \mem<50><7> , \mem<50><6> ,
         \mem<50><5> , \mem<50><4> , \mem<50><3> , \mem<50><2> , \mem<50><1> ,
         \mem<50><0> , \mem<51><7> , \mem<51><6> , \mem<51><5> , \mem<51><4> ,
         \mem<51><3> , \mem<51><2> , \mem<51><1> , \mem<51><0> , \mem<52><7> ,
         \mem<52><6> , \mem<52><5> , \mem<52><4> , \mem<52><3> , \mem<52><2> ,
         \mem<52><1> , \mem<52><0> , \mem<53><7> , \mem<53><6> , \mem<53><5> ,
         \mem<53><4> , \mem<53><3> , \mem<53><2> , \mem<53><1> , \mem<53><0> ,
         \mem<54><7> , \mem<54><6> , \mem<54><5> , \mem<54><4> , \mem<54><3> ,
         \mem<54><2> , \mem<54><1> , \mem<54><0> , \mem<55><7> , \mem<55><6> ,
         \mem<55><5> , \mem<55><4> , \mem<55><3> , \mem<55><2> , \mem<55><1> ,
         \mem<55><0> , \mem<56><7> , \mem<56><6> , \mem<56><5> , \mem<56><4> ,
         \mem<56><3> , \mem<56><2> , \mem<56><1> , \mem<56><0> , \mem<57><7> ,
         \mem<57><6> , \mem<57><5> , \mem<57><4> , \mem<57><3> , \mem<57><2> ,
         \mem<57><1> , \mem<57><0> , \mem<58><7> , \mem<58><6> , \mem<58><5> ,
         \mem<58><4> , \mem<58><3> , \mem<58><2> , \mem<58><1> , \mem<58><0> ,
         \mem<59><7> , \mem<59><6> , \mem<59><5> , \mem<59><4> , \mem<59><3> ,
         \mem<59><2> , \mem<59><1> , \mem<59><0> , \mem<60><7> , \mem<60><6> ,
         \mem<60><5> , \mem<60><4> , \mem<60><3> , \mem<60><2> , \mem<60><1> ,
         \mem<60><0> , \mem<61><7> , \mem<61><6> , \mem<61><5> , \mem<61><4> ,
         \mem<61><3> , \mem<61><2> , \mem<61><1> , \mem<61><0> , \mem<62><7> ,
         \mem<62><6> , \mem<62><5> , \mem<62><4> , \mem<62><3> , \mem<62><2> ,
         \mem<62><1> , \mem<62><0> , \mem<63><7> , \mem<63><6> , \mem<63><5> ,
         \mem<63><4> , \mem<63><3> , \mem<63><2> , \mem<63><1> , \mem<63><0> ,
         n599, n602, n603, n604, n605, n606, n607, n608, n625, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n600, n601, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007;
  assign N177 = \addr<0> ;
  assign N178 = \addr<1> ;
  assign N179 = \addr<2> ;
  assign N180 = \addr<3> ;
  assign N181 = \addr<4> ;
  assign N182 = \addr<5> ;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n2327), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2326), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2325), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2324), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2323), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2322), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2321), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2320), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2319), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2318), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2317), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2316), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2315), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2314), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2313), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2312), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2311), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2310), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2309), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2308), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2307), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2306), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2305), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2304), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2303), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2302), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2301), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2300), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2299), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2298), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2297), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2296), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2295), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2294), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2293), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2292), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2291), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2290), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2289), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2288), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2287), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2286), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2285), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2284), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2283), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2282), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2281), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2280), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2279), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2278), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2277), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2276), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2275), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2274), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2273), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2272), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2271), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2270), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2269), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2268), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2267), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2266), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2265), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2264), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2263), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2262), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2261), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2260), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2259), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2258), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2257), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2256), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2255), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2254), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2253), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2252), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2251), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2250), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2249), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2248), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2247), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2246), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2245), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2244), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2243), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2242), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2241), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2240), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2239), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2238), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2237), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2236), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2235), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2234), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2233), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2232), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2231), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2230), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2229), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2228), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2227), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2226), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2225), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2224), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2223), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2222), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2221), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2220), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2219), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2218), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2217), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2216), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2215), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2214), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2213), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2212), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2211), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2210), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2209), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2208), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2207), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2206), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2205), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2204), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2203), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2202), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2201), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2200), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2199), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2198), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2197), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2196), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2195), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2194), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2193), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2192), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2191), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2190), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2189), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2188), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2187), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2186), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2185), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2184), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2183), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2182), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2181), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2180), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2179), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2178), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2177), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2176), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2175), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2174), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2173), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2172), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2171), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2170), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2169), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2168), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2167), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2166), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2165), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2164), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2163), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2162), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2161), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2160), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2159), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2158), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2157), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2156), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2155), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2154), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2153), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2152), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2151), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2150), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2149), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2148), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2147), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2146), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2145), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2144), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2143), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2142), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2141), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2140), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2139), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2138), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2137), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2136), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2135), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2134), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2133), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2132), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2131), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2130), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2129), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2128), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2127), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2126), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2125), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2124), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2123), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2122), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2121), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2120), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2119), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2118), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2117), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2116), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2115), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2114), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2113), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2112), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2111), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2110), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2109), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2108), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2107), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2106), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2105), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2104), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2103), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2102), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2101), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2100), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2099), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2098), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2097), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2096), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2095), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2094), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2093), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2092), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2091), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2090), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2089), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2088), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2087), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2086), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2085), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2084), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2083), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2082), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2081), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2080), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2079), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2078), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2077), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2076), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2075), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2074), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2073), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2072), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n2071), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n2070), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n2069), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n2068), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n2067), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n2066), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n2065), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n2064), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n2063), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n2062), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n2061), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n2060), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n2059), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n2058), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n2057), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n2056), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n2055), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n2054), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n2053), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n2052), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n2051), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n2050), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n2049), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n2048), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n2047), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n2046), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n2045), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n2044), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n2043), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n2042), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n2041), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n2040), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n2039), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n2038), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n2037), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n2036), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n2035), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n2034), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n2033), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n2032), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n2031), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n2030), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n2029), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n2028), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n2027), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n2026), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n2025), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n2024), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n2023), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n2022), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n2021), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n2020), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n2019), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n2018), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n2017), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n2016), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n2015), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n2014), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n2013), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n2012), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n2011), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n2010), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n2009), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n2008), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n2007), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n2006), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n2005), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n2004), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n2003), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n2002), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n2001), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n2000), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n1999), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n1998), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n1997), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n1996), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n1995), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n1994), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n1993), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n1992), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n1991), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n1990), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n1989), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n1988), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n1987), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n1986), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n1985), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n1984), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n1983), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n1982), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n1981), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n1980), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n1979), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n1978), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n1977), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n1976), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n1975), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n1974), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n1973), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n1972), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n1971), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n1970), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n1969), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n1968), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n1967), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n1966), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n1965), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n1964), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n1963), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n1962), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n1961), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n1960), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n1959), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n1958), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n1957), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n1956), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n1955), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n1954), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n1953), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n1952), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n1951), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n1950), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n1949), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n1948), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n1947), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n1946), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n1945), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n1944), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n1943), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n1942), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n1941), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n1940), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n1939), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n1938), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n1937), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n1936), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n1935), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n1934), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n1933), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n1932), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n1931), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n1930), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n1929), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n1928), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n1927), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n1926), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n1925), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n1924), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n1923), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n1922), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n1921), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n1920), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n1919), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n1918), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n1917), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n1916), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n1915), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n1914), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n1913), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n1912), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n1911), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n1910), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n1909), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n1908), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n1907), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n1906), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n1905), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n1904), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n1903), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n1902), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n1901), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n1900), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n1899), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n1898), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n1897), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n1896), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n1895), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n1894), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n1893), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n1892), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n1891), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n1890), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n1889), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n1888), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n1887), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n1886), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n1885), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n1884), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n1883), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n1882), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n1881), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n1880), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n1879), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n1878), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n1877), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n1876), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n1875), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n1874), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n1873), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n1872), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n1871), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n1870), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n1869), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n1868), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n1867), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n1866), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n1865), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n1864), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n1863), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n1862), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n1861), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n1860), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n1859), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n1858), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n1857), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n1856), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n1855), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n1854), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n1853), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n1852), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n1851), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n1850), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n1849), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n1848), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n1847), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n1846), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n1845), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n1844), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n1843), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n1842), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n1841), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n1840), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n1839), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n1838), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n1837), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n1836), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n1835), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n1834), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n1833), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n1832), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n1831), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n1830), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n1829), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n1828), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n1827), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n1826), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n1825), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n1824), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n1823), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n1822), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n1821), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n1820), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n1819), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n1818), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n1817), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n1816), .CLK(clk), .Q(\mem<63><0> ) );
  OAI21X1 U817 ( .A(n4555), .B(n5007), .C(n955), .Y(n1816) );
  OAI21X1 U819 ( .A(n4555), .B(n5006), .C(n954), .Y(n1817) );
  OAI21X1 U821 ( .A(n4555), .B(n5005), .C(n953), .Y(n1818) );
  OAI21X1 U823 ( .A(n4555), .B(n5004), .C(n952), .Y(n1819) );
  OAI21X1 U825 ( .A(n4555), .B(n5003), .C(n951), .Y(n1820) );
  OAI21X1 U827 ( .A(n4555), .B(n5002), .C(n950), .Y(n1821) );
  OAI21X1 U829 ( .A(n4555), .B(n5001), .C(n949), .Y(n1822) );
  OAI21X1 U831 ( .A(n4555), .B(n5000), .C(n948), .Y(n1823) );
  NAND3X1 U1905 ( .A(enable), .B(n1580), .C(wr), .Y(n625) );
  MUX2X1 U3 ( .B(\mem<31><5> ), .A(\mem<30><5> ), .S(n1489), .Y(n2813) );
  INVX8 U4 ( .A(n1549), .Y(n1) );
  INVX8 U5 ( .A(n1534), .Y(n1549) );
  INVX1 U6 ( .A(n588), .Y(n2) );
  OR2X2 U7 ( .A(n1610), .B(n1609), .Y(n485) );
  INVX4 U8 ( .A(n655), .Y(n790) );
  INVX4 U9 ( .A(n657), .Y(n791) );
  INVX4 U10 ( .A(n1465), .Y(n1466) );
  INVX1 U11 ( .A(n585), .Y(n3) );
  INVX1 U12 ( .A(n713), .Y(n4) );
  INVX1 U13 ( .A(n1424), .Y(n5) );
  BUFX4 U14 ( .A(n698), .Y(n6) );
  INVX1 U15 ( .A(n661), .Y(n7) );
  INVX1 U16 ( .A(n7), .Y(n8) );
  INVX1 U17 ( .A(n691), .Y(n9) );
  INVX1 U18 ( .A(n828), .Y(n10) );
  AND2X2 U19 ( .A(n91), .B(n400), .Y(n11) );
  AND2X2 U20 ( .A(n439), .B(n360), .Y(n12) );
  AND2X2 U21 ( .A(n513), .B(n1651), .Y(n13) );
  AND2X2 U22 ( .A(n712), .B(n515), .Y(n14) );
  INVX4 U23 ( .A(n645), .Y(n1517) );
  INVX8 U24 ( .A(n850), .Y(n851) );
  INVX2 U25 ( .A(n1455), .Y(n850) );
  AND2X2 U26 ( .A(n861), .B(n1515), .Y(n15) );
  INVX1 U27 ( .A(n642), .Y(n16) );
  AND2X2 U28 ( .A(n361), .B(n440), .Y(n17) );
  INVX1 U29 ( .A(n690), .Y(n1486) );
  AND2X2 U30 ( .A(n248), .B(n291), .Y(n414) );
  INVX1 U31 ( .A(n688), .Y(n18) );
  INVX1 U32 ( .A(n688), .Y(n19) );
  INVX2 U33 ( .A(n687), .Y(n688) );
  INVX1 U34 ( .A(n828), .Y(n20) );
  INVX1 U35 ( .A(n702), .Y(n21) );
  INVX1 U36 ( .A(n714), .Y(n22) );
  INVX1 U37 ( .A(n636), .Y(n23) );
  INVX1 U38 ( .A(n637), .Y(n24) );
  INVX1 U39 ( .A(n56), .Y(n25) );
  INVX1 U40 ( .A(n25), .Y(n26) );
  INVX4 U41 ( .A(n825), .Y(n849) );
  INVX4 U42 ( .A(n706), .Y(n833) );
  INVX8 U43 ( .A(n697), .Y(n3296) );
  INVX4 U44 ( .A(n696), .Y(n697) );
  INVX4 U45 ( .A(n598), .Y(n831) );
  INVX4 U46 ( .A(n633), .Y(n634) );
  INVX4 U47 ( .A(n601), .Y(n797) );
  AND2X2 U48 ( .A(n82), .B(n405), .Y(n27) );
  INVX1 U49 ( .A(n3029), .Y(n3007) );
  INVX1 U50 ( .A(n3082), .Y(n3060) );
  INVX1 U51 ( .A(n1527), .Y(n3168) );
  INVX1 U52 ( .A(n612), .Y(n1283) );
  INVX1 U53 ( .A(n3843), .Y(n3821) );
  INVX1 U54 ( .A(n3895), .Y(n3873) );
  OR2X1 U55 ( .A(n2379), .B(n2378), .Y(n185) );
  INVX1 U56 ( .A(n3002), .Y(n2979) );
  INVX1 U57 ( .A(n3055), .Y(n3033) );
  INVX1 U58 ( .A(n3109), .Y(n3086) );
  INVX1 U59 ( .A(n3137), .Y(n3115) );
  INVX1 U60 ( .A(n3265), .Y(n3243) );
  INVX1 U61 ( .A(n3292), .Y(n3270) );
  INVX1 U62 ( .A(n3319), .Y(n3297) );
  INVX1 U63 ( .A(n3347), .Y(n3325) );
  INVX1 U64 ( .A(n3789), .Y(n3767) );
  INVX1 U65 ( .A(n3817), .Y(n3794) );
  INVX1 U66 ( .A(n3869), .Y(n3847) );
  INVX1 U67 ( .A(n3922), .Y(n3900) );
  INVX1 U68 ( .A(n3949), .Y(n3927) );
  BUFX2 U69 ( .A(n3190), .Y(n1527) );
  OR2X1 U70 ( .A(n2374), .B(n2373), .Y(n499) );
  OR2X1 U71 ( .A(n2408), .B(n2407), .Y(n199) );
  INVX1 U72 ( .A(n1629), .Y(n1497) );
  INVX1 U73 ( .A(n2787), .Y(n2788) );
  OR2X1 U74 ( .A(n2329), .B(n2328), .Y(n497) );
  OR2X1 U75 ( .A(n1715), .B(n1714), .Y(n149) );
  OR2X1 U76 ( .A(n1770), .B(n1769), .Y(n495) );
  AND2X1 U77 ( .A(n4496), .B(n863), .Y(n1174) );
  AND2X1 U78 ( .A(n4496), .B(n865), .Y(n1176) );
  AND2X1 U79 ( .A(n4496), .B(n867), .Y(n1178) );
  AND2X1 U80 ( .A(n4496), .B(n869), .Y(n1180) );
  AND2X1 U81 ( .A(n4496), .B(n871), .Y(n1182) );
  AND2X1 U82 ( .A(n4496), .B(n873), .Y(n1184) );
  AND2X1 U83 ( .A(n4496), .B(n875), .Y(n1186) );
  AND2X1 U84 ( .A(n4496), .B(n877), .Y(n1188) );
  AND2X1 U85 ( .A(n4496), .B(n879), .Y(n1190) );
  AND2X1 U86 ( .A(n4496), .B(n881), .Y(n1192) );
  AND2X1 U87 ( .A(n4496), .B(n883), .Y(n1194) );
  AND2X1 U88 ( .A(n4496), .B(n885), .Y(n1196) );
  AND2X1 U89 ( .A(n1528), .B(n887), .Y(n1198) );
  AND2X1 U90 ( .A(n1528), .B(n889), .Y(n1200) );
  AND2X1 U91 ( .A(n1528), .B(n891), .Y(n1202) );
  AND2X1 U92 ( .A(n1528), .B(n895), .Y(n1206) );
  AND2X1 U93 ( .A(n1528), .B(n899), .Y(n1210) );
  AND2X1 U94 ( .A(n1528), .B(n901), .Y(n1212) );
  AND2X1 U95 ( .A(n1528), .B(n903), .Y(n1214) );
  AND2X1 U96 ( .A(n1528), .B(n905), .Y(n1216) );
  AND2X1 U97 ( .A(n1528), .B(n907), .Y(n1218) );
  AND2X1 U98 ( .A(n1529), .B(n909), .Y(n1220) );
  AND2X1 U99 ( .A(n1529), .B(n911), .Y(n1222) );
  AND2X1 U100 ( .A(n1529), .B(n913), .Y(n1224) );
  AND2X1 U101 ( .A(n1529), .B(n915), .Y(n1226) );
  AND2X1 U102 ( .A(n1529), .B(n919), .Y(n1230) );
  AND2X1 U103 ( .A(n1529), .B(n921), .Y(n1232) );
  AND2X1 U104 ( .A(n1529), .B(n923), .Y(n1234) );
  AND2X1 U105 ( .A(n1529), .B(n925), .Y(n1236) );
  AND2X1 U106 ( .A(n1275), .B(n693), .Y(n924) );
  AND2X1 U107 ( .A(n1530), .B(n927), .Y(n1238) );
  AND2X1 U108 ( .A(n4272), .B(n693), .Y(n926) );
  AND2X1 U109 ( .A(n1530), .B(n929), .Y(n1240) );
  AND2X1 U110 ( .A(n1529), .B(n931), .Y(n1242) );
  AND2X1 U111 ( .A(n1530), .B(n935), .Y(n1246) );
  AND2X1 U112 ( .A(n1530), .B(n937), .Y(n1248) );
  AND2X1 U113 ( .A(n1530), .B(n941), .Y(n1252) );
  AND2X1 U114 ( .A(n1530), .B(n943), .Y(n1254) );
  AND2X1 U115 ( .A(n1530), .B(n945), .Y(n1256) );
  AND2X1 U116 ( .A(n1281), .B(n2976), .Y(n4555) );
  INVX1 U117 ( .A(\mem<61><0> ), .Y(n4999) );
  INVX1 U118 ( .A(\mem<61><1> ), .Y(n4998) );
  INVX1 U119 ( .A(\mem<61><2> ), .Y(n4997) );
  INVX1 U120 ( .A(\mem<61><3> ), .Y(n4996) );
  INVX1 U121 ( .A(\mem<61><4> ), .Y(n4995) );
  INVX1 U122 ( .A(\mem<61><5> ), .Y(n4994) );
  INVX1 U123 ( .A(\mem<61><6> ), .Y(n4993) );
  INVX1 U124 ( .A(\mem<61><7> ), .Y(n4992) );
  AND2X1 U125 ( .A(n827), .B(n3007), .Y(n1292) );
  INVX1 U126 ( .A(\mem<59><0> ), .Y(n4991) );
  INVX1 U127 ( .A(\mem<59><1> ), .Y(n4990) );
  INVX1 U128 ( .A(\mem<59><2> ), .Y(n4989) );
  INVX1 U129 ( .A(\mem<59><3> ), .Y(n4988) );
  INVX1 U130 ( .A(\mem<59><4> ), .Y(n4987) );
  INVX1 U131 ( .A(\mem<59><5> ), .Y(n4986) );
  INVX1 U132 ( .A(\mem<59><6> ), .Y(n4985) );
  INVX1 U133 ( .A(\mem<59><7> ), .Y(n4984) );
  AND2X1 U134 ( .A(n794), .B(n3060), .Y(n1296) );
  INVX1 U135 ( .A(\mem<56><0> ), .Y(n4983) );
  INVX1 U136 ( .A(\mem<56><1> ), .Y(n4982) );
  INVX1 U137 ( .A(\mem<56><2> ), .Y(n4981) );
  INVX1 U138 ( .A(\mem<56><3> ), .Y(n4980) );
  INVX1 U139 ( .A(\mem<56><4> ), .Y(n4979) );
  INVX1 U140 ( .A(\mem<56><5> ), .Y(n4978) );
  INVX1 U141 ( .A(\mem<56><6> ), .Y(n4977) );
  INVX1 U142 ( .A(\mem<56><7> ), .Y(n4976) );
  INVX1 U143 ( .A(\mem<55><0> ), .Y(n4975) );
  INVX1 U144 ( .A(\mem<55><1> ), .Y(n4974) );
  INVX1 U145 ( .A(\mem<55><2> ), .Y(n4973) );
  INVX1 U146 ( .A(\mem<55><3> ), .Y(n4972) );
  INVX1 U147 ( .A(\mem<55><4> ), .Y(n4971) );
  INVX1 U148 ( .A(\mem<55><5> ), .Y(n4970) );
  INVX1 U149 ( .A(\mem<55><6> ), .Y(n4969) );
  INVX1 U150 ( .A(\mem<55><7> ), .Y(n4968) );
  AND2X1 U151 ( .A(n831), .B(n3168), .Y(n1304) );
  INVX1 U152 ( .A(\mem<54><0> ), .Y(n4967) );
  INVX1 U153 ( .A(\mem<54><1> ), .Y(n4966) );
  INVX1 U154 ( .A(\mem<54><2> ), .Y(n4965) );
  INVX1 U155 ( .A(\mem<54><3> ), .Y(n4964) );
  INVX1 U156 ( .A(\mem<54><4> ), .Y(n4963) );
  INVX1 U157 ( .A(\mem<54><5> ), .Y(n4962) );
  INVX1 U158 ( .A(\mem<54><6> ), .Y(n4961) );
  INVX1 U159 ( .A(\mem<54><7> ), .Y(n4960) );
  INVX1 U160 ( .A(\mem<53><0> ), .Y(n4959) );
  INVX1 U161 ( .A(\mem<53><1> ), .Y(n4958) );
  INVX1 U162 ( .A(\mem<53><2> ), .Y(n4957) );
  INVX1 U163 ( .A(\mem<53><3> ), .Y(n4956) );
  INVX1 U164 ( .A(\mem<53><4> ), .Y(n4955) );
  INVX1 U165 ( .A(\mem<53><5> ), .Y(n4954) );
  INVX1 U166 ( .A(\mem<53><6> ), .Y(n4953) );
  INVX1 U167 ( .A(\mem<53><7> ), .Y(n4952) );
  INVX1 U168 ( .A(\mem<52><0> ), .Y(n4951) );
  INVX1 U169 ( .A(\mem<52><1> ), .Y(n4950) );
  INVX1 U170 ( .A(\mem<52><2> ), .Y(n4949) );
  INVX1 U171 ( .A(\mem<52><3> ), .Y(n4948) );
  INVX1 U172 ( .A(\mem<52><4> ), .Y(n4947) );
  INVX1 U173 ( .A(\mem<52><5> ), .Y(n4946) );
  INVX1 U174 ( .A(\mem<52><6> ), .Y(n4945) );
  INVX1 U175 ( .A(\mem<52><7> ), .Y(n4944) );
  INVX1 U176 ( .A(\mem<51><0> ), .Y(n4943) );
  INVX1 U177 ( .A(\mem<51><1> ), .Y(n4942) );
  INVX1 U178 ( .A(\mem<51><2> ), .Y(n4941) );
  INVX1 U179 ( .A(\mem<51><3> ), .Y(n4940) );
  INVX1 U180 ( .A(\mem<51><4> ), .Y(n4939) );
  INVX1 U181 ( .A(\mem<51><5> ), .Y(n4938) );
  INVX1 U182 ( .A(\mem<51><6> ), .Y(n4937) );
  INVX1 U183 ( .A(\mem<51><7> ), .Y(n4936) );
  INVX1 U184 ( .A(\mem<50><0> ), .Y(n4935) );
  INVX1 U185 ( .A(\mem<50><1> ), .Y(n4934) );
  INVX1 U186 ( .A(\mem<50><2> ), .Y(n4933) );
  INVX1 U187 ( .A(\mem<50><3> ), .Y(n4932) );
  INVX1 U188 ( .A(\mem<50><4> ), .Y(n4931) );
  INVX1 U189 ( .A(\mem<50><5> ), .Y(n4930) );
  INVX1 U190 ( .A(\mem<50><6> ), .Y(n4929) );
  INVX1 U191 ( .A(\mem<50><7> ), .Y(n4928) );
  INVX1 U192 ( .A(\mem<49><0> ), .Y(n4927) );
  INVX1 U193 ( .A(\mem<49><1> ), .Y(n4926) );
  INVX1 U194 ( .A(\mem<49><2> ), .Y(n4925) );
  INVX1 U195 ( .A(\mem<49><3> ), .Y(n4924) );
  INVX1 U196 ( .A(\mem<49><4> ), .Y(n4923) );
  INVX1 U197 ( .A(\mem<49><5> ), .Y(n4922) );
  INVX1 U198 ( .A(\mem<49><6> ), .Y(n4921) );
  INVX1 U199 ( .A(\mem<49><7> ), .Y(n4920) );
  INVX1 U200 ( .A(\mem<48><0> ), .Y(n4919) );
  INVX1 U201 ( .A(\mem<48><1> ), .Y(n4918) );
  INVX1 U202 ( .A(\mem<48><2> ), .Y(n4917) );
  INVX1 U203 ( .A(\mem<48><3> ), .Y(n4916) );
  INVX1 U204 ( .A(\mem<48><4> ), .Y(n4915) );
  INVX1 U205 ( .A(\mem<48><5> ), .Y(n4914) );
  INVX1 U206 ( .A(\mem<48><6> ), .Y(n4913) );
  INVX1 U207 ( .A(\mem<48><7> ), .Y(n4912) );
  INVX1 U208 ( .A(\mem<47><0> ), .Y(n4911) );
  INVX1 U209 ( .A(\mem<47><1> ), .Y(n4910) );
  INVX1 U210 ( .A(\mem<47><2> ), .Y(n4909) );
  INVX1 U211 ( .A(\mem<47><3> ), .Y(n4908) );
  INVX1 U212 ( .A(\mem<47><4> ), .Y(n4907) );
  INVX1 U213 ( .A(\mem<47><5> ), .Y(n4906) );
  INVX1 U214 ( .A(\mem<47><6> ), .Y(n4905) );
  INVX1 U215 ( .A(\mem<47><7> ), .Y(n4904) );
  INVX1 U216 ( .A(\mem<46><0> ), .Y(n4903) );
  INVX1 U217 ( .A(\mem<46><1> ), .Y(n4902) );
  INVX1 U218 ( .A(\mem<46><2> ), .Y(n4901) );
  INVX1 U219 ( .A(\mem<46><3> ), .Y(n4900) );
  INVX1 U220 ( .A(\mem<46><4> ), .Y(n4899) );
  INVX1 U221 ( .A(\mem<46><5> ), .Y(n4898) );
  INVX1 U222 ( .A(\mem<46><6> ), .Y(n4897) );
  INVX1 U223 ( .A(\mem<46><7> ), .Y(n4896) );
  INVX1 U224 ( .A(\mem<45><0> ), .Y(n4895) );
  INVX1 U225 ( .A(\mem<45><1> ), .Y(n4894) );
  INVX1 U226 ( .A(\mem<45><2> ), .Y(n4893) );
  INVX1 U227 ( .A(\mem<45><3> ), .Y(n4892) );
  INVX1 U228 ( .A(\mem<45><4> ), .Y(n4891) );
  INVX1 U229 ( .A(\mem<45><5> ), .Y(n4890) );
  INVX1 U230 ( .A(\mem<45><6> ), .Y(n4889) );
  INVX1 U231 ( .A(\mem<45><7> ), .Y(n4888) );
  INVX1 U232 ( .A(\mem<44><0> ), .Y(n4887) );
  INVX1 U233 ( .A(\mem<44><1> ), .Y(n4886) );
  INVX1 U234 ( .A(\mem<44><2> ), .Y(n4885) );
  INVX1 U235 ( .A(\mem<44><3> ), .Y(n4884) );
  INVX1 U236 ( .A(\mem<44><4> ), .Y(n4883) );
  INVX1 U237 ( .A(\mem<44><5> ), .Y(n4882) );
  INVX1 U238 ( .A(\mem<44><6> ), .Y(n4881) );
  INVX1 U239 ( .A(\mem<44><7> ), .Y(n4880) );
  INVX1 U240 ( .A(\mem<43><0> ), .Y(n4879) );
  INVX1 U241 ( .A(\mem<43><1> ), .Y(n4878) );
  INVX1 U242 ( .A(\mem<43><2> ), .Y(n4877) );
  INVX1 U243 ( .A(\mem<43><3> ), .Y(n4876) );
  INVX1 U244 ( .A(\mem<43><4> ), .Y(n4875) );
  INVX1 U245 ( .A(\mem<43><5> ), .Y(n4874) );
  INVX1 U246 ( .A(\mem<43><6> ), .Y(n4873) );
  INVX1 U247 ( .A(\mem<43><7> ), .Y(n4872) );
  INVX1 U248 ( .A(\mem<42><0> ), .Y(n4871) );
  INVX1 U249 ( .A(\mem<42><1> ), .Y(n4870) );
  INVX1 U250 ( .A(\mem<42><2> ), .Y(n4869) );
  INVX1 U251 ( .A(\mem<42><3> ), .Y(n4868) );
  INVX1 U252 ( .A(\mem<42><4> ), .Y(n4867) );
  INVX1 U253 ( .A(\mem<42><5> ), .Y(n4866) );
  INVX1 U254 ( .A(\mem<42><6> ), .Y(n4865) );
  INVX1 U255 ( .A(\mem<42><7> ), .Y(n4864) );
  INVX1 U256 ( .A(\mem<41><1> ), .Y(n4862) );
  INVX1 U257 ( .A(\mem<41><2> ), .Y(n4861) );
  INVX1 U258 ( .A(\mem<41><3> ), .Y(n4860) );
  INVX1 U259 ( .A(\mem<41><4> ), .Y(n4859) );
  INVX1 U260 ( .A(\mem<41><5> ), .Y(n4858) );
  INVX1 U261 ( .A(\mem<41><6> ), .Y(n4857) );
  INVX1 U262 ( .A(\mem<41><7> ), .Y(n4856) );
  INVX1 U263 ( .A(\mem<40><0> ), .Y(n4855) );
  INVX1 U264 ( .A(\mem<40><1> ), .Y(n4854) );
  INVX1 U265 ( .A(\mem<40><2> ), .Y(n4853) );
  INVX1 U266 ( .A(\mem<40><3> ), .Y(n4852) );
  INVX1 U267 ( .A(\mem<40><4> ), .Y(n4851) );
  INVX1 U268 ( .A(\mem<40><5> ), .Y(n4850) );
  INVX1 U269 ( .A(\mem<40><6> ), .Y(n4849) );
  INVX1 U270 ( .A(\mem<40><7> ), .Y(n4848) );
  INVX1 U271 ( .A(\mem<39><0> ), .Y(n4847) );
  INVX1 U272 ( .A(\mem<39><1> ), .Y(n4846) );
  INVX1 U273 ( .A(\mem<39><2> ), .Y(n4845) );
  INVX1 U274 ( .A(\mem<39><3> ), .Y(n4844) );
  INVX1 U275 ( .A(\mem<39><4> ), .Y(n4843) );
  INVX1 U276 ( .A(\mem<39><5> ), .Y(n4842) );
  INVX1 U277 ( .A(\mem<39><6> ), .Y(n4841) );
  INVX1 U278 ( .A(\mem<39><7> ), .Y(n4840) );
  INVX1 U279 ( .A(\mem<38><0> ), .Y(n4839) );
  INVX1 U280 ( .A(\mem<38><1> ), .Y(n4838) );
  INVX1 U281 ( .A(\mem<38><2> ), .Y(n4837) );
  INVX1 U282 ( .A(\mem<38><3> ), .Y(n4836) );
  INVX1 U283 ( .A(\mem<38><4> ), .Y(n4835) );
  INVX1 U284 ( .A(\mem<38><5> ), .Y(n4834) );
  INVX1 U285 ( .A(\mem<38><6> ), .Y(n4833) );
  INVX1 U286 ( .A(\mem<38><7> ), .Y(n4832) );
  INVX1 U287 ( .A(\mem<37><0> ), .Y(n4831) );
  INVX1 U288 ( .A(\mem<37><1> ), .Y(n4830) );
  INVX1 U289 ( .A(\mem<37><2> ), .Y(n4829) );
  INVX1 U290 ( .A(\mem<37><3> ), .Y(n4828) );
  INVX1 U291 ( .A(\mem<37><4> ), .Y(n4827) );
  INVX1 U292 ( .A(\mem<37><5> ), .Y(n4826) );
  INVX1 U293 ( .A(\mem<37><6> ), .Y(n4825) );
  INVX1 U294 ( .A(\mem<37><7> ), .Y(n4824) );
  INVX1 U295 ( .A(\mem<36><0> ), .Y(n4823) );
  INVX1 U296 ( .A(\mem<36><1> ), .Y(n4822) );
  INVX1 U297 ( .A(\mem<36><2> ), .Y(n4821) );
  INVX1 U298 ( .A(\mem<36><3> ), .Y(n4820) );
  INVX1 U299 ( .A(\mem<36><4> ), .Y(n4819) );
  INVX1 U300 ( .A(\mem<36><5> ), .Y(n4818) );
  INVX1 U301 ( .A(\mem<36><6> ), .Y(n4817) );
  INVX1 U302 ( .A(\mem<36><7> ), .Y(n4816) );
  INVX1 U303 ( .A(\mem<35><0> ), .Y(n4815) );
  INVX1 U304 ( .A(\mem<35><1> ), .Y(n4814) );
  INVX1 U305 ( .A(\mem<35><2> ), .Y(n4813) );
  INVX1 U306 ( .A(\mem<35><3> ), .Y(n4812) );
  INVX1 U307 ( .A(\mem<35><4> ), .Y(n4811) );
  INVX1 U308 ( .A(\mem<35><5> ), .Y(n4810) );
  INVX1 U309 ( .A(\mem<35><6> ), .Y(n4809) );
  INVX1 U310 ( .A(\mem<35><7> ), .Y(n4808) );
  INVX1 U311 ( .A(\mem<34><0> ), .Y(n4807) );
  INVX1 U312 ( .A(\mem<34><1> ), .Y(n4806) );
  INVX1 U313 ( .A(\mem<34><2> ), .Y(n4805) );
  INVX1 U314 ( .A(\mem<34><3> ), .Y(n4804) );
  INVX1 U315 ( .A(\mem<34><4> ), .Y(n4803) );
  INVX1 U316 ( .A(\mem<34><5> ), .Y(n4802) );
  INVX1 U317 ( .A(\mem<34><6> ), .Y(n4801) );
  INVX1 U318 ( .A(\mem<34><7> ), .Y(n4800) );
  INVX1 U319 ( .A(\mem<33><0> ), .Y(n4799) );
  INVX1 U320 ( .A(\mem<33><1> ), .Y(n4798) );
  INVX1 U321 ( .A(\mem<33><2> ), .Y(n4797) );
  INVX1 U322 ( .A(\mem<33><3> ), .Y(n4796) );
  INVX1 U323 ( .A(\mem<33><4> ), .Y(n4795) );
  INVX1 U324 ( .A(\mem<33><5> ), .Y(n4794) );
  INVX1 U325 ( .A(\mem<33><6> ), .Y(n4793) );
  INVX1 U326 ( .A(\mem<33><7> ), .Y(n4792) );
  INVX1 U327 ( .A(\mem<32><0> ), .Y(n4791) );
  INVX1 U328 ( .A(\mem<32><1> ), .Y(n4790) );
  INVX1 U329 ( .A(\mem<32><2> ), .Y(n4789) );
  INVX1 U330 ( .A(\mem<32><3> ), .Y(n4788) );
  INVX1 U331 ( .A(\mem<32><4> ), .Y(n4787) );
  INVX1 U332 ( .A(\mem<32><5> ), .Y(n4786) );
  INVX1 U333 ( .A(\mem<32><6> ), .Y(n4785) );
  INVX1 U334 ( .A(\mem<32><7> ), .Y(n4784) );
  INVX1 U335 ( .A(\mem<31><2> ), .Y(n4782) );
  INVX1 U336 ( .A(\mem<31><3> ), .Y(n4781) );
  INVX1 U337 ( .A(\mem<31><4> ), .Y(n4780) );
  INVX1 U338 ( .A(\mem<31><5> ), .Y(n4779) );
  INVX1 U339 ( .A(\mem<31><6> ), .Y(n4778) );
  INVX1 U340 ( .A(\mem<31><7> ), .Y(n4777) );
  INVX1 U341 ( .A(\mem<30><0> ), .Y(n4776) );
  INVX1 U342 ( .A(\mem<30><1> ), .Y(n4775) );
  INVX1 U343 ( .A(\mem<29><2> ), .Y(n4773) );
  INVX1 U344 ( .A(\mem<29><3> ), .Y(n4772) );
  INVX1 U345 ( .A(\mem<29><4> ), .Y(n4771) );
  INVX1 U346 ( .A(\mem<29><5> ), .Y(n4770) );
  INVX1 U347 ( .A(\mem<29><6> ), .Y(n4769) );
  INVX1 U348 ( .A(\mem<29><7> ), .Y(n4768) );
  AND2X1 U349 ( .A(n804), .B(n3821), .Y(n1356) );
  INVX1 U350 ( .A(\mem<28><0> ), .Y(n4767) );
  INVX1 U351 ( .A(\mem<28><1> ), .Y(n4766) );
  INVX1 U352 ( .A(\mem<27><2> ), .Y(n4765) );
  INVX1 U353 ( .A(\mem<27><3> ), .Y(n4764) );
  INVX1 U354 ( .A(\mem<27><4> ), .Y(n4763) );
  INVX1 U355 ( .A(\mem<27><5> ), .Y(n4762) );
  INVX1 U356 ( .A(\mem<27><6> ), .Y(n4761) );
  INVX1 U357 ( .A(\mem<27><7> ), .Y(n4760) );
  AND2X1 U358 ( .A(n836), .B(n3873), .Y(n1360) );
  INVX1 U359 ( .A(\mem<26><0> ), .Y(n4759) );
  INVX1 U360 ( .A(\mem<26><1> ), .Y(n4758) );
  INVX1 U361 ( .A(\mem<24><0> ), .Y(n4757) );
  INVX1 U362 ( .A(\mem<24><1> ), .Y(n4756) );
  INVX1 U363 ( .A(\mem<24><2> ), .Y(n4755) );
  INVX1 U364 ( .A(\mem<24><3> ), .Y(n4754) );
  INVX1 U365 ( .A(\mem<24><4> ), .Y(n4753) );
  INVX1 U366 ( .A(\mem<24><5> ), .Y(n4752) );
  INVX1 U367 ( .A(\mem<24><6> ), .Y(n4751) );
  INVX1 U368 ( .A(\mem<24><7> ), .Y(n4750) );
  INVX1 U369 ( .A(\mem<23><0> ), .Y(n4749) );
  INVX1 U370 ( .A(\mem<23><1> ), .Y(n4748) );
  INVX1 U371 ( .A(\mem<23><2> ), .Y(n4747) );
  INVX1 U372 ( .A(\mem<23><3> ), .Y(n4746) );
  INVX1 U373 ( .A(\mem<23><4> ), .Y(n4745) );
  INVX1 U374 ( .A(\mem<23><5> ), .Y(n4744) );
  INVX1 U375 ( .A(\mem<23><6> ), .Y(n4743) );
  INVX1 U376 ( .A(\mem<23><7> ), .Y(n4742) );
  INVX1 U377 ( .A(\mem<22><0> ), .Y(n4741) );
  INVX1 U378 ( .A(\mem<22><1> ), .Y(n4740) );
  INVX1 U379 ( .A(\mem<22><2> ), .Y(n4739) );
  INVX1 U380 ( .A(\mem<22><3> ), .Y(n4738) );
  INVX1 U381 ( .A(\mem<22><4> ), .Y(n4737) );
  INVX1 U382 ( .A(\mem<22><5> ), .Y(n4736) );
  INVX1 U383 ( .A(\mem<22><6> ), .Y(n4735) );
  INVX1 U384 ( .A(\mem<22><7> ), .Y(n4734) );
  INVX1 U385 ( .A(\mem<21><0> ), .Y(n4733) );
  INVX1 U386 ( .A(\mem<21><1> ), .Y(n4732) );
  INVX1 U387 ( .A(\mem<21><2> ), .Y(n4731) );
  INVX1 U388 ( .A(\mem<21><3> ), .Y(n4730) );
  INVX1 U389 ( .A(\mem<21><4> ), .Y(n4729) );
  INVX1 U390 ( .A(\mem<21><5> ), .Y(n4728) );
  INVX1 U391 ( .A(\mem<21><6> ), .Y(n4727) );
  INVX1 U392 ( .A(\mem<21><7> ), .Y(n4726) );
  INVX1 U393 ( .A(\mem<20><0> ), .Y(n4725) );
  INVX1 U394 ( .A(\mem<20><1> ), .Y(n4724) );
  INVX1 U395 ( .A(\mem<20><2> ), .Y(n4723) );
  INVX1 U396 ( .A(\mem<20><3> ), .Y(n4722) );
  INVX1 U397 ( .A(\mem<20><4> ), .Y(n4721) );
  INVX1 U398 ( .A(\mem<20><5> ), .Y(n4720) );
  INVX1 U399 ( .A(\mem<20><6> ), .Y(n4719) );
  INVX1 U400 ( .A(\mem<20><7> ), .Y(n4718) );
  INVX1 U401 ( .A(\mem<19><0> ), .Y(n4717) );
  INVX1 U402 ( .A(\mem<19><1> ), .Y(n4716) );
  INVX1 U403 ( .A(\mem<19><2> ), .Y(n4715) );
  INVX1 U404 ( .A(\mem<19><3> ), .Y(n4714) );
  INVX1 U405 ( .A(\mem<19><4> ), .Y(n4713) );
  INVX1 U406 ( .A(\mem<19><5> ), .Y(n4712) );
  INVX1 U407 ( .A(\mem<19><6> ), .Y(n4711) );
  INVX1 U408 ( .A(\mem<19><7> ), .Y(n4710) );
  INVX1 U409 ( .A(\mem<18><0> ), .Y(n4709) );
  INVX1 U410 ( .A(\mem<18><1> ), .Y(n4708) );
  INVX1 U411 ( .A(\mem<18><2> ), .Y(n4707) );
  INVX1 U412 ( .A(\mem<18><3> ), .Y(n4706) );
  INVX1 U413 ( .A(\mem<18><4> ), .Y(n4705) );
  INVX1 U414 ( .A(\mem<18><5> ), .Y(n4704) );
  INVX1 U415 ( .A(\mem<18><6> ), .Y(n4703) );
  INVX1 U416 ( .A(\mem<18><7> ), .Y(n4702) );
  INVX1 U417 ( .A(\mem<17><0> ), .Y(n4701) );
  INVX1 U418 ( .A(\mem<17><1> ), .Y(n4700) );
  INVX1 U419 ( .A(\mem<17><2> ), .Y(n4699) );
  INVX1 U420 ( .A(\mem<17><3> ), .Y(n4698) );
  INVX1 U421 ( .A(\mem<17><4> ), .Y(n4697) );
  INVX1 U422 ( .A(\mem<17><5> ), .Y(n4696) );
  INVX1 U423 ( .A(\mem<17><6> ), .Y(n4695) );
  INVX1 U424 ( .A(\mem<17><7> ), .Y(n4694) );
  INVX1 U425 ( .A(\mem<16><0> ), .Y(n4693) );
  INVX1 U426 ( .A(\mem<16><1> ), .Y(n4692) );
  INVX1 U427 ( .A(\mem<16><2> ), .Y(n4691) );
  INVX1 U428 ( .A(\mem<16><3> ), .Y(n4690) );
  INVX1 U429 ( .A(\mem<16><4> ), .Y(n4689) );
  INVX1 U430 ( .A(\mem<16><5> ), .Y(n4688) );
  INVX1 U431 ( .A(\mem<16><6> ), .Y(n4687) );
  INVX1 U432 ( .A(\mem<16><7> ), .Y(n4686) );
  INVX1 U433 ( .A(\mem<15><0> ), .Y(n4685) );
  INVX1 U434 ( .A(\mem<15><1> ), .Y(n4684) );
  INVX1 U435 ( .A(\mem<15><2> ), .Y(n4683) );
  INVX1 U436 ( .A(\mem<15><3> ), .Y(n4682) );
  INVX1 U437 ( .A(\mem<15><4> ), .Y(n4681) );
  INVX1 U438 ( .A(\mem<15><5> ), .Y(n4680) );
  INVX1 U439 ( .A(\mem<15><6> ), .Y(n4679) );
  INVX1 U440 ( .A(\mem<15><7> ), .Y(n4678) );
  INVX1 U441 ( .A(\mem<14><0> ), .Y(n4677) );
  INVX1 U442 ( .A(\mem<14><1> ), .Y(n4676) );
  INVX1 U443 ( .A(\mem<14><2> ), .Y(n4675) );
  INVX1 U444 ( .A(\mem<14><3> ), .Y(n4674) );
  INVX1 U445 ( .A(\mem<14><4> ), .Y(n4673) );
  INVX1 U446 ( .A(\mem<14><5> ), .Y(n4672) );
  INVX1 U447 ( .A(\mem<14><6> ), .Y(n4671) );
  INVX1 U448 ( .A(\mem<14><7> ), .Y(n4670) );
  INVX1 U449 ( .A(\mem<13><0> ), .Y(n4669) );
  INVX1 U450 ( .A(\mem<13><1> ), .Y(n4668) );
  INVX1 U451 ( .A(\mem<13><2> ), .Y(n4667) );
  INVX1 U452 ( .A(\mem<13><3> ), .Y(n4666) );
  INVX1 U453 ( .A(\mem<13><4> ), .Y(n4665) );
  INVX1 U454 ( .A(\mem<13><5> ), .Y(n4664) );
  INVX1 U455 ( .A(\mem<13><6> ), .Y(n4663) );
  INVX1 U456 ( .A(\mem<13><7> ), .Y(n4662) );
  INVX1 U457 ( .A(\mem<12><0> ), .Y(n4661) );
  INVX1 U458 ( .A(\mem<12><1> ), .Y(n4660) );
  INVX1 U459 ( .A(\mem<12><2> ), .Y(n4659) );
  INVX1 U460 ( .A(\mem<12><3> ), .Y(n4658) );
  INVX1 U461 ( .A(\mem<12><4> ), .Y(n4657) );
  INVX1 U462 ( .A(\mem<12><5> ), .Y(n4656) );
  INVX1 U463 ( .A(\mem<12><6> ), .Y(n4655) );
  INVX1 U464 ( .A(\mem<12><7> ), .Y(n4654) );
  INVX1 U465 ( .A(\mem<11><0> ), .Y(n4653) );
  INVX1 U466 ( .A(\mem<11><1> ), .Y(n4652) );
  INVX1 U467 ( .A(\mem<11><2> ), .Y(n4651) );
  INVX1 U468 ( .A(\mem<11><3> ), .Y(n4650) );
  INVX1 U469 ( .A(\mem<11><4> ), .Y(n4649) );
  INVX1 U470 ( .A(\mem<11><5> ), .Y(n4648) );
  INVX1 U471 ( .A(\mem<11><6> ), .Y(n4647) );
  INVX1 U472 ( .A(\mem<11><7> ), .Y(n4646) );
  INVX1 U473 ( .A(\mem<10><0> ), .Y(n4645) );
  INVX1 U474 ( .A(\mem<10><1> ), .Y(n4644) );
  INVX1 U475 ( .A(\mem<10><2> ), .Y(n4643) );
  INVX1 U476 ( .A(\mem<10><3> ), .Y(n4642) );
  INVX1 U477 ( .A(\mem<10><4> ), .Y(n4641) );
  INVX1 U478 ( .A(\mem<10><5> ), .Y(n4640) );
  INVX1 U479 ( .A(\mem<10><6> ), .Y(n4639) );
  INVX1 U480 ( .A(\mem<10><7> ), .Y(n4638) );
  INVX1 U481 ( .A(\mem<9><0> ), .Y(n4637) );
  INVX1 U482 ( .A(\mem<9><1> ), .Y(n4636) );
  INVX1 U483 ( .A(\mem<9><2> ), .Y(n4635) );
  INVX1 U484 ( .A(\mem<9><3> ), .Y(n4634) );
  INVX1 U485 ( .A(\mem<9><4> ), .Y(n4633) );
  INVX1 U486 ( .A(\mem<9><5> ), .Y(n4632) );
  INVX1 U487 ( .A(\mem<9><6> ), .Y(n4631) );
  INVX1 U488 ( .A(\mem<9><7> ), .Y(n4630) );
  INVX1 U489 ( .A(\mem<8><0> ), .Y(n4629) );
  INVX1 U490 ( .A(\mem<8><1> ), .Y(n4628) );
  INVX1 U491 ( .A(\mem<8><2> ), .Y(n4627) );
  INVX1 U492 ( .A(\mem<8><3> ), .Y(n4626) );
  INVX1 U493 ( .A(\mem<8><4> ), .Y(n4625) );
  INVX1 U494 ( .A(\mem<8><5> ), .Y(n4624) );
  INVX1 U495 ( .A(\mem<8><6> ), .Y(n4623) );
  INVX1 U496 ( .A(\mem<8><7> ), .Y(n4622) );
  INVX1 U497 ( .A(\mem<7><0> ), .Y(n4621) );
  INVX1 U498 ( .A(\mem<7><1> ), .Y(n4620) );
  INVX1 U499 ( .A(\mem<7><2> ), .Y(n4619) );
  INVX1 U500 ( .A(\mem<7><3> ), .Y(n4618) );
  INVX1 U501 ( .A(\mem<7><4> ), .Y(n4617) );
  INVX1 U502 ( .A(\mem<7><5> ), .Y(n4616) );
  INVX1 U503 ( .A(\mem<7><6> ), .Y(n4615) );
  INVX1 U504 ( .A(\mem<7><7> ), .Y(n4614) );
  INVX1 U505 ( .A(\mem<6><0> ), .Y(n4613) );
  INVX1 U506 ( .A(\mem<6><1> ), .Y(n4612) );
  INVX1 U507 ( .A(\mem<6><2> ), .Y(n4611) );
  INVX1 U508 ( .A(\mem<6><3> ), .Y(n4610) );
  INVX1 U509 ( .A(\mem<6><4> ), .Y(n4609) );
  INVX1 U510 ( .A(\mem<6><5> ), .Y(n4608) );
  INVX1 U511 ( .A(\mem<6><6> ), .Y(n4607) );
  INVX1 U512 ( .A(\mem<6><7> ), .Y(n4606) );
  INVX1 U513 ( .A(\mem<5><0> ), .Y(n4605) );
  INVX1 U514 ( .A(\mem<5><1> ), .Y(n4604) );
  INVX1 U515 ( .A(\mem<5><2> ), .Y(n4603) );
  INVX1 U516 ( .A(\mem<5><3> ), .Y(n4602) );
  INVX1 U517 ( .A(\mem<5><4> ), .Y(n4601) );
  INVX1 U518 ( .A(\mem<5><5> ), .Y(n4600) );
  INVX1 U519 ( .A(\mem<5><6> ), .Y(n4599) );
  INVX1 U520 ( .A(\mem<5><7> ), .Y(n4598) );
  INVX1 U521 ( .A(\mem<4><0> ), .Y(n4597) );
  INVX1 U522 ( .A(\mem<4><1> ), .Y(n4596) );
  INVX1 U523 ( .A(\mem<4><2> ), .Y(n4595) );
  INVX1 U524 ( .A(\mem<4><3> ), .Y(n4594) );
  INVX1 U525 ( .A(\mem<4><4> ), .Y(n4593) );
  INVX1 U526 ( .A(\mem<4><5> ), .Y(n4592) );
  INVX1 U527 ( .A(\mem<4><6> ), .Y(n4591) );
  INVX1 U528 ( .A(\mem<4><7> ), .Y(n4590) );
  INVX1 U529 ( .A(\mem<3><0> ), .Y(n4589) );
  INVX1 U530 ( .A(\mem<3><1> ), .Y(n4588) );
  INVX1 U531 ( .A(\mem<3><2> ), .Y(n4587) );
  INVX1 U532 ( .A(\mem<3><3> ), .Y(n4586) );
  INVX1 U533 ( .A(\mem<3><4> ), .Y(n4585) );
  INVX1 U534 ( .A(\mem<3><5> ), .Y(n4584) );
  INVX1 U535 ( .A(\mem<3><6> ), .Y(n4583) );
  INVX1 U536 ( .A(\mem<3><7> ), .Y(n4582) );
  INVX1 U537 ( .A(\mem<2><0> ), .Y(n4581) );
  INVX1 U538 ( .A(\mem<2><1> ), .Y(n4580) );
  INVX1 U539 ( .A(\mem<2><2> ), .Y(n4579) );
  INVX1 U540 ( .A(\mem<2><3> ), .Y(n4578) );
  INVX1 U541 ( .A(\mem<2><4> ), .Y(n4577) );
  INVX1 U542 ( .A(\mem<2><5> ), .Y(n4576) );
  INVX1 U543 ( .A(\mem<2><6> ), .Y(n4575) );
  INVX1 U544 ( .A(\mem<2><7> ), .Y(n4574) );
  INVX1 U545 ( .A(\mem<1><0> ), .Y(n4573) );
  INVX1 U546 ( .A(\mem<1><1> ), .Y(n4572) );
  INVX1 U547 ( .A(\mem<1><2> ), .Y(n4571) );
  INVX1 U548 ( .A(\mem<1><3> ), .Y(n4570) );
  INVX1 U549 ( .A(\mem<1><4> ), .Y(n4569) );
  INVX1 U550 ( .A(\mem<1><5> ), .Y(n4568) );
  INVX1 U551 ( .A(\mem<1><6> ), .Y(n4567) );
  INVX1 U552 ( .A(\mem<1><7> ), .Y(n4566) );
  INVX1 U553 ( .A(n2777), .Y(n2781) );
  AND2X1 U554 ( .A(n271), .B(n97), .Y(n463) );
  AND2X1 U555 ( .A(n273), .B(n307), .Y(n1082) );
  INVX1 U556 ( .A(n705), .Y(n3269) );
  INVX1 U557 ( .A(n708), .Y(n3323) );
  INVX1 U558 ( .A(n2712), .Y(n2767) );
  AND2X1 U559 ( .A(n267), .B(n180), .Y(n424) );
  AND2X1 U560 ( .A(n275), .B(n226), .Y(n430) );
  AND2X1 U561 ( .A(n257), .B(n297), .Y(n1052) );
  INVX1 U562 ( .A(wr), .Y(n1658) );
  AND2X1 U563 ( .A(n261), .B(n301), .Y(n1064) );
  INVX1 U564 ( .A(n1531), .Y(n1529) );
  INVX1 U565 ( .A(n1532), .Y(n1528) );
  INVX1 U566 ( .A(n634), .Y(n3059) );
  INVX2 U567 ( .A(n1531), .Y(n1530) );
  INVX1 U568 ( .A(\mem<63><0> ), .Y(n5007) );
  INVX1 U569 ( .A(\mem<63><1> ), .Y(n5006) );
  INVX1 U570 ( .A(\mem<63><2> ), .Y(n5005) );
  INVX1 U571 ( .A(\mem<63><3> ), .Y(n5004) );
  INVX1 U572 ( .A(\mem<63><4> ), .Y(n5003) );
  INVX1 U573 ( .A(\mem<63><5> ), .Y(n5002) );
  INVX1 U574 ( .A(\mem<63><6> ), .Y(n5001) );
  INVX1 U575 ( .A(\mem<63><7> ), .Y(n5000) );
  INVX1 U576 ( .A(\data_in<0> ), .Y(n2983) );
  INVX1 U577 ( .A(n1621), .Y(n2981) );
  INVX1 U578 ( .A(\data_in<1> ), .Y(n2986) );
  INVX1 U579 ( .A(n1679), .Y(n2984) );
  INVX1 U580 ( .A(\data_in<2> ), .Y(n2989) );
  INVX1 U581 ( .A(n1709), .Y(n2987) );
  INVX1 U582 ( .A(\data_in<3> ), .Y(n2992) );
  INVX1 U583 ( .A(n1753), .Y(n2990) );
  INVX1 U584 ( .A(\data_in<4> ), .Y(n2995) );
  INVX1 U585 ( .A(n1800), .Y(n2993) );
  INVX1 U586 ( .A(\data_in<5> ), .Y(n2998) );
  INVX1 U587 ( .A(n2357), .Y(n2996) );
  INVX1 U588 ( .A(\data_in<6> ), .Y(n3001) );
  INVX1 U589 ( .A(n2402), .Y(n2999) );
  INVX1 U590 ( .A(\data_in<7> ), .Y(n3005) );
  INVX1 U591 ( .A(n2448), .Y(n3003) );
  INVX1 U592 ( .A(\data_in<0> ), .Y(n3010) );
  INVX1 U593 ( .A(n4999), .Y(n3008) );
  INVX1 U594 ( .A(\data_in<1> ), .Y(n3013) );
  INVX1 U595 ( .A(n4998), .Y(n3011) );
  INVX1 U596 ( .A(\data_in<2> ), .Y(n3016) );
  INVX1 U597 ( .A(n4997), .Y(n3014) );
  INVX1 U598 ( .A(\data_in<3> ), .Y(n3019) );
  INVX1 U599 ( .A(n4996), .Y(n3017) );
  INVX1 U600 ( .A(\data_in<4> ), .Y(n3022) );
  INVX1 U601 ( .A(n4995), .Y(n3020) );
  INVX1 U602 ( .A(\data_in<5> ), .Y(n3025) );
  INVX1 U603 ( .A(n4994), .Y(n3023) );
  INVX1 U604 ( .A(\data_in<6> ), .Y(n3028) );
  INVX1 U605 ( .A(n4993), .Y(n3026) );
  INVX1 U606 ( .A(\data_in<7> ), .Y(n3032) );
  INVX1 U607 ( .A(n4992), .Y(n3030) );
  INVX1 U608 ( .A(\data_in<0> ), .Y(n3036) );
  INVX1 U609 ( .A(n1618), .Y(n3034) );
  INVX1 U610 ( .A(\data_in<1> ), .Y(n3039) );
  INVX1 U611 ( .A(n1677), .Y(n3037) );
  INVX1 U612 ( .A(\data_in<2> ), .Y(n3042) );
  INVX1 U613 ( .A(n1708), .Y(n3040) );
  INVX1 U614 ( .A(\data_in<3> ), .Y(n3045) );
  INVX1 U615 ( .A(n1752), .Y(n3043) );
  INVX1 U616 ( .A(\data_in<4> ), .Y(n3048) );
  INVX1 U617 ( .A(n1798), .Y(n3046) );
  INVX1 U618 ( .A(\data_in<5> ), .Y(n3051) );
  INVX1 U619 ( .A(n2356), .Y(n3049) );
  INVX1 U620 ( .A(\data_in<6> ), .Y(n3054) );
  INVX1 U621 ( .A(n2401), .Y(n3052) );
  INVX1 U622 ( .A(\data_in<7> ), .Y(n3058) );
  INVX1 U623 ( .A(n2446), .Y(n3056) );
  INVX1 U624 ( .A(\data_in<0> ), .Y(n3063) );
  INVX1 U625 ( .A(n4991), .Y(n3061) );
  INVX1 U626 ( .A(\data_in<1> ), .Y(n3066) );
  INVX1 U627 ( .A(n4990), .Y(n3064) );
  INVX1 U628 ( .A(\data_in<2> ), .Y(n3069) );
  INVX1 U629 ( .A(n4989), .Y(n3067) );
  INVX1 U630 ( .A(\data_in<3> ), .Y(n3072) );
  INVX1 U631 ( .A(n4988), .Y(n3070) );
  INVX1 U632 ( .A(\data_in<4> ), .Y(n3075) );
  INVX1 U633 ( .A(n4987), .Y(n3073) );
  INVX1 U634 ( .A(\data_in<5> ), .Y(n3078) );
  INVX1 U635 ( .A(n4986), .Y(n3076) );
  INVX1 U636 ( .A(\data_in<6> ), .Y(n3081) );
  INVX1 U637 ( .A(n4985), .Y(n3079) );
  INVX1 U638 ( .A(\data_in<7> ), .Y(n3085) );
  INVX1 U639 ( .A(n4984), .Y(n3083) );
  INVX1 U640 ( .A(\data_in<0> ), .Y(n3090) );
  INVX1 U641 ( .A(n1608), .Y(n3088) );
  INVX1 U642 ( .A(\data_in<1> ), .Y(n3093) );
  INVX1 U643 ( .A(n1669), .Y(n3091) );
  INVX1 U644 ( .A(\data_in<2> ), .Y(n3096) );
  INVX1 U645 ( .A(n1713), .Y(n3094) );
  INVX1 U646 ( .A(\data_in<3> ), .Y(n3099) );
  INVX1 U647 ( .A(n1758), .Y(n3097) );
  INVX1 U648 ( .A(\data_in<4> ), .Y(n3102) );
  INVX1 U649 ( .A(n1806), .Y(n3100) );
  INVX1 U650 ( .A(\data_in<5> ), .Y(n3105) );
  INVX1 U651 ( .A(n2362), .Y(n3103) );
  INVX1 U652 ( .A(\data_in<6> ), .Y(n3108) );
  INVX1 U653 ( .A(n2406), .Y(n3106) );
  INVX1 U654 ( .A(\data_in<7> ), .Y(n3112) );
  INVX1 U655 ( .A(n2453), .Y(n3110) );
  INVX1 U656 ( .A(\data_in<0> ), .Y(n3118) );
  INVX1 U657 ( .A(n1605), .Y(n3116) );
  INVX1 U658 ( .A(\data_in<1> ), .Y(n3121) );
  INVX1 U659 ( .A(n1668), .Y(n3119) );
  INVX1 U660 ( .A(\data_in<2> ), .Y(n3124) );
  INVX1 U661 ( .A(n1712), .Y(n3122) );
  INVX1 U662 ( .A(\data_in<3> ), .Y(n3127) );
  INVX1 U663 ( .A(n1757), .Y(n3125) );
  INVX1 U664 ( .A(\data_in<4> ), .Y(n3130) );
  INVX1 U665 ( .A(n1804), .Y(n3128) );
  INVX1 U666 ( .A(\data_in<5> ), .Y(n3133) );
  INVX1 U667 ( .A(n2361), .Y(n3131) );
  INVX1 U668 ( .A(\data_in<6> ), .Y(n3136) );
  INVX1 U669 ( .A(n2405), .Y(n3134) );
  INVX1 U670 ( .A(\data_in<7> ), .Y(n3140) );
  INVX1 U671 ( .A(n2451), .Y(n3138) );
  INVX1 U672 ( .A(\data_in<0> ), .Y(n3144) );
  INVX1 U673 ( .A(n4983), .Y(n3142) );
  INVX1 U674 ( .A(\data_in<1> ), .Y(n3147) );
  INVX1 U675 ( .A(n4982), .Y(n3145) );
  INVX1 U676 ( .A(\data_in<2> ), .Y(n3150) );
  INVX1 U677 ( .A(n4981), .Y(n3148) );
  INVX1 U678 ( .A(\data_in<3> ), .Y(n3153) );
  INVX1 U679 ( .A(n4980), .Y(n3151) );
  INVX1 U680 ( .A(\data_in<4> ), .Y(n3156) );
  INVX1 U681 ( .A(n4979), .Y(n3154) );
  INVX1 U682 ( .A(\data_in<5> ), .Y(n3159) );
  INVX1 U683 ( .A(n4978), .Y(n3157) );
  INVX1 U684 ( .A(\data_in<6> ), .Y(n3162) );
  INVX1 U685 ( .A(n4977), .Y(n3160) );
  INVX1 U686 ( .A(\data_in<7> ), .Y(n3165) );
  INVX1 U687 ( .A(n4976), .Y(n3163) );
  INVX1 U688 ( .A(\data_in<0> ), .Y(n3171) );
  INVX1 U689 ( .A(n4975), .Y(n3169) );
  INVX1 U690 ( .A(\data_in<1> ), .Y(n3174) );
  INVX1 U691 ( .A(n4974), .Y(n3172) );
  INVX1 U692 ( .A(\data_in<2> ), .Y(n3177) );
  INVX1 U693 ( .A(n4973), .Y(n3175) );
  INVX1 U694 ( .A(\data_in<3> ), .Y(n3180) );
  INVX1 U695 ( .A(n4972), .Y(n3178) );
  INVX1 U696 ( .A(\data_in<4> ), .Y(n3183) );
  INVX1 U697 ( .A(n4971), .Y(n3181) );
  INVX1 U698 ( .A(\data_in<5> ), .Y(n3186) );
  INVX1 U699 ( .A(n4970), .Y(n3184) );
  INVX1 U700 ( .A(\data_in<6> ), .Y(n3189) );
  INVX1 U701 ( .A(n4969), .Y(n3187) );
  INVX1 U702 ( .A(\data_in<7> ), .Y(n3193) );
  INVX1 U703 ( .A(n4968), .Y(n3191) );
  INVX1 U704 ( .A(\data_in<0> ), .Y(n3196) );
  INVX1 U705 ( .A(n4967), .Y(n3194) );
  INVX1 U706 ( .A(\data_in<1> ), .Y(n3199) );
  INVX1 U707 ( .A(n4966), .Y(n3197) );
  INVX1 U708 ( .A(\data_in<2> ), .Y(n3202) );
  INVX1 U709 ( .A(n4965), .Y(n3200) );
  INVX1 U710 ( .A(\data_in<3> ), .Y(n3205) );
  INVX1 U711 ( .A(n4964), .Y(n3203) );
  INVX1 U712 ( .A(\data_in<4> ), .Y(n3208) );
  INVX1 U713 ( .A(n4963), .Y(n3206) );
  INVX1 U714 ( .A(\data_in<5> ), .Y(n3211) );
  INVX1 U715 ( .A(n4962), .Y(n3209) );
  INVX1 U716 ( .A(\data_in<6> ), .Y(n3214) );
  INVX1 U717 ( .A(n4961), .Y(n3212) );
  INVX1 U718 ( .A(\data_in<7> ), .Y(n3217) );
  INVX1 U719 ( .A(n4960), .Y(n3215) );
  INVX1 U720 ( .A(\data_in<0> ), .Y(n3221) );
  INVX1 U721 ( .A(n4959), .Y(n3219) );
  INVX1 U722 ( .A(\data_in<1> ), .Y(n3224) );
  INVX1 U723 ( .A(n4958), .Y(n3222) );
  INVX1 U724 ( .A(\data_in<2> ), .Y(n3227) );
  INVX1 U725 ( .A(n4957), .Y(n3225) );
  INVX1 U726 ( .A(\data_in<3> ), .Y(n3230) );
  INVX1 U727 ( .A(n4956), .Y(n3228) );
  INVX1 U728 ( .A(\data_in<4> ), .Y(n3233) );
  INVX1 U729 ( .A(n4955), .Y(n3231) );
  INVX1 U730 ( .A(\data_in<5> ), .Y(n3236) );
  INVX1 U731 ( .A(n4954), .Y(n3234) );
  INVX1 U732 ( .A(\data_in<6> ), .Y(n3239) );
  INVX1 U733 ( .A(n4953), .Y(n3237) );
  INVX1 U734 ( .A(\data_in<7> ), .Y(n3242) );
  INVX1 U735 ( .A(n4952), .Y(n3240) );
  INVX1 U736 ( .A(\data_in<0> ), .Y(n3246) );
  INVX1 U737 ( .A(n4951), .Y(n3244) );
  INVX1 U738 ( .A(\data_in<1> ), .Y(n3249) );
  INVX1 U739 ( .A(n4950), .Y(n3247) );
  INVX1 U740 ( .A(\data_in<2> ), .Y(n3252) );
  INVX1 U741 ( .A(n4949), .Y(n3250) );
  INVX1 U742 ( .A(\data_in<3> ), .Y(n3255) );
  INVX1 U743 ( .A(n4948), .Y(n3253) );
  INVX1 U744 ( .A(\data_in<4> ), .Y(n3258) );
  INVX1 U745 ( .A(n4947), .Y(n3256) );
  INVX1 U746 ( .A(\data_in<5> ), .Y(n3261) );
  INVX1 U747 ( .A(n4946), .Y(n3259) );
  INVX1 U748 ( .A(\data_in<6> ), .Y(n3264) );
  INVX1 U749 ( .A(n4945), .Y(n3262) );
  INVX1 U750 ( .A(\data_in<7> ), .Y(n3268) );
  INVX1 U751 ( .A(n4944), .Y(n3266) );
  INVX1 U752 ( .A(\data_in<0> ), .Y(n3273) );
  INVX1 U753 ( .A(n4943), .Y(n3271) );
  INVX1 U754 ( .A(\data_in<1> ), .Y(n3276) );
  INVX1 U755 ( .A(n4942), .Y(n3274) );
  INVX1 U756 ( .A(\data_in<2> ), .Y(n3279) );
  INVX1 U757 ( .A(n4941), .Y(n3277) );
  INVX1 U758 ( .A(\data_in<3> ), .Y(n3282) );
  INVX1 U759 ( .A(n4940), .Y(n3280) );
  INVX1 U760 ( .A(\data_in<4> ), .Y(n3285) );
  INVX1 U761 ( .A(n4939), .Y(n3283) );
  INVX1 U762 ( .A(\data_in<5> ), .Y(n3288) );
  INVX1 U763 ( .A(n4938), .Y(n3286) );
  INVX1 U764 ( .A(\data_in<6> ), .Y(n3291) );
  INVX1 U765 ( .A(n4937), .Y(n3289) );
  INVX1 U766 ( .A(\data_in<7> ), .Y(n3295) );
  INVX1 U767 ( .A(n4936), .Y(n3293) );
  INVX1 U768 ( .A(\data_in<0> ), .Y(n3300) );
  INVX1 U769 ( .A(n4935), .Y(n3298) );
  INVX1 U770 ( .A(\data_in<1> ), .Y(n3303) );
  INVX1 U771 ( .A(n4934), .Y(n3301) );
  INVX1 U772 ( .A(\data_in<2> ), .Y(n3306) );
  INVX1 U773 ( .A(n4933), .Y(n3304) );
  INVX1 U774 ( .A(\data_in<3> ), .Y(n3309) );
  INVX1 U775 ( .A(n4932), .Y(n3307) );
  INVX1 U776 ( .A(\data_in<4> ), .Y(n3312) );
  INVX1 U777 ( .A(n4931), .Y(n3310) );
  INVX1 U778 ( .A(\data_in<5> ), .Y(n3315) );
  INVX1 U779 ( .A(n4930), .Y(n3313) );
  INVX1 U780 ( .A(\data_in<6> ), .Y(n3318) );
  INVX1 U781 ( .A(n4929), .Y(n3316) );
  INVX1 U782 ( .A(\data_in<7> ), .Y(n3322) );
  INVX1 U783 ( .A(n4928), .Y(n3320) );
  INVX1 U784 ( .A(\data_in<0> ), .Y(n3328) );
  INVX1 U785 ( .A(n4927), .Y(n3326) );
  INVX1 U786 ( .A(\data_in<1> ), .Y(n3331) );
  INVX1 U787 ( .A(n4926), .Y(n3329) );
  INVX1 U788 ( .A(\data_in<2> ), .Y(n3334) );
  INVX1 U789 ( .A(n4925), .Y(n3332) );
  INVX1 U790 ( .A(\data_in<3> ), .Y(n3337) );
  INVX1 U791 ( .A(n4924), .Y(n3335) );
  INVX1 U792 ( .A(\data_in<4> ), .Y(n3340) );
  INVX1 U793 ( .A(n4923), .Y(n3338) );
  INVX1 U794 ( .A(\data_in<5> ), .Y(n3343) );
  INVX1 U795 ( .A(n4922), .Y(n3341) );
  INVX1 U796 ( .A(\data_in<6> ), .Y(n3346) );
  INVX1 U797 ( .A(n4921), .Y(n3344) );
  INVX1 U798 ( .A(\data_in<7> ), .Y(n3350) );
  INVX1 U799 ( .A(n4920), .Y(n3348) );
  INVX1 U800 ( .A(\data_in<0> ), .Y(n3353) );
  INVX1 U801 ( .A(n4919), .Y(n3351) );
  INVX1 U802 ( .A(\data_in<1> ), .Y(n3356) );
  INVX1 U803 ( .A(n4918), .Y(n3354) );
  INVX1 U804 ( .A(\data_in<2> ), .Y(n3359) );
  INVX1 U805 ( .A(n4917), .Y(n3357) );
  INVX1 U806 ( .A(\data_in<3> ), .Y(n3362) );
  INVX1 U807 ( .A(n4916), .Y(n3360) );
  INVX1 U808 ( .A(\data_in<4> ), .Y(n3365) );
  INVX1 U809 ( .A(n4915), .Y(n3363) );
  INVX1 U810 ( .A(\data_in<5> ), .Y(n3368) );
  INVX1 U811 ( .A(n4914), .Y(n3366) );
  INVX1 U812 ( .A(\data_in<6> ), .Y(n3371) );
  INVX1 U813 ( .A(n4913), .Y(n3369) );
  INVX1 U814 ( .A(\data_in<7> ), .Y(n3374) );
  INVX1 U815 ( .A(n4912), .Y(n3372) );
  INVX1 U816 ( .A(\data_in<0> ), .Y(n3378) );
  INVX1 U818 ( .A(n4911), .Y(n3376) );
  INVX1 U820 ( .A(\data_in<1> ), .Y(n3381) );
  INVX1 U822 ( .A(n4910), .Y(n3379) );
  INVX1 U824 ( .A(\data_in<2> ), .Y(n3384) );
  INVX1 U826 ( .A(n4909), .Y(n3382) );
  INVX1 U828 ( .A(\data_in<3> ), .Y(n3387) );
  INVX1 U830 ( .A(n4908), .Y(n3385) );
  INVX1 U832 ( .A(\data_in<4> ), .Y(n3390) );
  INVX1 U833 ( .A(n4907), .Y(n3388) );
  INVX1 U834 ( .A(\data_in<5> ), .Y(n3393) );
  INVX1 U835 ( .A(n4906), .Y(n3391) );
  INVX1 U836 ( .A(\data_in<6> ), .Y(n3396) );
  INVX1 U837 ( .A(n4905), .Y(n3394) );
  INVX1 U838 ( .A(\data_in<7> ), .Y(n3399) );
  INVX1 U839 ( .A(n4904), .Y(n3397) );
  INVX1 U840 ( .A(\data_in<0> ), .Y(n3402) );
  INVX1 U841 ( .A(n4903), .Y(n3400) );
  INVX1 U842 ( .A(\data_in<1> ), .Y(n3405) );
  INVX1 U843 ( .A(n4902), .Y(n3403) );
  INVX1 U844 ( .A(\data_in<2> ), .Y(n3408) );
  INVX1 U845 ( .A(n4901), .Y(n3406) );
  INVX1 U846 ( .A(\data_in<3> ), .Y(n3411) );
  INVX1 U847 ( .A(n4900), .Y(n3409) );
  INVX1 U848 ( .A(\data_in<4> ), .Y(n3414) );
  INVX1 U849 ( .A(n4899), .Y(n3412) );
  INVX1 U850 ( .A(\data_in<5> ), .Y(n3417) );
  INVX1 U851 ( .A(n4898), .Y(n3415) );
  INVX1 U852 ( .A(\data_in<6> ), .Y(n3420) );
  INVX1 U853 ( .A(n4897), .Y(n3418) );
  INVX1 U854 ( .A(\data_in<7> ), .Y(n3423) );
  INVX1 U855 ( .A(n4896), .Y(n3421) );
  INVX1 U856 ( .A(\data_in<0> ), .Y(n3426) );
  INVX1 U857 ( .A(n4895), .Y(n3424) );
  INVX1 U858 ( .A(\data_in<1> ), .Y(n3429) );
  INVX1 U859 ( .A(n4894), .Y(n3427) );
  INVX1 U860 ( .A(\data_in<2> ), .Y(n3432) );
  INVX1 U861 ( .A(n4893), .Y(n3430) );
  INVX1 U862 ( .A(\data_in<3> ), .Y(n3435) );
  INVX1 U863 ( .A(n4892), .Y(n3433) );
  INVX1 U864 ( .A(\data_in<4> ), .Y(n3438) );
  INVX1 U865 ( .A(n4891), .Y(n3436) );
  INVX1 U866 ( .A(\data_in<5> ), .Y(n3441) );
  INVX1 U867 ( .A(n4890), .Y(n3439) );
  INVX1 U868 ( .A(\data_in<6> ), .Y(n3444) );
  INVX1 U869 ( .A(n4889), .Y(n3442) );
  INVX1 U870 ( .A(\data_in<7> ), .Y(n3447) );
  INVX1 U871 ( .A(n4888), .Y(n3445) );
  INVX1 U872 ( .A(\data_in<0> ), .Y(n3450) );
  INVX1 U873 ( .A(n4887), .Y(n3448) );
  INVX1 U874 ( .A(\data_in<1> ), .Y(n3453) );
  INVX1 U875 ( .A(n4886), .Y(n3451) );
  INVX1 U876 ( .A(\data_in<2> ), .Y(n3456) );
  INVX1 U877 ( .A(n4885), .Y(n3454) );
  INVX1 U878 ( .A(\data_in<3> ), .Y(n3459) );
  INVX1 U879 ( .A(n4884), .Y(n3457) );
  INVX1 U880 ( .A(\data_in<4> ), .Y(n3462) );
  INVX1 U881 ( .A(n4883), .Y(n3460) );
  INVX1 U882 ( .A(\data_in<5> ), .Y(n3465) );
  INVX1 U883 ( .A(n4882), .Y(n3463) );
  INVX1 U884 ( .A(\data_in<6> ), .Y(n3468) );
  INVX1 U885 ( .A(n4881), .Y(n3466) );
  INVX1 U886 ( .A(\data_in<7> ), .Y(n3471) );
  INVX1 U887 ( .A(n4880), .Y(n3469) );
  INVX1 U888 ( .A(\data_in<0> ), .Y(n3475) );
  INVX1 U889 ( .A(n4879), .Y(n3473) );
  INVX1 U890 ( .A(\data_in<1> ), .Y(n3478) );
  INVX1 U891 ( .A(n4878), .Y(n3476) );
  INVX1 U892 ( .A(\data_in<2> ), .Y(n3481) );
  INVX1 U893 ( .A(n4877), .Y(n3479) );
  INVX1 U894 ( .A(\data_in<3> ), .Y(n3484) );
  INVX1 U895 ( .A(n4876), .Y(n3482) );
  INVX1 U896 ( .A(\data_in<4> ), .Y(n3487) );
  INVX1 U897 ( .A(n4875), .Y(n3485) );
  INVX1 U898 ( .A(\data_in<5> ), .Y(n3490) );
  INVX1 U899 ( .A(n4874), .Y(n3488) );
  INVX1 U900 ( .A(\data_in<6> ), .Y(n3493) );
  INVX1 U901 ( .A(n4873), .Y(n3491) );
  INVX1 U902 ( .A(\data_in<7> ), .Y(n3496) );
  INVX1 U903 ( .A(n4872), .Y(n3494) );
  INVX1 U904 ( .A(\data_in<0> ), .Y(n3500) );
  INVX1 U905 ( .A(n4871), .Y(n3498) );
  INVX1 U906 ( .A(\data_in<1> ), .Y(n3503) );
  INVX1 U907 ( .A(n4870), .Y(n3501) );
  INVX1 U908 ( .A(\data_in<2> ), .Y(n3506) );
  INVX1 U909 ( .A(n4869), .Y(n3504) );
  INVX1 U910 ( .A(\data_in<3> ), .Y(n3509) );
  INVX1 U911 ( .A(n4868), .Y(n3507) );
  INVX1 U912 ( .A(\data_in<4> ), .Y(n3512) );
  INVX1 U913 ( .A(n4867), .Y(n3510) );
  INVX1 U914 ( .A(\data_in<5> ), .Y(n3515) );
  INVX1 U915 ( .A(n4866), .Y(n3513) );
  INVX1 U916 ( .A(\data_in<6> ), .Y(n3518) );
  INVX1 U917 ( .A(n4865), .Y(n3516) );
  INVX1 U918 ( .A(\data_in<7> ), .Y(n3521) );
  INVX1 U919 ( .A(n4864), .Y(n3519) );
  INVX1 U920 ( .A(\data_in<0> ), .Y(n3524) );
  INVX1 U921 ( .A(n4863), .Y(n3522) );
  INVX1 U922 ( .A(\data_in<1> ), .Y(n3527) );
  INVX1 U923 ( .A(n4862), .Y(n3525) );
  INVX1 U924 ( .A(\data_in<2> ), .Y(n3530) );
  INVX1 U925 ( .A(n4861), .Y(n3528) );
  INVX1 U926 ( .A(\data_in<3> ), .Y(n3533) );
  INVX1 U927 ( .A(n4860), .Y(n3531) );
  INVX1 U928 ( .A(\data_in<4> ), .Y(n3536) );
  INVX1 U929 ( .A(n4859), .Y(n3534) );
  INVX1 U930 ( .A(\data_in<5> ), .Y(n3539) );
  INVX1 U931 ( .A(n4858), .Y(n3537) );
  INVX1 U932 ( .A(\data_in<6> ), .Y(n3542) );
  INVX1 U933 ( .A(n4857), .Y(n3540) );
  INVX1 U934 ( .A(\data_in<7> ), .Y(n3545) );
  INVX1 U935 ( .A(n4856), .Y(n3543) );
  INVX1 U936 ( .A(\data_in<0> ), .Y(n3549) );
  INVX1 U937 ( .A(n4855), .Y(n3547) );
  INVX1 U938 ( .A(\data_in<1> ), .Y(n3552) );
  INVX1 U939 ( .A(n4854), .Y(n3550) );
  INVX1 U940 ( .A(\data_in<2> ), .Y(n3555) );
  INVX1 U941 ( .A(n4853), .Y(n3553) );
  INVX1 U942 ( .A(\data_in<3> ), .Y(n3558) );
  INVX1 U943 ( .A(n4852), .Y(n3556) );
  INVX1 U944 ( .A(\data_in<4> ), .Y(n3561) );
  INVX1 U945 ( .A(n4851), .Y(n3559) );
  INVX1 U946 ( .A(\data_in<5> ), .Y(n3564) );
  INVX1 U947 ( .A(n4850), .Y(n3562) );
  INVX1 U948 ( .A(\data_in<6> ), .Y(n3567) );
  INVX1 U949 ( .A(n4849), .Y(n3565) );
  INVX1 U950 ( .A(\data_in<7> ), .Y(n3570) );
  INVX1 U951 ( .A(n4848), .Y(n3568) );
  INVX1 U952 ( .A(\data_in<0> ), .Y(n3574) );
  INVX1 U953 ( .A(n4847), .Y(n3572) );
  INVX1 U954 ( .A(\data_in<1> ), .Y(n3577) );
  INVX1 U955 ( .A(n4846), .Y(n3575) );
  INVX1 U956 ( .A(\data_in<2> ), .Y(n3580) );
  INVX1 U957 ( .A(n4845), .Y(n3578) );
  INVX1 U958 ( .A(\data_in<3> ), .Y(n3583) );
  INVX1 U959 ( .A(n4844), .Y(n3581) );
  INVX1 U960 ( .A(\data_in<4> ), .Y(n3586) );
  INVX1 U961 ( .A(n4843), .Y(n3584) );
  INVX1 U962 ( .A(\data_in<5> ), .Y(n3589) );
  INVX1 U963 ( .A(n4842), .Y(n3587) );
  INVX1 U964 ( .A(\data_in<6> ), .Y(n3592) );
  INVX1 U965 ( .A(n4841), .Y(n3590) );
  INVX1 U966 ( .A(\data_in<7> ), .Y(n3595) );
  INVX1 U967 ( .A(n4840), .Y(n3593) );
  INVX1 U968 ( .A(\data_in<0> ), .Y(n3598) );
  INVX1 U969 ( .A(n4839), .Y(n3596) );
  INVX1 U970 ( .A(\data_in<1> ), .Y(n3601) );
  INVX1 U971 ( .A(n4838), .Y(n3599) );
  INVX1 U972 ( .A(\data_in<2> ), .Y(n3604) );
  INVX1 U973 ( .A(n4837), .Y(n3602) );
  INVX1 U974 ( .A(\data_in<3> ), .Y(n3607) );
  INVX1 U975 ( .A(n4836), .Y(n3605) );
  INVX1 U976 ( .A(\data_in<4> ), .Y(n3610) );
  INVX1 U977 ( .A(n4835), .Y(n3608) );
  INVX1 U978 ( .A(\data_in<5> ), .Y(n3613) );
  INVX1 U979 ( .A(n4834), .Y(n3611) );
  INVX1 U980 ( .A(\data_in<6> ), .Y(n3616) );
  INVX1 U981 ( .A(n4833), .Y(n3614) );
  INVX1 U982 ( .A(\data_in<7> ), .Y(n3619) );
  INVX1 U983 ( .A(n4832), .Y(n3617) );
  INVX1 U984 ( .A(\data_in<0> ), .Y(n3623) );
  INVX1 U985 ( .A(n4831), .Y(n3621) );
  INVX1 U986 ( .A(\data_in<1> ), .Y(n3626) );
  INVX1 U987 ( .A(n4830), .Y(n3624) );
  INVX1 U988 ( .A(\data_in<2> ), .Y(n3629) );
  INVX1 U989 ( .A(n4829), .Y(n3627) );
  INVX1 U990 ( .A(\data_in<3> ), .Y(n3632) );
  INVX1 U991 ( .A(n4828), .Y(n3630) );
  INVX1 U992 ( .A(\data_in<4> ), .Y(n3635) );
  INVX1 U993 ( .A(n4827), .Y(n3633) );
  INVX1 U994 ( .A(\data_in<5> ), .Y(n3638) );
  INVX1 U995 ( .A(n4826), .Y(n3636) );
  INVX1 U996 ( .A(\data_in<6> ), .Y(n3641) );
  INVX1 U997 ( .A(n4825), .Y(n3639) );
  INVX1 U998 ( .A(\data_in<7> ), .Y(n3644) );
  INVX1 U999 ( .A(n4824), .Y(n3642) );
  INVX1 U1000 ( .A(\data_in<0> ), .Y(n3647) );
  INVX1 U1001 ( .A(n4823), .Y(n3645) );
  INVX1 U1002 ( .A(\data_in<1> ), .Y(n3650) );
  INVX1 U1003 ( .A(n4822), .Y(n3648) );
  INVX1 U1004 ( .A(\data_in<2> ), .Y(n3653) );
  INVX1 U1005 ( .A(n4821), .Y(n3651) );
  INVX1 U1006 ( .A(\data_in<3> ), .Y(n3656) );
  INVX1 U1007 ( .A(n4820), .Y(n3654) );
  INVX1 U1008 ( .A(\data_in<4> ), .Y(n3659) );
  INVX1 U1009 ( .A(n4819), .Y(n3657) );
  INVX1 U1010 ( .A(\data_in<5> ), .Y(n3662) );
  INVX1 U1011 ( .A(n4818), .Y(n3660) );
  INVX1 U1012 ( .A(\data_in<6> ), .Y(n3665) );
  INVX1 U1013 ( .A(n4817), .Y(n3663) );
  INVX1 U1014 ( .A(\data_in<7> ), .Y(n3668) );
  INVX1 U1015 ( .A(n4816), .Y(n3666) );
  INVX1 U1016 ( .A(\data_in<0> ), .Y(n3672) );
  INVX1 U1017 ( .A(n4815), .Y(n3670) );
  INVX1 U1018 ( .A(\data_in<1> ), .Y(n3675) );
  INVX1 U1019 ( .A(n4814), .Y(n3673) );
  INVX1 U1020 ( .A(\data_in<2> ), .Y(n3678) );
  INVX1 U1021 ( .A(n4813), .Y(n3676) );
  INVX1 U1022 ( .A(\data_in<3> ), .Y(n3681) );
  INVX1 U1023 ( .A(n4812), .Y(n3679) );
  INVX1 U1024 ( .A(\data_in<4> ), .Y(n3684) );
  INVX1 U1025 ( .A(n4811), .Y(n3682) );
  INVX1 U1026 ( .A(\data_in<5> ), .Y(n3687) );
  INVX1 U1027 ( .A(n4810), .Y(n3685) );
  INVX1 U1028 ( .A(\data_in<6> ), .Y(n3690) );
  INVX1 U1029 ( .A(n4809), .Y(n3688) );
  INVX1 U1030 ( .A(\data_in<7> ), .Y(n3693) );
  INVX1 U1031 ( .A(n4808), .Y(n3691) );
  INVX1 U1032 ( .A(\data_in<0> ), .Y(n3696) );
  INVX1 U1033 ( .A(n4807), .Y(n3694) );
  INVX1 U1034 ( .A(\data_in<1> ), .Y(n3699) );
  INVX1 U1035 ( .A(n4806), .Y(n3697) );
  INVX1 U1036 ( .A(\data_in<2> ), .Y(n3702) );
  INVX1 U1037 ( .A(n4805), .Y(n3700) );
  INVX1 U1038 ( .A(\data_in<3> ), .Y(n3705) );
  INVX1 U1039 ( .A(n4804), .Y(n3703) );
  INVX1 U1040 ( .A(\data_in<4> ), .Y(n3708) );
  INVX1 U1041 ( .A(n4803), .Y(n3706) );
  INVX1 U1042 ( .A(\data_in<5> ), .Y(n3711) );
  INVX1 U1043 ( .A(n4802), .Y(n3709) );
  INVX1 U1044 ( .A(\data_in<6> ), .Y(n3714) );
  INVX1 U1045 ( .A(n4801), .Y(n3712) );
  INVX1 U1046 ( .A(\data_in<7> ), .Y(n3717) );
  INVX1 U1047 ( .A(n4800), .Y(n3715) );
  INVX1 U1048 ( .A(\data_in<0> ), .Y(n3721) );
  INVX1 U1049 ( .A(n4799), .Y(n3719) );
  INVX1 U1050 ( .A(\data_in<1> ), .Y(n3724) );
  INVX1 U1051 ( .A(n4798), .Y(n3722) );
  INVX1 U1052 ( .A(\data_in<2> ), .Y(n3727) );
  INVX1 U1053 ( .A(n4797), .Y(n3725) );
  INVX1 U1054 ( .A(\data_in<3> ), .Y(n3730) );
  INVX1 U1055 ( .A(n4796), .Y(n3728) );
  INVX1 U1056 ( .A(\data_in<4> ), .Y(n3733) );
  INVX1 U1057 ( .A(n4795), .Y(n3731) );
  INVX1 U1058 ( .A(\data_in<5> ), .Y(n3736) );
  INVX1 U1059 ( .A(n4794), .Y(n3734) );
  INVX1 U1060 ( .A(\data_in<6> ), .Y(n3739) );
  INVX1 U1061 ( .A(n4793), .Y(n3737) );
  INVX1 U1062 ( .A(\data_in<7> ), .Y(n3742) );
  INVX1 U1063 ( .A(n4792), .Y(n3740) );
  INVX1 U1064 ( .A(\data_in<0> ), .Y(n3745) );
  INVX1 U1065 ( .A(n4791), .Y(n3743) );
  INVX1 U1066 ( .A(\data_in<1> ), .Y(n3748) );
  INVX1 U1067 ( .A(n4790), .Y(n3746) );
  INVX1 U1068 ( .A(\data_in<2> ), .Y(n3751) );
  INVX1 U1069 ( .A(n4789), .Y(n3749) );
  INVX1 U1070 ( .A(\data_in<3> ), .Y(n3754) );
  INVX1 U1071 ( .A(n4788), .Y(n3752) );
  INVX1 U1072 ( .A(\data_in<4> ), .Y(n3757) );
  INVX1 U1073 ( .A(n4787), .Y(n3755) );
  INVX1 U1074 ( .A(\data_in<5> ), .Y(n3760) );
  INVX1 U1075 ( .A(n4786), .Y(n3758) );
  INVX1 U1076 ( .A(\data_in<6> ), .Y(n3763) );
  INVX1 U1077 ( .A(n4785), .Y(n3761) );
  INVX1 U1078 ( .A(\data_in<7> ), .Y(n3766) );
  INVX1 U1079 ( .A(n4784), .Y(n3764) );
  INVX1 U1080 ( .A(\data_in<0> ), .Y(n3770) );
  INVX1 U1081 ( .A(n1641), .Y(n3768) );
  INVX1 U1082 ( .A(\data_in<1> ), .Y(n3773) );
  INVX1 U1083 ( .A(n4783), .Y(n3771) );
  INVX1 U1084 ( .A(\data_in<2> ), .Y(n3776) );
  INVX1 U1085 ( .A(n4782), .Y(n3774) );
  INVX1 U1086 ( .A(\data_in<3> ), .Y(n3779) );
  INVX1 U1087 ( .A(n4781), .Y(n3777) );
  INVX1 U1088 ( .A(\data_in<4> ), .Y(n3782) );
  INVX1 U1089 ( .A(n4780), .Y(n3780) );
  INVX1 U1090 ( .A(\data_in<5> ), .Y(n3785) );
  INVX1 U1091 ( .A(n4779), .Y(n3783) );
  INVX1 U1092 ( .A(\data_in<6> ), .Y(n3788) );
  INVX1 U1093 ( .A(n4778), .Y(n3786) );
  INVX1 U1094 ( .A(\data_in<7> ), .Y(n3792) );
  INVX1 U1095 ( .A(n4777), .Y(n3790) );
  INVX1 U1096 ( .A(\data_in<0> ), .Y(n3798) );
  INVX1 U1097 ( .A(n4776), .Y(n3796) );
  INVX1 U1098 ( .A(\data_in<1> ), .Y(n3801) );
  INVX1 U1099 ( .A(n4775), .Y(n3799) );
  INVX1 U1100 ( .A(\data_in<2> ), .Y(n3804) );
  INVX1 U1101 ( .A(n1723), .Y(n3802) );
  INVX1 U1102 ( .A(\data_in<3> ), .Y(n3807) );
  INVX1 U1103 ( .A(n1768), .Y(n3805) );
  INVX1 U1104 ( .A(\data_in<4> ), .Y(n3810) );
  INVX1 U1105 ( .A(n1815), .Y(n3808) );
  INVX1 U1106 ( .A(\data_in<5> ), .Y(n3813) );
  INVX1 U1107 ( .A(n2372), .Y(n3811) );
  INVX1 U1108 ( .A(\data_in<6> ), .Y(n3816) );
  INVX1 U1109 ( .A(n2416), .Y(n3814) );
  INVX1 U1110 ( .A(\data_in<7> ), .Y(n3820) );
  INVX1 U1111 ( .A(n2463), .Y(n3818) );
  INVX1 U1112 ( .A(\data_in<0> ), .Y(n3824) );
  INVX1 U1113 ( .A(n1639), .Y(n3822) );
  INVX1 U1114 ( .A(\data_in<1> ), .Y(n3827) );
  INVX1 U1115 ( .A(n4774), .Y(n3825) );
  INVX1 U1116 ( .A(\data_in<2> ), .Y(n3830) );
  INVX1 U1117 ( .A(n4773), .Y(n3828) );
  INVX1 U1118 ( .A(\data_in<3> ), .Y(n3833) );
  INVX1 U1119 ( .A(n4772), .Y(n3831) );
  INVX1 U1120 ( .A(\data_in<4> ), .Y(n3836) );
  INVX1 U1121 ( .A(n4771), .Y(n3834) );
  INVX1 U1122 ( .A(\data_in<5> ), .Y(n3839) );
  INVX1 U1123 ( .A(n4770), .Y(n3837) );
  INVX1 U1124 ( .A(\data_in<6> ), .Y(n3842) );
  INVX1 U1125 ( .A(n4769), .Y(n3840) );
  INVX1 U1126 ( .A(\data_in<7> ), .Y(n3846) );
  INVX1 U1127 ( .A(n4768), .Y(n3844) );
  INVX1 U1128 ( .A(\data_in<0> ), .Y(n3850) );
  INVX1 U1129 ( .A(n4767), .Y(n3848) );
  INVX1 U1130 ( .A(\data_in<1> ), .Y(n3853) );
  INVX1 U1131 ( .A(n4766), .Y(n3851) );
  INVX1 U1132 ( .A(\data_in<2> ), .Y(n3856) );
  INVX1 U1133 ( .A(n1721), .Y(n3854) );
  INVX1 U1134 ( .A(\data_in<3> ), .Y(n3859) );
  INVX1 U1135 ( .A(n1766), .Y(n3857) );
  INVX1 U1136 ( .A(\data_in<4> ), .Y(n3862) );
  INVX1 U1137 ( .A(n1813), .Y(n3860) );
  INVX1 U1138 ( .A(\data_in<5> ), .Y(n3865) );
  INVX1 U1139 ( .A(n2370), .Y(n3863) );
  INVX1 U1140 ( .A(\data_in<6> ), .Y(n3868) );
  INVX1 U1141 ( .A(n2414), .Y(n3866) );
  INVX1 U1142 ( .A(\data_in<7> ), .Y(n3872) );
  INVX1 U1143 ( .A(n2461), .Y(n3870) );
  INVX1 U1144 ( .A(\data_in<0> ), .Y(n3876) );
  INVX1 U1145 ( .A(n1631), .Y(n3874) );
  INVX1 U1146 ( .A(\data_in<1> ), .Y(n3879) );
  INVX1 U1147 ( .A(n1684), .Y(n3877) );
  INVX1 U1148 ( .A(\data_in<2> ), .Y(n3882) );
  INVX1 U1149 ( .A(n4765), .Y(n3880) );
  INVX1 U1150 ( .A(\data_in<3> ), .Y(n3885) );
  INVX1 U1151 ( .A(n4764), .Y(n3883) );
  INVX1 U1152 ( .A(\data_in<4> ), .Y(n3888) );
  INVX1 U1153 ( .A(n4763), .Y(n3886) );
  INVX1 U1154 ( .A(\data_in<5> ), .Y(n3891) );
  INVX1 U1155 ( .A(n4762), .Y(n3889) );
  INVX1 U1156 ( .A(\data_in<6> ), .Y(n3894) );
  INVX1 U1157 ( .A(n4761), .Y(n3892) );
  INVX1 U1158 ( .A(\data_in<7> ), .Y(n3898) );
  INVX1 U1159 ( .A(n4760), .Y(n3896) );
  INVX1 U1160 ( .A(\data_in<0> ), .Y(n3903) );
  INVX1 U1161 ( .A(n4759), .Y(n3901) );
  INVX1 U1162 ( .A(\data_in<1> ), .Y(n3906) );
  INVX1 U1163 ( .A(n4758), .Y(n3904) );
  INVX1 U1164 ( .A(\data_in<2> ), .Y(n3909) );
  INVX1 U1165 ( .A(n1727), .Y(n3907) );
  INVX1 U1166 ( .A(\data_in<3> ), .Y(n3912) );
  INVX1 U1167 ( .A(n1772), .Y(n3910) );
  INVX1 U1168 ( .A(\data_in<4> ), .Y(n3915) );
  INVX1 U1169 ( .A(n2331), .Y(n3913) );
  INVX1 U1170 ( .A(\data_in<5> ), .Y(n3918) );
  INVX1 U1171 ( .A(n2377), .Y(n3916) );
  INVX1 U1172 ( .A(\data_in<6> ), .Y(n3921) );
  INVX1 U1173 ( .A(n2421), .Y(n3919) );
  INVX1 U1174 ( .A(\data_in<7> ), .Y(n3925) );
  INVX1 U1175 ( .A(n2468), .Y(n3923) );
  INVX1 U1176 ( .A(\data_in<0> ), .Y(n3930) );
  INVX1 U1177 ( .A(n1630), .Y(n3928) );
  INVX1 U1178 ( .A(\data_in<1> ), .Y(n3933) );
  INVX1 U1179 ( .A(n1683), .Y(n3931) );
  INVX1 U1180 ( .A(\data_in<2> ), .Y(n3936) );
  INVX1 U1181 ( .A(n1726), .Y(n3934) );
  INVX1 U1182 ( .A(\data_in<3> ), .Y(n3939) );
  INVX1 U1183 ( .A(n1771), .Y(n3937) );
  INVX1 U1184 ( .A(\data_in<4> ), .Y(n3942) );
  INVX1 U1185 ( .A(n2330), .Y(n3940) );
  INVX1 U1186 ( .A(\data_in<5> ), .Y(n3945) );
  INVX1 U1187 ( .A(n2375), .Y(n3943) );
  INVX1 U1188 ( .A(\data_in<6> ), .Y(n3948) );
  INVX1 U1189 ( .A(n2419), .Y(n3946) );
  INVX1 U1190 ( .A(\data_in<7> ), .Y(n3952) );
  INVX1 U1191 ( .A(n2466), .Y(n3950) );
  INVX1 U1192 ( .A(\data_in<0> ), .Y(n3955) );
  INVX1 U1193 ( .A(n4757), .Y(n3953) );
  INVX1 U1194 ( .A(\data_in<1> ), .Y(n3958) );
  INVX1 U1195 ( .A(n4756), .Y(n3956) );
  INVX1 U1196 ( .A(\data_in<2> ), .Y(n3961) );
  INVX1 U1197 ( .A(n4755), .Y(n3959) );
  INVX1 U1198 ( .A(\data_in<3> ), .Y(n3964) );
  INVX1 U1199 ( .A(n4754), .Y(n3962) );
  INVX1 U1200 ( .A(\data_in<4> ), .Y(n3967) );
  INVX1 U1201 ( .A(n4753), .Y(n3965) );
  INVX1 U1202 ( .A(\data_in<5> ), .Y(n3970) );
  INVX1 U1203 ( .A(n4752), .Y(n3968) );
  INVX1 U1204 ( .A(\data_in<6> ), .Y(n3973) );
  INVX1 U1205 ( .A(n4751), .Y(n3971) );
  INVX1 U1206 ( .A(\data_in<7> ), .Y(n3976) );
  INVX1 U1207 ( .A(n4750), .Y(n3974) );
  INVX1 U1208 ( .A(\data_in<0> ), .Y(n3979) );
  INVX1 U1209 ( .A(n4749), .Y(n3977) );
  INVX1 U1210 ( .A(\data_in<1> ), .Y(n3982) );
  INVX1 U1211 ( .A(n4748), .Y(n3980) );
  INVX1 U1212 ( .A(\data_in<2> ), .Y(n3985) );
  INVX1 U1213 ( .A(n4747), .Y(n3983) );
  INVX1 U1214 ( .A(\data_in<3> ), .Y(n3988) );
  INVX1 U1215 ( .A(n4746), .Y(n3986) );
  INVX1 U1216 ( .A(\data_in<4> ), .Y(n3991) );
  INVX1 U1217 ( .A(n4745), .Y(n3989) );
  INVX1 U1218 ( .A(\data_in<5> ), .Y(n3994) );
  INVX1 U1219 ( .A(n4744), .Y(n3992) );
  INVX1 U1220 ( .A(\data_in<6> ), .Y(n3997) );
  INVX1 U1221 ( .A(n4743), .Y(n3995) );
  INVX1 U1222 ( .A(\data_in<7> ), .Y(n4000) );
  INVX1 U1223 ( .A(n4742), .Y(n3998) );
  INVX1 U1224 ( .A(\data_in<0> ), .Y(n4003) );
  INVX1 U1225 ( .A(n4741), .Y(n4001) );
  INVX1 U1226 ( .A(\data_in<1> ), .Y(n4006) );
  INVX1 U1227 ( .A(n4740), .Y(n4004) );
  INVX1 U1228 ( .A(\data_in<2> ), .Y(n4009) );
  INVX1 U1229 ( .A(n4739), .Y(n4007) );
  INVX1 U1230 ( .A(\data_in<3> ), .Y(n4012) );
  INVX1 U1231 ( .A(n4738), .Y(n4010) );
  INVX1 U1232 ( .A(\data_in<4> ), .Y(n4015) );
  INVX1 U1233 ( .A(n4737), .Y(n4013) );
  INVX1 U1234 ( .A(\data_in<5> ), .Y(n4018) );
  INVX1 U1235 ( .A(n4736), .Y(n4016) );
  INVX1 U1236 ( .A(\data_in<6> ), .Y(n4021) );
  INVX1 U1237 ( .A(n4735), .Y(n4019) );
  INVX1 U1238 ( .A(\data_in<7> ), .Y(n4024) );
  INVX1 U1239 ( .A(n4734), .Y(n4022) );
  INVX1 U1240 ( .A(\data_in<0> ), .Y(n4028) );
  INVX1 U1241 ( .A(n4733), .Y(n4026) );
  INVX1 U1242 ( .A(\data_in<1> ), .Y(n4031) );
  INVX1 U1243 ( .A(n4732), .Y(n4029) );
  INVX1 U1244 ( .A(\data_in<2> ), .Y(n4034) );
  INVX1 U1245 ( .A(n4731), .Y(n4032) );
  INVX1 U1246 ( .A(\data_in<3> ), .Y(n4037) );
  INVX1 U1247 ( .A(n4730), .Y(n4035) );
  INVX1 U1248 ( .A(\data_in<4> ), .Y(n4040) );
  INVX1 U1249 ( .A(n4729), .Y(n4038) );
  INVX1 U1250 ( .A(\data_in<5> ), .Y(n4043) );
  INVX1 U1251 ( .A(n4728), .Y(n4041) );
  INVX1 U1252 ( .A(\data_in<6> ), .Y(n4046) );
  INVX1 U1253 ( .A(n4727), .Y(n4044) );
  INVX1 U1254 ( .A(\data_in<7> ), .Y(n4049) );
  INVX1 U1255 ( .A(n4726), .Y(n4047) );
  INVX1 U1256 ( .A(\data_in<0> ), .Y(n4053) );
  INVX1 U1257 ( .A(n4725), .Y(n4051) );
  INVX1 U1258 ( .A(\data_in<1> ), .Y(n4056) );
  INVX1 U1259 ( .A(n4724), .Y(n4054) );
  INVX1 U1260 ( .A(\data_in<2> ), .Y(n4059) );
  INVX1 U1261 ( .A(n4723), .Y(n4057) );
  INVX1 U1262 ( .A(\data_in<3> ), .Y(n4062) );
  INVX1 U1263 ( .A(n4722), .Y(n4060) );
  INVX1 U1264 ( .A(\data_in<4> ), .Y(n4065) );
  INVX1 U1265 ( .A(n4721), .Y(n4063) );
  INVX1 U1266 ( .A(\data_in<5> ), .Y(n4068) );
  INVX1 U1267 ( .A(n4720), .Y(n4066) );
  INVX1 U1268 ( .A(\data_in<6> ), .Y(n4071) );
  INVX1 U1269 ( .A(n4719), .Y(n4069) );
  INVX1 U1270 ( .A(\data_in<7> ), .Y(n4074) );
  INVX1 U1271 ( .A(n4718), .Y(n4072) );
  INVX1 U1272 ( .A(\data_in<0> ), .Y(n4078) );
  INVX1 U1273 ( .A(n4717), .Y(n4076) );
  INVX1 U1274 ( .A(\data_in<1> ), .Y(n4081) );
  INVX1 U1275 ( .A(n4716), .Y(n4079) );
  INVX1 U1276 ( .A(\data_in<2> ), .Y(n4084) );
  INVX1 U1277 ( .A(n4715), .Y(n4082) );
  INVX1 U1278 ( .A(\data_in<3> ), .Y(n4087) );
  INVX1 U1279 ( .A(n4714), .Y(n4085) );
  INVX1 U1280 ( .A(\data_in<4> ), .Y(n4090) );
  INVX1 U1281 ( .A(n4713), .Y(n4088) );
  INVX1 U1282 ( .A(\data_in<5> ), .Y(n4093) );
  INVX1 U1283 ( .A(n4712), .Y(n4091) );
  INVX1 U1284 ( .A(\data_in<6> ), .Y(n4096) );
  INVX1 U1285 ( .A(n4711), .Y(n4094) );
  INVX1 U1286 ( .A(\data_in<7> ), .Y(n4099) );
  INVX1 U1287 ( .A(n4710), .Y(n4097) );
  INVX1 U1288 ( .A(\data_in<0> ), .Y(n4102) );
  INVX1 U1289 ( .A(n4709), .Y(n4100) );
  INVX1 U1290 ( .A(\data_in<1> ), .Y(n4105) );
  INVX1 U1291 ( .A(n4708), .Y(n4103) );
  INVX1 U1292 ( .A(\data_in<2> ), .Y(n4108) );
  INVX1 U1293 ( .A(n4707), .Y(n4106) );
  INVX1 U1294 ( .A(\data_in<3> ), .Y(n4111) );
  INVX1 U1295 ( .A(n4706), .Y(n4109) );
  INVX1 U1296 ( .A(\data_in<4> ), .Y(n4114) );
  INVX1 U1297 ( .A(n4705), .Y(n4112) );
  INVX1 U1298 ( .A(\data_in<5> ), .Y(n4117) );
  INVX1 U1299 ( .A(n4704), .Y(n4115) );
  INVX1 U1300 ( .A(\data_in<6> ), .Y(n4120) );
  INVX1 U1301 ( .A(n4703), .Y(n4118) );
  INVX1 U1302 ( .A(\data_in<7> ), .Y(n4123) );
  INVX1 U1303 ( .A(n4702), .Y(n4121) );
  INVX1 U1304 ( .A(\data_in<0> ), .Y(n4126) );
  INVX1 U1305 ( .A(n4701), .Y(n4124) );
  INVX1 U1306 ( .A(\data_in<1> ), .Y(n4129) );
  INVX1 U1307 ( .A(n4700), .Y(n4127) );
  INVX1 U1308 ( .A(\data_in<2> ), .Y(n4132) );
  INVX1 U1309 ( .A(n4699), .Y(n4130) );
  INVX1 U1310 ( .A(\data_in<3> ), .Y(n4135) );
  INVX1 U1311 ( .A(n4698), .Y(n4133) );
  INVX1 U1312 ( .A(\data_in<4> ), .Y(n4138) );
  INVX1 U1313 ( .A(n4697), .Y(n4136) );
  INVX1 U1314 ( .A(\data_in<5> ), .Y(n4141) );
  INVX1 U1315 ( .A(n4696), .Y(n4139) );
  INVX1 U1316 ( .A(\data_in<6> ), .Y(n4144) );
  INVX1 U1317 ( .A(n4695), .Y(n4142) );
  INVX1 U1318 ( .A(\data_in<7> ), .Y(n4147) );
  INVX1 U1319 ( .A(n4694), .Y(n4145) );
  INVX1 U1320 ( .A(\data_in<0> ), .Y(n4152) );
  INVX1 U1321 ( .A(n4693), .Y(n4150) );
  INVX1 U1322 ( .A(\data_in<1> ), .Y(n4155) );
  INVX1 U1323 ( .A(n4692), .Y(n4153) );
  INVX1 U1324 ( .A(\data_in<2> ), .Y(n4158) );
  INVX1 U1325 ( .A(n4691), .Y(n4156) );
  INVX1 U1326 ( .A(\data_in<3> ), .Y(n4161) );
  INVX1 U1327 ( .A(n4690), .Y(n4159) );
  INVX1 U1328 ( .A(\data_in<4> ), .Y(n4164) );
  INVX1 U1329 ( .A(n4689), .Y(n4162) );
  INVX1 U1330 ( .A(\data_in<5> ), .Y(n4167) );
  INVX1 U1331 ( .A(n4688), .Y(n4165) );
  INVX1 U1332 ( .A(\data_in<6> ), .Y(n4170) );
  INVX1 U1333 ( .A(n4687), .Y(n4168) );
  INVX1 U1334 ( .A(\data_in<7> ), .Y(n4173) );
  INVX1 U1335 ( .A(n4686), .Y(n4171) );
  INVX1 U1336 ( .A(\data_in<0> ), .Y(n4176) );
  INVX1 U1337 ( .A(n4685), .Y(n4174) );
  INVX1 U1338 ( .A(\data_in<1> ), .Y(n4179) );
  INVX1 U1339 ( .A(n4684), .Y(n4177) );
  INVX1 U1340 ( .A(\data_in<2> ), .Y(n4182) );
  INVX1 U1341 ( .A(n4683), .Y(n4180) );
  INVX1 U1342 ( .A(\data_in<3> ), .Y(n4185) );
  INVX1 U1343 ( .A(n4682), .Y(n4183) );
  INVX1 U1344 ( .A(\data_in<4> ), .Y(n4188) );
  INVX1 U1345 ( .A(n4681), .Y(n4186) );
  INVX1 U1346 ( .A(\data_in<5> ), .Y(n4191) );
  INVX1 U1347 ( .A(n4680), .Y(n4189) );
  INVX1 U1348 ( .A(\data_in<6> ), .Y(n4194) );
  INVX1 U1349 ( .A(n4679), .Y(n4192) );
  INVX1 U1350 ( .A(\data_in<7> ), .Y(n4197) );
  INVX1 U1351 ( .A(n4678), .Y(n4195) );
  INVX1 U1352 ( .A(\data_in<0> ), .Y(n4202) );
  INVX1 U1353 ( .A(n4677), .Y(n4200) );
  INVX1 U1354 ( .A(\data_in<1> ), .Y(n4205) );
  INVX1 U1355 ( .A(n4676), .Y(n4203) );
  INVX1 U1356 ( .A(\data_in<2> ), .Y(n4208) );
  INVX1 U1357 ( .A(n4675), .Y(n4206) );
  INVX1 U1358 ( .A(\data_in<3> ), .Y(n4211) );
  INVX1 U1359 ( .A(n4674), .Y(n4209) );
  INVX1 U1360 ( .A(\data_in<4> ), .Y(n4214) );
  INVX1 U1361 ( .A(n4673), .Y(n4212) );
  INVX1 U1362 ( .A(\data_in<5> ), .Y(n4217) );
  INVX1 U1363 ( .A(n4672), .Y(n4215) );
  INVX1 U1364 ( .A(\data_in<6> ), .Y(n4220) );
  INVX1 U1365 ( .A(n4671), .Y(n4218) );
  INVX1 U1366 ( .A(\data_in<7> ), .Y(n4223) );
  INVX1 U1367 ( .A(n4670), .Y(n4221) );
  INVX1 U1368 ( .A(\data_in<0> ), .Y(n4226) );
  INVX1 U1369 ( .A(n4669), .Y(n4224) );
  INVX1 U1370 ( .A(\data_in<1> ), .Y(n4229) );
  INVX1 U1371 ( .A(n4668), .Y(n4227) );
  INVX1 U1372 ( .A(\data_in<2> ), .Y(n4232) );
  INVX1 U1373 ( .A(n4667), .Y(n4230) );
  INVX1 U1374 ( .A(\data_in<3> ), .Y(n4235) );
  INVX1 U1375 ( .A(n4666), .Y(n4233) );
  INVX1 U1376 ( .A(\data_in<4> ), .Y(n4238) );
  INVX1 U1377 ( .A(n4665), .Y(n4236) );
  INVX1 U1378 ( .A(\data_in<5> ), .Y(n4241) );
  INVX1 U1379 ( .A(n4664), .Y(n4239) );
  INVX1 U1380 ( .A(\data_in<6> ), .Y(n4244) );
  INVX1 U1381 ( .A(n4663), .Y(n4242) );
  INVX1 U1382 ( .A(\data_in<7> ), .Y(n4247) );
  INVX1 U1383 ( .A(n4662), .Y(n4245) );
  INVX1 U1384 ( .A(\data_in<0> ), .Y(n4250) );
  INVX1 U1385 ( .A(n4661), .Y(n4248) );
  INVX1 U1386 ( .A(\data_in<1> ), .Y(n4253) );
  INVX1 U1387 ( .A(n4660), .Y(n4251) );
  INVX1 U1388 ( .A(\data_in<2> ), .Y(n4256) );
  INVX1 U1389 ( .A(n4659), .Y(n4254) );
  INVX1 U1390 ( .A(\data_in<3> ), .Y(n4259) );
  INVX1 U1391 ( .A(n4658), .Y(n4257) );
  INVX1 U1392 ( .A(\data_in<4> ), .Y(n4262) );
  INVX1 U1393 ( .A(n4657), .Y(n4260) );
  INVX1 U1394 ( .A(\data_in<5> ), .Y(n4265) );
  INVX1 U1395 ( .A(n4656), .Y(n4263) );
  INVX1 U1396 ( .A(\data_in<6> ), .Y(n4268) );
  INVX1 U1397 ( .A(n4655), .Y(n4266) );
  INVX1 U1398 ( .A(\data_in<7> ), .Y(n4271) );
  INVX1 U1399 ( .A(n4654), .Y(n4269) );
  INVX1 U1400 ( .A(\data_in<0> ), .Y(n4275) );
  INVX1 U1401 ( .A(n4653), .Y(n4273) );
  INVX1 U1402 ( .A(\data_in<1> ), .Y(n4278) );
  INVX1 U1403 ( .A(n4652), .Y(n4276) );
  INVX1 U1404 ( .A(\data_in<2> ), .Y(n4281) );
  INVX1 U1405 ( .A(n4651), .Y(n4279) );
  INVX1 U1406 ( .A(\data_in<3> ), .Y(n4284) );
  INVX1 U1407 ( .A(n4650), .Y(n4282) );
  INVX1 U1408 ( .A(\data_in<4> ), .Y(n4287) );
  INVX1 U1409 ( .A(n4649), .Y(n4285) );
  INVX1 U1410 ( .A(\data_in<5> ), .Y(n4290) );
  INVX1 U1411 ( .A(n4648), .Y(n4288) );
  INVX1 U1412 ( .A(\data_in<6> ), .Y(n4293) );
  INVX1 U1413 ( .A(n4647), .Y(n4291) );
  INVX1 U1414 ( .A(\data_in<7> ), .Y(n4296) );
  INVX1 U1415 ( .A(n4646), .Y(n4294) );
  INVX1 U1416 ( .A(\data_in<0> ), .Y(n4300) );
  INVX1 U1417 ( .A(n4645), .Y(n4298) );
  INVX1 U1418 ( .A(\data_in<1> ), .Y(n4303) );
  INVX1 U1419 ( .A(n4644), .Y(n4301) );
  INVX1 U1420 ( .A(\data_in<2> ), .Y(n4306) );
  INVX1 U1421 ( .A(n4643), .Y(n4304) );
  INVX1 U1422 ( .A(\data_in<3> ), .Y(n4309) );
  INVX1 U1423 ( .A(n4642), .Y(n4307) );
  INVX1 U1424 ( .A(\data_in<4> ), .Y(n4312) );
  INVX1 U1425 ( .A(n4641), .Y(n4310) );
  INVX1 U1426 ( .A(\data_in<5> ), .Y(n4315) );
  INVX1 U1427 ( .A(n4640), .Y(n4313) );
  INVX1 U1428 ( .A(\data_in<6> ), .Y(n4318) );
  INVX1 U1429 ( .A(n4639), .Y(n4316) );
  INVX1 U1430 ( .A(\data_in<7> ), .Y(n4321) );
  INVX1 U1431 ( .A(n4638), .Y(n4319) );
  INVX1 U1432 ( .A(\data_in<0> ), .Y(n4324) );
  INVX1 U1433 ( .A(n4637), .Y(n4322) );
  INVX1 U1434 ( .A(\data_in<1> ), .Y(n4327) );
  INVX1 U1435 ( .A(n4636), .Y(n4325) );
  INVX1 U1436 ( .A(\data_in<2> ), .Y(n4330) );
  INVX1 U1437 ( .A(n4635), .Y(n4328) );
  INVX1 U1438 ( .A(\data_in<3> ), .Y(n4333) );
  INVX1 U1439 ( .A(n4634), .Y(n4331) );
  INVX1 U1440 ( .A(\data_in<4> ), .Y(n4336) );
  INVX1 U1441 ( .A(n4633), .Y(n4334) );
  INVX1 U1442 ( .A(\data_in<5> ), .Y(n4339) );
  INVX1 U1443 ( .A(n4632), .Y(n4337) );
  INVX1 U1444 ( .A(\data_in<6> ), .Y(n4342) );
  INVX1 U1445 ( .A(n4631), .Y(n4340) );
  INVX1 U1446 ( .A(\data_in<7> ), .Y(n4345) );
  INVX1 U1447 ( .A(n4630), .Y(n4343) );
  INVX1 U1448 ( .A(\data_in<0> ), .Y(n4349) );
  INVX1 U1449 ( .A(n4629), .Y(n4347) );
  INVX1 U1450 ( .A(\data_in<1> ), .Y(n4352) );
  INVX1 U1451 ( .A(n4628), .Y(n4350) );
  INVX1 U1452 ( .A(\data_in<2> ), .Y(n4355) );
  INVX1 U1453 ( .A(n4627), .Y(n4353) );
  INVX1 U1454 ( .A(\data_in<3> ), .Y(n4358) );
  INVX1 U1455 ( .A(n4626), .Y(n4356) );
  INVX1 U1456 ( .A(\data_in<4> ), .Y(n4361) );
  INVX1 U1457 ( .A(n4625), .Y(n4359) );
  INVX1 U1458 ( .A(\data_in<5> ), .Y(n4364) );
  INVX1 U1459 ( .A(n4624), .Y(n4362) );
  INVX1 U1460 ( .A(\data_in<6> ), .Y(n4367) );
  INVX1 U1461 ( .A(n4623), .Y(n4365) );
  INVX1 U1462 ( .A(\data_in<7> ), .Y(n4370) );
  INVX1 U1463 ( .A(n4622), .Y(n4368) );
  INVX1 U1464 ( .A(\data_in<0> ), .Y(n4374) );
  INVX1 U1465 ( .A(n4621), .Y(n4372) );
  INVX1 U1466 ( .A(\data_in<1> ), .Y(n4377) );
  INVX1 U1467 ( .A(n4620), .Y(n4375) );
  INVX1 U1468 ( .A(\data_in<2> ), .Y(n4380) );
  INVX1 U1469 ( .A(n4619), .Y(n4378) );
  INVX1 U1470 ( .A(\data_in<3> ), .Y(n4383) );
  INVX1 U1471 ( .A(n4618), .Y(n4381) );
  INVX1 U1472 ( .A(\data_in<4> ), .Y(n4386) );
  INVX1 U1473 ( .A(n4617), .Y(n4384) );
  INVX1 U1474 ( .A(\data_in<5> ), .Y(n4389) );
  INVX1 U1475 ( .A(n4616), .Y(n4387) );
  INVX1 U1476 ( .A(\data_in<6> ), .Y(n4392) );
  INVX1 U1477 ( .A(n4615), .Y(n4390) );
  INVX1 U1478 ( .A(\data_in<7> ), .Y(n4395) );
  INVX1 U1479 ( .A(n4614), .Y(n4393) );
  INVX1 U1480 ( .A(\data_in<0> ), .Y(n4399) );
  INVX1 U1481 ( .A(n4613), .Y(n4397) );
  INVX1 U1482 ( .A(\data_in<1> ), .Y(n4402) );
  INVX1 U1483 ( .A(n4612), .Y(n4400) );
  INVX1 U1484 ( .A(\data_in<2> ), .Y(n4405) );
  INVX1 U1485 ( .A(n4611), .Y(n4403) );
  INVX1 U1486 ( .A(\data_in<3> ), .Y(n4408) );
  INVX1 U1487 ( .A(n4610), .Y(n4406) );
  INVX1 U1488 ( .A(\data_in<4> ), .Y(n4411) );
  INVX1 U1489 ( .A(n4609), .Y(n4409) );
  INVX1 U1490 ( .A(\data_in<5> ), .Y(n4414) );
  INVX1 U1491 ( .A(n4608), .Y(n4412) );
  INVX1 U1492 ( .A(\data_in<6> ), .Y(n4417) );
  INVX1 U1493 ( .A(n4607), .Y(n4415) );
  INVX1 U1494 ( .A(\data_in<7> ), .Y(n4420) );
  INVX1 U1495 ( .A(n4606), .Y(n4418) );
  INVX1 U1496 ( .A(\data_in<0> ), .Y(n4423) );
  INVX1 U1497 ( .A(n4605), .Y(n4421) );
  INVX1 U1498 ( .A(\data_in<1> ), .Y(n4426) );
  INVX1 U1499 ( .A(n4604), .Y(n4424) );
  INVX1 U1500 ( .A(\data_in<2> ), .Y(n4429) );
  INVX1 U1501 ( .A(n4603), .Y(n4427) );
  INVX1 U1502 ( .A(\data_in<3> ), .Y(n4432) );
  INVX1 U1503 ( .A(n4602), .Y(n4430) );
  INVX1 U1504 ( .A(\data_in<4> ), .Y(n4435) );
  INVX1 U1505 ( .A(n4601), .Y(n4433) );
  INVX1 U1506 ( .A(\data_in<5> ), .Y(n4438) );
  INVX1 U1507 ( .A(n4600), .Y(n4436) );
  INVX1 U1508 ( .A(\data_in<6> ), .Y(n4441) );
  INVX1 U1509 ( .A(n4599), .Y(n4439) );
  INVX1 U1510 ( .A(\data_in<7> ), .Y(n4444) );
  INVX1 U1511 ( .A(n4598), .Y(n4442) );
  INVX1 U1512 ( .A(\data_in<0> ), .Y(n4448) );
  INVX1 U1513 ( .A(n4597), .Y(n4446) );
  INVX1 U1514 ( .A(\data_in<1> ), .Y(n4451) );
  INVX1 U1515 ( .A(n4596), .Y(n4449) );
  INVX1 U1516 ( .A(\data_in<2> ), .Y(n4454) );
  INVX1 U1517 ( .A(n4595), .Y(n4452) );
  INVX1 U1518 ( .A(\data_in<3> ), .Y(n4457) );
  INVX1 U1519 ( .A(n4594), .Y(n4455) );
  INVX1 U1520 ( .A(\data_in<4> ), .Y(n4460) );
  INVX1 U1521 ( .A(n4593), .Y(n4458) );
  INVX1 U1522 ( .A(\data_in<5> ), .Y(n4463) );
  INVX1 U1523 ( .A(n4592), .Y(n4461) );
  INVX1 U1524 ( .A(\data_in<6> ), .Y(n4466) );
  INVX1 U1525 ( .A(n4591), .Y(n4464) );
  INVX1 U1526 ( .A(\data_in<7> ), .Y(n4469) );
  INVX1 U1527 ( .A(n4590), .Y(n4467) );
  INVX1 U1528 ( .A(\data_in<0> ), .Y(n4474) );
  INVX1 U1529 ( .A(n4589), .Y(n4472) );
  INVX1 U1530 ( .A(\data_in<1> ), .Y(n4477) );
  INVX1 U1531 ( .A(n4588), .Y(n4475) );
  INVX1 U1532 ( .A(\data_in<2> ), .Y(n4480) );
  INVX1 U1533 ( .A(n4587), .Y(n4478) );
  INVX1 U1534 ( .A(\data_in<3> ), .Y(n4483) );
  INVX1 U1535 ( .A(n4586), .Y(n4481) );
  INVX1 U1536 ( .A(\data_in<4> ), .Y(n4486) );
  INVX1 U1537 ( .A(n4585), .Y(n4484) );
  INVX1 U1538 ( .A(\data_in<5> ), .Y(n4489) );
  INVX1 U1539 ( .A(n4584), .Y(n4487) );
  INVX1 U1540 ( .A(\data_in<6> ), .Y(n4492) );
  INVX1 U1541 ( .A(n4583), .Y(n4490) );
  INVX1 U1542 ( .A(\data_in<7> ), .Y(n4495) );
  INVX1 U1543 ( .A(n4582), .Y(n4493) );
  INVX1 U1544 ( .A(\data_in<0> ), .Y(n4499) );
  INVX1 U1545 ( .A(n4581), .Y(n4497) );
  INVX1 U1546 ( .A(\data_in<1> ), .Y(n4502) );
  INVX1 U1547 ( .A(n4580), .Y(n4500) );
  INVX1 U1548 ( .A(\data_in<2> ), .Y(n4505) );
  INVX1 U1549 ( .A(n4579), .Y(n4503) );
  INVX1 U1550 ( .A(\data_in<3> ), .Y(n4508) );
  INVX1 U1551 ( .A(n4578), .Y(n4506) );
  INVX1 U1552 ( .A(\data_in<4> ), .Y(n4511) );
  INVX1 U1553 ( .A(n4577), .Y(n4509) );
  INVX1 U1554 ( .A(\data_in<5> ), .Y(n4514) );
  INVX1 U1555 ( .A(n4576), .Y(n4512) );
  INVX1 U1556 ( .A(\data_in<6> ), .Y(n4517) );
  INVX1 U1557 ( .A(n4575), .Y(n4515) );
  INVX1 U1558 ( .A(\data_in<7> ), .Y(n4520) );
  INVX1 U1559 ( .A(n4574), .Y(n4518) );
  INVX1 U1560 ( .A(\data_in<0> ), .Y(n4524) );
  INVX1 U1561 ( .A(\data_in<1> ), .Y(n4527) );
  INVX1 U1562 ( .A(\data_in<2> ), .Y(n4530) );
  INVX1 U1563 ( .A(\data_in<3> ), .Y(n4533) );
  INVX1 U1564 ( .A(\data_in<4> ), .Y(n4536) );
  INVX1 U1565 ( .A(\data_in<5> ), .Y(n4539) );
  INVX1 U1566 ( .A(\data_in<6> ), .Y(n4542) );
  INVX1 U1567 ( .A(\data_in<7> ), .Y(n4546) );
  INVX1 U1568 ( .A(\data_in<8> ), .Y(n4547) );
  INVX1 U1569 ( .A(\mem<0><0> ), .Y(n4565) );
  INVX1 U1570 ( .A(\data_in<9> ), .Y(n4548) );
  INVX1 U1571 ( .A(\mem<0><1> ), .Y(n4564) );
  INVX1 U1572 ( .A(\data_in<10> ), .Y(n4549) );
  INVX1 U1573 ( .A(\data_in<11> ), .Y(n4550) );
  INVX1 U1574 ( .A(\data_in<12> ), .Y(n4551) );
  INVX1 U1575 ( .A(\data_in<13> ), .Y(n4552) );
  INVX1 U1576 ( .A(\data_in<14> ), .Y(n4553) );
  INVX1 U1577 ( .A(\data_in<15> ), .Y(n4554) );
  INVX8 U1578 ( .A(n1534), .Y(n1548) );
  INVX8 U1579 ( .A(n1574), .Y(n1570) );
  INVX1 U1580 ( .A(N177), .Y(n1432) );
  INVX1 U1581 ( .A(n1570), .Y(n812) );
  INVX4 U1582 ( .A(n1570), .Y(n1427) );
  INVX1 U1583 ( .A(n1570), .Y(n1437) );
  INVX4 U1584 ( .A(n1552), .Y(n1564) );
  AND2X1 U1585 ( .A(n1528), .B(n897), .Y(n1208) );
  INVX1 U1586 ( .A(n1556), .Y(n58) );
  AND2X2 U1587 ( .A(n2973), .B(n1575), .Y(n28) );
  AND2X2 U1588 ( .A(n1575), .B(n2832), .Y(n29) );
  AND2X2 U1589 ( .A(n1525), .B(n1576), .Y(n30) );
  AND2X2 U1590 ( .A(n1414), .B(n1424), .Y(n31) );
  INVX1 U1591 ( .A(n1559), .Y(n1430) );
  AND2X1 U1592 ( .A(n693), .B(n1236), .Y(n1145) );
  AND2X1 U1593 ( .A(n1529), .B(n933), .Y(n1244) );
  AND2X1 U1594 ( .A(n1528), .B(n893), .Y(n1204) );
  AND2X1 U1595 ( .A(n1529), .B(n917), .Y(n1228) );
  AND2X1 U1596 ( .A(n1529), .B(n939), .Y(n1250) );
  AND2X1 U1597 ( .A(n1528), .B(n947), .Y(n1258) );
  INVX1 U1598 ( .A(\mem<41><0> ), .Y(n4863) );
  INVX1 U1599 ( .A(n4496), .Y(n1531) );
  INVX1 U1600 ( .A(\mem<31><1> ), .Y(n4783) );
  INVX1 U1601 ( .A(\mem<29><1> ), .Y(n4774) );
  INVX1 U1602 ( .A(n4496), .Y(n1532) );
  INVX1 U1603 ( .A(\mem<60><4> ), .Y(n1798) );
  INVX1 U1604 ( .A(\mem<58><6> ), .Y(n2406) );
  INVX1 U1605 ( .A(\mem<57><4> ), .Y(n1804) );
  INVX1 U1606 ( .A(\mem<28><4> ), .Y(n1813) );
  INVX1 U1607 ( .A(\mem<26><5> ), .Y(n2377) );
  INVX1 U1608 ( .A(\mem<26><7> ), .Y(n2468) );
  INVX1 U1609 ( .A(\mem<62><0> ), .Y(n1621) );
  INVX1 U1610 ( .A(\mem<62><1> ), .Y(n1679) );
  INVX1 U1611 ( .A(\mem<62><2> ), .Y(n1709) );
  INVX1 U1612 ( .A(\mem<62><3> ), .Y(n1753) );
  INVX1 U1613 ( .A(\mem<62><4> ), .Y(n1800) );
  INVX1 U1614 ( .A(\mem<62><6> ), .Y(n2402) );
  INVX1 U1615 ( .A(\mem<62><7> ), .Y(n2448) );
  INVX1 U1616 ( .A(\mem<60><0> ), .Y(n1618) );
  INVX1 U1617 ( .A(\mem<60><1> ), .Y(n1677) );
  INVX1 U1618 ( .A(\mem<60><2> ), .Y(n1708) );
  INVX1 U1619 ( .A(\mem<60><3> ), .Y(n1752) );
  INVX1 U1620 ( .A(\mem<60><5> ), .Y(n2356) );
  INVX1 U1621 ( .A(\mem<60><6> ), .Y(n2401) );
  INVX1 U1622 ( .A(\mem<58><0> ), .Y(n1608) );
  INVX1 U1623 ( .A(\mem<58><2> ), .Y(n1713) );
  INVX1 U1624 ( .A(\mem<58><3> ), .Y(n1758) );
  INVX1 U1625 ( .A(\mem<58><4> ), .Y(n1806) );
  INVX1 U1626 ( .A(\mem<58><5> ), .Y(n2362) );
  INVX1 U1627 ( .A(\mem<58><7> ), .Y(n2453) );
  INVX1 U1628 ( .A(\mem<57><7> ), .Y(n2451) );
  INVX1 U1629 ( .A(\mem<30><2> ), .Y(n1723) );
  INVX1 U1630 ( .A(\mem<30><3> ), .Y(n1768) );
  INVX1 U1631 ( .A(\mem<30><4> ), .Y(n1815) );
  INVX1 U1632 ( .A(\mem<28><2> ), .Y(n1721) );
  INVX1 U1633 ( .A(\mem<28><3> ), .Y(n1766) );
  INVX1 U1634 ( .A(\mem<28><5> ), .Y(n2370) );
  INVX1 U1635 ( .A(\mem<28><6> ), .Y(n2414) );
  INVX1 U1636 ( .A(\mem<26><2> ), .Y(n1727) );
  INVX1 U1637 ( .A(\mem<26><3> ), .Y(n1772) );
  INVX1 U1638 ( .A(\mem<25><6> ), .Y(n2419) );
  INVX1 U1639 ( .A(\mem<25><7> ), .Y(n2466) );
  INVX1 U1640 ( .A(\mem<0><6> ), .Y(n4559) );
  INVX1 U1641 ( .A(\mem<0><7> ), .Y(n4558) );
  INVX1 U1642 ( .A(\mem<0><5> ), .Y(n4560) );
  INVX1 U1643 ( .A(\mem<0><2> ), .Y(n4563) );
  INVX1 U1644 ( .A(\mem<0><3> ), .Y(n4562) );
  INVX1 U1645 ( .A(\mem<0><4> ), .Y(n4561) );
  INVX1 U1646 ( .A(\mem<62><5> ), .Y(n2357) );
  INVX1 U1647 ( .A(\mem<60><7> ), .Y(n2446) );
  INVX1 U1648 ( .A(\mem<57><0> ), .Y(n1605) );
  INVX1 U1649 ( .A(\mem<57><2> ), .Y(n1712) );
  INVX1 U1650 ( .A(\mem<57><3> ), .Y(n1757) );
  INVX1 U1651 ( .A(\mem<57><5> ), .Y(n2361) );
  INVX1 U1652 ( .A(\mem<57><6> ), .Y(n2405) );
  INVX1 U1653 ( .A(\mem<31><0> ), .Y(n1641) );
  INVX1 U1654 ( .A(\mem<30><6> ), .Y(n2416) );
  INVX1 U1655 ( .A(\mem<30><7> ), .Y(n2463) );
  INVX1 U1656 ( .A(\mem<29><0> ), .Y(n1639) );
  INVX1 U1657 ( .A(\mem<27><0> ), .Y(n1631) );
  INVX1 U1658 ( .A(\mem<27><1> ), .Y(n1684) );
  INVX1 U1659 ( .A(\mem<26><4> ), .Y(n2331) );
  INVX1 U1660 ( .A(\mem<26><6> ), .Y(n2421) );
  INVX1 U1661 ( .A(\mem<25><0> ), .Y(n1630) );
  INVX1 U1662 ( .A(\mem<25><2> ), .Y(n1726) );
  INVX1 U1663 ( .A(\mem<25><3> ), .Y(n1771) );
  INVX1 U1664 ( .A(\mem<25><5> ), .Y(n2375) );
  INVX1 U1665 ( .A(\mem<30><5> ), .Y(n2372) );
  INVX1 U1666 ( .A(\mem<28><7> ), .Y(n2461) );
  INVX1 U1667 ( .A(\mem<25><4> ), .Y(n2330) );
  INVX1 U1668 ( .A(n41), .Y(n32) );
  INVX2 U1669 ( .A(n1534), .Y(n826) );
  INVX1 U1670 ( .A(n1557), .Y(n1421) );
  MUX2X1 U1671 ( .B(\mem<51><4> ), .A(\mem<50><4> ), .S(n1550), .Y(n2778) );
  MUX2X1 U1672 ( .B(n2778), .A(n2779), .S(n1566), .Y(n2780) );
  INVX4 U1673 ( .A(n1566), .Y(n1558) );
  INVX1 U1674 ( .A(n41), .Y(n1538) );
  MUX2X1 U1675 ( .B(n2758), .A(n2757), .S(n1570), .Y(n2759) );
  INVX4 U1676 ( .A(n1549), .Y(n1537) );
  MUX2X1 U1677 ( .B(\mem<58><4> ), .A(\mem<59><4> ), .S(n1534), .Y(n2791) );
  MUX2X1 U1678 ( .B(\mem<56><4> ), .A(\mem<57><4> ), .S(n1534), .Y(n2792) );
  INVX1 U1679 ( .A(n1485), .Y(n1493) );
  MUX2X1 U1680 ( .B(\mem<45><7> ), .A(\mem<44><7> ), .S(n1489), .Y(n2970) );
  INVX4 U1681 ( .A(n1550), .Y(n33) );
  INVX1 U1682 ( .A(n626), .Y(n34) );
  INVX4 U1683 ( .A(N179), .Y(n1573) );
  INVX4 U1684 ( .A(n1573), .Y(n1572) );
  MUX2X1 U1685 ( .B(\mem<29><4> ), .A(\mem<28><4> ), .S(n1490), .Y(n2742) );
  BUFX4 U1686 ( .A(n700), .Y(n35) );
  MUX2X1 U1687 ( .B(\mem<62><4> ), .A(\mem<63><4> ), .S(n39), .Y(n2795) );
  INVX1 U1688 ( .A(n652), .Y(n36) );
  OR2X2 U1689 ( .A(n1643), .B(n1642), .Y(n560) );
  INVX1 U1690 ( .A(n588), .Y(n37) );
  INVX4 U1691 ( .A(n1424), .Y(n1578) );
  MUX2X1 U1692 ( .B(\mem<19><5> ), .A(\mem<18><5> ), .S(n41), .Y(n2823) );
  INVX1 U1693 ( .A(n1533), .Y(n38) );
  INVX1 U1694 ( .A(n1533), .Y(n1483) );
  MUX2X1 U1695 ( .B(\mem<56><5> ), .A(\mem<57><5> ), .S(n1475), .Y(n2835) );
  MUX2X1 U1696 ( .B(n2795), .A(n2796), .S(n1525), .Y(n2797) );
  MUX2X1 U1697 ( .B(\mem<44><5> ), .A(\mem<45><5> ), .S(n1539), .Y(n2850) );
  INVX1 U1698 ( .A(n1483), .Y(n39) );
  INVX1 U1699 ( .A(n39), .Y(n40) );
  MUX2X1 U1700 ( .B(\mem<49><4> ), .A(\mem<48><4> ), .S(n1548), .Y(n2779) );
  MUX2X1 U1701 ( .B(\mem<52><7> ), .A(\mem<53><7> ), .S(n1475), .Y(n2964) );
  MUX2X1 U1702 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1485), .Y(n2939) );
  INVX1 U1703 ( .A(n1555), .Y(n46) );
  MUX2X1 U1704 ( .B(\mem<36><5> ), .A(\mem<37><5> ), .S(n1485), .Y(n2828) );
  INVX8 U1705 ( .A(n1489), .Y(n1485) );
  INVX1 U1706 ( .A(n47), .Y(n41) );
  INVX1 U1707 ( .A(n9), .Y(n42) );
  INVX1 U1708 ( .A(n692), .Y(n43) );
  INVX1 U1709 ( .A(n692), .Y(n1471) );
  INVX2 U1710 ( .A(n1440), .Y(n44) );
  INVX4 U1711 ( .A(n47), .Y(n1440) );
  INVX1 U1712 ( .A(n714), .Y(n45) );
  INVX4 U1713 ( .A(n664), .Y(n813) );
  MUX2X1 U1714 ( .B(n2949), .A(n2950), .S(n46), .Y(n2951) );
  INVX4 U1715 ( .A(n1573), .Y(n1571) );
  INVX2 U1716 ( .A(n1568), .Y(n1574) );
  INVX2 U1717 ( .A(n1431), .Y(n47) );
  INVX1 U1718 ( .A(n1431), .Y(n1533) );
  MUX2X1 U1719 ( .B(\mem<61><4> ), .A(\mem<60><4> ), .S(n826), .Y(n2796) );
  INVX1 U1720 ( .A(n1440), .Y(n48) );
  INVX1 U1721 ( .A(n1440), .Y(n1484) );
  INVX1 U1722 ( .A(n50), .Y(n49) );
  INVX1 U1723 ( .A(n1518), .Y(n50) );
  MUX2X1 U1724 ( .B(\mem<42><7> ), .A(\mem<43><7> ), .S(n1485), .Y(n2971) );
  INVX1 U1725 ( .A(n595), .Y(n51) );
  INVX1 U1726 ( .A(n636), .Y(n52) );
  AND2X2 U1727 ( .A(n631), .B(n629), .Y(n53) );
  INVX1 U1728 ( .A(n686), .Y(n54) );
  BUFX4 U1729 ( .A(n700), .Y(n55) );
  AND2X2 U1730 ( .A(n624), .B(n521), .Y(n56) );
  INVX1 U1731 ( .A(n26), .Y(n693) );
  INVX2 U1732 ( .A(n128), .Y(n803) );
  BUFX4 U1733 ( .A(n1451), .Y(n57) );
  INVX1 U1734 ( .A(n1451), .Y(n828) );
  INVX2 U1735 ( .A(n1440), .Y(n1536) );
  MUX2X1 U1736 ( .B(n2866), .A(n2867), .S(n58), .Y(n2868) );
  AND2X2 U1737 ( .A(n92), .B(n414), .Y(n59) );
  AND2X2 U1738 ( .A(n31), .B(n1601), .Y(n60) );
  INVX1 U1739 ( .A(n1547), .Y(n1551) );
  INVX1 U1740 ( .A(n715), .Y(n61) );
  INVX1 U1741 ( .A(n61), .Y(n62) );
  INVX1 U1742 ( .A(n828), .Y(n829) );
  AND2X2 U1743 ( .A(n2968), .B(n1575), .Y(n70) );
  MUX2X1 U1744 ( .B(\mem<27><7> ), .A(\mem<26><7> ), .S(n1488), .Y(n2941) );
  MUX2X1 U1745 ( .B(\mem<48><7> ), .A(\mem<49><7> ), .S(n1534), .Y(n2967) );
  INVX4 U1746 ( .A(n1554), .Y(n1553) );
  INVX1 U1747 ( .A(n691), .Y(n63) );
  INVX1 U1748 ( .A(n722), .Y(n557) );
  AND2X2 U1749 ( .A(n1428), .B(n227), .Y(n722) );
  NOR2X1 U1750 ( .A(n64), .B(n65), .Y(n124) );
  AND2X2 U1751 ( .A(\mem<32><1> ), .B(n649), .Y(n64) );
  AND2X2 U1752 ( .A(\mem<33><1> ), .B(n1659), .Y(n65) );
  INVX1 U1753 ( .A(n88), .Y(n2955) );
  MUX2X1 U1754 ( .B(n2814), .A(n2813), .S(n1557), .Y(n2815) );
  MUX2X1 U1755 ( .B(\mem<46><7> ), .A(\mem<47><7> ), .S(n47), .Y(n2969) );
  INVX1 U1756 ( .A(n1534), .Y(n1487) );
  AND2X2 U1757 ( .A(n2829), .B(n1571), .Y(n68) );
  INVX2 U1758 ( .A(n1441), .Y(n1539) );
  AND2X1 U1759 ( .A(n2818), .B(n1575), .Y(n66) );
  AND2X2 U1760 ( .A(n2822), .B(n1570), .Y(n67) );
  AND2X2 U1761 ( .A(n2965), .B(n1571), .Y(n69) );
  AND2X2 U1762 ( .A(\mem<23><0> ), .B(n663), .Y(n71) );
  INVX1 U1763 ( .A(n71), .Y(n72) );
  AND2X2 U1764 ( .A(\mem<44><1> ), .B(n1468), .Y(n73) );
  INVX1 U1765 ( .A(n73), .Y(n74) );
  AND2X2 U1766 ( .A(\mem<30><0> ), .B(n1523), .Y(n75) );
  INVX1 U1767 ( .A(n75), .Y(n76) );
  AND2X2 U1768 ( .A(\mem<26><1> ), .B(n825), .Y(n77) );
  INVX1 U1769 ( .A(n77), .Y(n78) );
  INVX4 U1770 ( .A(n1432), .Y(n1534) );
  INVX1 U1771 ( .A(n691), .Y(n692) );
  INVX1 U1772 ( .A(n1441), .Y(n1541) );
  INVX1 U1773 ( .A(n1489), .Y(n1547) );
  MUX2X1 U1774 ( .B(n2823), .A(n2824), .S(n1566), .Y(n2825) );
  MUX2X1 U1775 ( .B(\mem<39><5> ), .A(\mem<38><5> ), .S(n1488), .Y(n2827) );
  MUX2X1 U1776 ( .B(\mem<27><5> ), .A(\mem<26><5> ), .S(n1440), .Y(n2816) );
  AND2X2 U1777 ( .A(n714), .B(n2688), .Y(n79) );
  INVX1 U1778 ( .A(n637), .Y(n1648) );
  INVX1 U1779 ( .A(n702), .Y(n1447) );
  AND2X2 U1780 ( .A(n715), .B(n1042), .Y(n80) );
  INVX2 U1781 ( .A(n689), .Y(n690) );
  INVX1 U1782 ( .A(n137), .Y(n81) );
  NOR3X1 U1783 ( .A(n561), .B(n551), .C(n488), .Y(n82) );
  AND2X2 U1784 ( .A(n710), .B(n2688), .Y(n83) );
  INVX4 U1785 ( .A(n648), .Y(n783) );
  INVX1 U1786 ( .A(n639), .Y(n84) );
  INVX1 U1787 ( .A(n639), .Y(n85) );
  INVX1 U1788 ( .A(n638), .Y(n639) );
  OR2X2 U1789 ( .A(n68), .B(n557), .Y(n117) );
  NOR3X1 U1790 ( .A(n487), .B(n550), .C(n558), .Y(n86) );
  INVX1 U1791 ( .A(n86), .Y(n1682) );
  INVX1 U1792 ( .A(n652), .Y(n1595) );
  INVX1 U1793 ( .A(n1523), .Y(n3795) );
  AND2X2 U1794 ( .A(n1043), .B(n715), .Y(n87) );
  NOR3X1 U1795 ( .A(n109), .B(n114), .C(n89), .Y(n88) );
  INVX1 U1796 ( .A(n2954), .Y(n89) );
  INVX1 U1797 ( .A(n610), .Y(n90) );
  INVX1 U1798 ( .A(n661), .Y(n1289) );
  NOR3X1 U1799 ( .A(n486), .B(n549), .C(n560), .Y(n91) );
  OR2X2 U1800 ( .A(n4863), .B(n63), .Y(n1513) );
  AND2X2 U1801 ( .A(n714), .B(n1424), .Y(n822) );
  NOR3X1 U1802 ( .A(n485), .B(n548), .C(n559), .Y(n92) );
  AND2X2 U1803 ( .A(n62), .B(n415), .Y(n93) );
  INVX1 U1804 ( .A(n1585), .Y(n94) );
  INVX1 U1805 ( .A(n94), .Y(n95) );
  INVX1 U1806 ( .A(n1516), .Y(n1518) );
  OR2X2 U1807 ( .A(n1029), .B(n758), .Y(n96) );
  INVX1 U1808 ( .A(n96), .Y(n97) );
  OR2X2 U1809 ( .A(n387), .B(n432), .Y(n98) );
  INVX1 U1810 ( .A(n98), .Y(\data_out<14> ) );
  OR2X2 U1811 ( .A(n239), .B(n101), .Y(n100) );
  OR2X2 U1812 ( .A(n237), .B(n238), .Y(n101) );
  OR2X2 U1813 ( .A(n242), .B(n103), .Y(n102) );
  OR2X2 U1814 ( .A(n69), .B(n70), .Y(n103) );
  OR2X2 U1815 ( .A(n1280), .B(n105), .Y(n104) );
  OR2X2 U1816 ( .A(n28), .B(n287), .Y(n105) );
  OR2X2 U1817 ( .A(n67), .B(n107), .Y(n106) );
  OR2X2 U1818 ( .A(n481), .B(n482), .Y(n107) );
  OR2X2 U1819 ( .A(n481), .B(n110), .Y(n108) );
  INVX1 U1820 ( .A(n108), .Y(n109) );
  OR2X2 U1821 ( .A(n483), .B(n484), .Y(n110) );
  OR2X2 U1822 ( .A(n545), .B(n112), .Y(n111) );
  OR2X2 U1823 ( .A(n66), .B(n544), .Y(n112) );
  OR2X2 U1824 ( .A(n545), .B(n115), .Y(n113) );
  INVX1 U1825 ( .A(n113), .Y(n114) );
  OR2X2 U1826 ( .A(n546), .B(n547), .Y(n115) );
  OR2X2 U1827 ( .A(n29), .B(n117), .Y(n116) );
  OR2X2 U1828 ( .A(n229), .B(n119), .Y(n118) );
  OR2X2 U1829 ( .A(n230), .B(n228), .Y(n119) );
  OR2X2 U1830 ( .A(n617), .B(n121), .Y(n120) );
  OR2X2 U1831 ( .A(n615), .B(n616), .Y(n121) );
  OR2X2 U1832 ( .A(n620), .B(n123), .Y(n122) );
  OR2X2 U1833 ( .A(n618), .B(n619), .Y(n123) );
  INVX1 U1834 ( .A(n124), .Y(n125) );
  AND2X2 U1835 ( .A(n815), .B(n337), .Y(n126) );
  INVX1 U1836 ( .A(n126), .Y(n127) );
  AND2X2 U1837 ( .A(n1650), .B(n1417), .Y(n128) );
  AND2X2 U1838 ( .A(n341), .B(n339), .Y(n129) );
  AND2X2 U1839 ( .A(n76), .B(n741), .Y(n130) );
  AND2X2 U1840 ( .A(n1462), .B(n1463), .Y(n131) );
  AND2X2 U1841 ( .A(n1492), .B(n1491), .Y(n132) );
  AND2X2 U1842 ( .A(n1494), .B(n1495), .Y(n133) );
  AND2X2 U1843 ( .A(n1588), .B(n1589), .Y(n134) );
  AND2X2 U1844 ( .A(n1511), .B(n1510), .Y(n135) );
  AND2X2 U1845 ( .A(n1521), .B(n1520), .Y(n136) );
  AND2X2 U1846 ( .A(n1650), .B(n651), .Y(n137) );
  OR2X2 U1847 ( .A(n1624), .B(n359), .Y(n138) );
  AND2X2 U1848 ( .A(n1093), .B(n54), .Y(n139) );
  AND2X2 U1849 ( .A(n1655), .B(n1505), .Y(n140) );
  AND2X2 U1850 ( .A(n1701), .B(n1700), .Y(n141) );
  INVX1 U1851 ( .A(n141), .Y(n142) );
  AND2X2 U1852 ( .A(n1705), .B(n1704), .Y(n143) );
  INVX1 U1853 ( .A(n143), .Y(n144) );
  OR2X2 U1854 ( .A(n144), .B(n448), .Y(n145) );
  INVX1 U1855 ( .A(n145), .Y(n146) );
  OR2X2 U1856 ( .A(n1711), .B(n1710), .Y(n147) );
  INVX1 U1857 ( .A(n147), .Y(n148) );
  INVX1 U1858 ( .A(n149), .Y(n150) );
  OR2X2 U1859 ( .A(n1729), .B(n1728), .Y(n151) );
  INVX1 U1860 ( .A(n151), .Y(n152) );
  OR2X2 U1861 ( .A(n1017), .B(n1051), .Y(n153) );
  INVX1 U1862 ( .A(n153), .Y(n154) );
  AND2X2 U1863 ( .A(n1737), .B(n1736), .Y(n155) );
  INVX1 U1864 ( .A(n155), .Y(n156) );
  AND2X2 U1865 ( .A(n1749), .B(n1748), .Y(n157) );
  INVX1 U1866 ( .A(n157), .Y(n158) );
  OR2X2 U1867 ( .A(n1755), .B(n1754), .Y(n159) );
  INVX1 U1868 ( .A(n159), .Y(n160) );
  OR2X2 U1869 ( .A(n1760), .B(n1759), .Y(n161) );
  INVX1 U1870 ( .A(n161), .Y(n162) );
  OR2X2 U1871 ( .A(n1774), .B(n1773), .Y(n163) );
  INVX1 U1872 ( .A(n163), .Y(n164) );
  OR2X2 U1873 ( .A(n1021), .B(n1063), .Y(n165) );
  INVX1 U1874 ( .A(n165), .Y(n166) );
  AND2X2 U1875 ( .A(n1792), .B(n1791), .Y(n167) );
  INVX1 U1876 ( .A(n167), .Y(n168) );
  AND2X2 U1877 ( .A(n1794), .B(n1793), .Y(n169) );
  INVX1 U1878 ( .A(n169), .Y(n170) );
  AND2X2 U1879 ( .A(n1810), .B(n1809), .Y(n171) );
  INVX1 U1880 ( .A(n171), .Y(n172) );
  OR2X2 U1881 ( .A(n353), .B(n456), .Y(n173) );
  INVX1 U1882 ( .A(n173), .Y(n174) );
  OR2X2 U1883 ( .A(n2333), .B(n2332), .Y(n175) );
  INVX1 U1884 ( .A(n175), .Y(n176) );
  AND2X2 U1885 ( .A(n2341), .B(n2340), .Y(n177) );
  INVX1 U1886 ( .A(n177), .Y(n178) );
  OR2X2 U1887 ( .A(n373), .B(n460), .Y(n179) );
  INVX1 U1888 ( .A(n179), .Y(n180) );
  OR2X2 U1889 ( .A(n2359), .B(n2358), .Y(n181) );
  INVX1 U1890 ( .A(n181), .Y(n182) );
  OR2X2 U1891 ( .A(n2364), .B(n2363), .Y(n183) );
  INVX1 U1892 ( .A(n183), .Y(n184) );
  INVX1 U1893 ( .A(n185), .Y(n186) );
  OR2X2 U1894 ( .A(n1027), .B(n1073), .Y(n187) );
  INVX1 U1895 ( .A(n187), .Y(n188) );
  OR2X2 U1896 ( .A(n743), .B(n464), .Y(n189) );
  INVX1 U1897 ( .A(n189), .Y(n190) );
  OR2X2 U1898 ( .A(n375), .B(n1075), .Y(n191) );
  INVX1 U1899 ( .A(n191), .Y(n192) );
  OR2X2 U1900 ( .A(n1031), .B(n466), .Y(n193) );
  INVX1 U1901 ( .A(n193), .Y(n194) );
  AND2X2 U1902 ( .A(n192), .B(n194), .Y(n195) );
  INVX1 U1903 ( .A(n195), .Y(n196) );
  OR2X2 U1904 ( .A(n2404), .B(n2403), .Y(n197) );
  INVX1 U1906 ( .A(n197), .Y(n198) );
  INVX1 U1907 ( .A(n199), .Y(n200) );
  OR2X2 U1908 ( .A(n2423), .B(n2422), .Y(n201) );
  INVX1 U1909 ( .A(n201), .Y(n202) );
  OR2X2 U1910 ( .A(n1033), .B(n1081), .Y(n203) );
  INVX1 U1911 ( .A(n203), .Y(n204) );
  AND2X2 U1912 ( .A(n2431), .B(n2430), .Y(n205) );
  INVX1 U1913 ( .A(n205), .Y(n206) );
  OR2X2 U1914 ( .A(n348), .B(n1083), .Y(n207) );
  INVX1 U1915 ( .A(n207), .Y(n208) );
  AND2X2 U1916 ( .A(n2441), .B(n2440), .Y(n209) );
  INVX1 U1917 ( .A(n209), .Y(n210) );
  OR2X2 U1918 ( .A(n381), .B(n470), .Y(n211) );
  INVX1 U1919 ( .A(n211), .Y(n212) );
  AND2X2 U1920 ( .A(n343), .B(n212), .Y(n213) );
  INVX1 U1921 ( .A(n213), .Y(n214) );
  OR2X2 U1922 ( .A(n2450), .B(n2449), .Y(n215) );
  INVX1 U1923 ( .A(n215), .Y(n216) );
  OR2X1 U1924 ( .A(n2455), .B(n2454), .Y(n217) );
  INVX1 U1925 ( .A(n217), .Y(n218) );
  AND2X2 U1926 ( .A(n2457), .B(n2456), .Y(n219) );
  INVX1 U1927 ( .A(n219), .Y(n220) );
  OR2X2 U1928 ( .A(n2470), .B(n2469), .Y(n221) );
  INVX1 U1929 ( .A(n221), .Y(n222) );
  AND2X2 U1930 ( .A(n2479), .B(n2478), .Y(n223) );
  INVX1 U1931 ( .A(n223), .Y(n224) );
  OR2X2 U1932 ( .A(n383), .B(n472), .Y(n225) );
  INVX1 U1933 ( .A(n225), .Y(n226) );
  AND2X2 U1934 ( .A(n2688), .B(N182), .Y(n227) );
  AND2X2 U1935 ( .A(n723), .B(n2745), .Y(n228) );
  AND2X2 U1936 ( .A(n724), .B(n2752), .Y(n229) );
  AND2X2 U1937 ( .A(n722), .B(n2759), .Y(n230) );
  AND2X2 U1938 ( .A(n1578), .B(n2767), .Y(n231) );
  OR2X2 U1939 ( .A(n2780), .B(n474), .Y(n232) );
  INVX1 U1940 ( .A(n232), .Y(n233) );
  OR2X2 U1941 ( .A(n1085), .B(n2797), .Y(n234) );
  INVX1 U1942 ( .A(n234), .Y(n235) );
  BUFX2 U1943 ( .A(n2917), .Y(n236) );
  INVX1 U1944 ( .A(n2841), .Y(n237) );
  INVX1 U1945 ( .A(n2840), .Y(n238) );
  INVX1 U1946 ( .A(n768), .Y(n239) );
  BUFX2 U1947 ( .A(n2857), .Y(n240) );
  BUFX2 U1948 ( .A(n2962), .Y(n241) );
  INVX1 U1949 ( .A(n767), .Y(n242) );
  AND2X2 U1950 ( .A(\mem<44><0> ), .B(n1468), .Y(n243) );
  INVX1 U1951 ( .A(n243), .Y(n244) );
  AND2X2 U1952 ( .A(n723), .B(n2914), .Y(n245) );
  INVX1 U1953 ( .A(n245), .Y(n246) );
  OR2X2 U1954 ( .A(n357), .B(n438), .Y(n247) );
  INVX1 U1955 ( .A(n247), .Y(n248) );
  INVX1 U1956 ( .A(n630), .Y(n249) );
  OR2X2 U1957 ( .A(n442), .B(n365), .Y(n250) );
  INVX1 U1958 ( .A(n250), .Y(n251) );
  OR2X2 U1959 ( .A(n367), .B(n444), .Y(n252) );
  INVX1 U1960 ( .A(n252), .Y(n253) );
  OR2X2 U1961 ( .A(n142), .B(n1045), .Y(n254) );
  INVX1 U1962 ( .A(n254), .Y(n255) );
  OR2X2 U1963 ( .A(n344), .B(n156), .Y(n256) );
  INVX1 U1964 ( .A(n256), .Y(n257) );
  OR2X2 U1965 ( .A(n747), .B(n1055), .Y(n258) );
  INVX1 U1966 ( .A(n258), .Y(n259) );
  OR2X2 U1967 ( .A(n345), .B(n754), .Y(n260) );
  INVX1 U1968 ( .A(n260), .Y(n261) );
  OR2X2 U1969 ( .A(n371), .B(n168), .Y(n262) );
  INVX1 U1970 ( .A(n262), .Y(n263) );
  OR2X2 U1971 ( .A(n172), .B(n458), .Y(n264) );
  INVX1 U1972 ( .A(n264), .Y(n265) );
  OR2X2 U1973 ( .A(n346), .B(n178), .Y(n266) );
  INVX1 U1974 ( .A(n266), .Y(n267) );
  OR2X2 U1975 ( .A(n749), .B(n1067), .Y(n268) );
  INVX1 U1976 ( .A(n268), .Y(n269) );
  OR2X2 U1977 ( .A(n347), .B(n756), .Y(n270) );
  INVX1 U1978 ( .A(n270), .Y(n271) );
  OR2X2 U1979 ( .A(n349), .B(n206), .Y(n272) );
  INVX1 U1980 ( .A(n272), .Y(n273) );
  OR2X2 U1981 ( .A(n350), .B(n224), .Y(n274) );
  INVX1 U1982 ( .A(n274), .Y(n275) );
  AND2X2 U1983 ( .A(n725), .B(n2766), .Y(n276) );
  INVX1 U1984 ( .A(n276), .Y(n277) );
  AND2X2 U1985 ( .A(n725), .B(n2806), .Y(n278) );
  INVX1 U1986 ( .A(n278), .Y(n279) );
  OR2X2 U1987 ( .A(n351), .B(n476), .Y(n280) );
  INVX1 U1988 ( .A(n280), .Y(n281) );
  AND2X2 U1989 ( .A(n725), .B(n2925), .Y(n282) );
  INVX1 U1990 ( .A(n282), .Y(n283) );
  OR2X2 U1991 ( .A(n389), .B(n2955), .Y(n284) );
  INVX1 U1992 ( .A(n284), .Y(n285) );
  BUFX2 U1993 ( .A(n2856), .Y(n286) );
  INVX1 U1994 ( .A(n2974), .Y(n287) );
  AND2X2 U1995 ( .A(n722), .B(n2915), .Y(n288) );
  INVX1 U1996 ( .A(n288), .Y(n289) );
  OR2X2 U1997 ( .A(n355), .B(n436), .Y(n290) );
  INVX1 U1998 ( .A(n290), .Y(n291) );
  OR2X2 U1999 ( .A(n363), .B(n434), .Y(n292) );
  INVX1 U2000 ( .A(n292), .Y(n293) );
  OR2X2 U2001 ( .A(n446), .B(n369), .Y(n294) );
  INVX1 U2002 ( .A(n294), .Y(n295) );
  OR2X2 U2003 ( .A(n745), .B(n450), .Y(n296) );
  INVX1 U2004 ( .A(n296), .Y(n297) );
  OR2X2 U2005 ( .A(n1057), .B(n158), .Y(n298) );
  INVX1 U2006 ( .A(n298), .Y(n299) );
  OR2X2 U2007 ( .A(n1023), .B(n452), .Y(n300) );
  INVX1 U2008 ( .A(n300), .Y(n301) );
  OR2X2 U2009 ( .A(n170), .B(n454), .Y(n302) );
  INVX1 U2010 ( .A(n302), .Y(n303) );
  OR2X2 U2011 ( .A(n1025), .B(n462), .Y(n304) );
  INVX1 U2012 ( .A(n304), .Y(n305) );
  OR2X2 U2013 ( .A(n377), .B(n468), .Y(n306) );
  INVX1 U2014 ( .A(n306), .Y(n307) );
  AND2X2 U2015 ( .A(n231), .B(n2774), .Y(n308) );
  INVX1 U2016 ( .A(n308), .Y(n309) );
  AND2X2 U2017 ( .A(n231), .B(n2812), .Y(n310) );
  INVX1 U2018 ( .A(n310), .Y(n311) );
  OR2X2 U2019 ( .A(n385), .B(n478), .Y(n312) );
  INVX1 U2020 ( .A(n312), .Y(n313) );
  AND2X2 U2021 ( .A(n231), .B(n2932), .Y(n314) );
  INVX1 U2022 ( .A(n314), .Y(n315) );
  OR2X2 U2023 ( .A(n391), .B(n480), .Y(n316) );
  INVX1 U2024 ( .A(n316), .Y(n317) );
  AND2X2 U2025 ( .A(\mem<26><0> ), .B(n825), .Y(n318) );
  INVX1 U2026 ( .A(n318), .Y(n319) );
  AND2X2 U2027 ( .A(\mem<56><2> ), .B(n793), .Y(n320) );
  INVX1 U2028 ( .A(n320), .Y(n321) );
  AND2X2 U2029 ( .A(\mem<27><2> ), .B(n3899), .Y(n322) );
  INVX1 U2030 ( .A(n322), .Y(n323) );
  AND2X2 U2031 ( .A(\mem<27><3> ), .B(n3899), .Y(n324) );
  INVX1 U2032 ( .A(n324), .Y(n325) );
  AND2X2 U2033 ( .A(\mem<27><4> ), .B(n3899), .Y(n326) );
  INVX1 U2034 ( .A(n326), .Y(n327) );
  AND2X2 U2035 ( .A(\mem<56><6> ), .B(n793), .Y(n328) );
  INVX1 U2036 ( .A(n328), .Y(n329) );
  AND2X2 U2037 ( .A(\mem<61><7> ), .B(n662), .Y(n330) );
  INVX1 U2038 ( .A(n330), .Y(n331) );
  AND2X2 U2039 ( .A(\mem<56><7> ), .B(n793), .Y(n332) );
  INVX1 U2040 ( .A(n332), .Y(n333) );
  AND2X2 U2041 ( .A(\mem<29><7> ), .B(n798), .Y(n334) );
  INVX1 U2042 ( .A(n334), .Y(n335) );
  AND2X2 U2043 ( .A(n2783), .B(n1558), .Y(n336) );
  INVX1 U2044 ( .A(n336), .Y(n337) );
  OR2X2 U2045 ( .A(n1808), .B(n1807), .Y(n338) );
  INVX1 U2046 ( .A(n338), .Y(n339) );
  OR2X2 U2047 ( .A(n1802), .B(n1801), .Y(n340) );
  INVX1 U2048 ( .A(n340), .Y(n341) );
  OR2X2 U2049 ( .A(n379), .B(n210), .Y(n342) );
  INVX1 U2050 ( .A(n342), .Y(n343) );
  BUFX2 U2051 ( .A(n1738), .Y(n344) );
  BUFX2 U2052 ( .A(n1783), .Y(n345) );
  BUFX2 U2053 ( .A(n2342), .Y(n346) );
  BUFX2 U2054 ( .A(n2387), .Y(n347) );
  BUFX2 U2055 ( .A(n2437), .Y(n348) );
  BUFX2 U2056 ( .A(n2432), .Y(n349) );
  BUFX2 U2057 ( .A(n2480), .Y(n350) );
  BUFX2 U2058 ( .A(n2833), .Y(n351) );
  AND2X2 U2059 ( .A(n265), .B(n129), .Y(n352) );
  INVX1 U2060 ( .A(n352), .Y(n353) );
  AND2X2 U2061 ( .A(n134), .B(n1587), .Y(n354) );
  INVX1 U2062 ( .A(n354), .Y(n355) );
  AND2X2 U2063 ( .A(n1597), .B(n1596), .Y(n356) );
  INVX1 U2064 ( .A(n356), .Y(n357) );
  AND2X2 U2065 ( .A(\addr<12> ), .B(\addr<13> ), .Y(n358) );
  INVX1 U2066 ( .A(n358), .Y(n359) );
  AND2X2 U2067 ( .A(n1645), .B(n1644), .Y(n360) );
  AND2X2 U2068 ( .A(n1652), .B(n1653), .Y(n361) );
  AND2X2 U2069 ( .A(n1661), .B(n1662), .Y(n362) );
  INVX1 U2070 ( .A(n362), .Y(n363) );
  AND2X2 U2071 ( .A(n1664), .B(n1663), .Y(n364) );
  INVX1 U2072 ( .A(n364), .Y(n365) );
  AND2X2 U2073 ( .A(n1695), .B(n1694), .Y(n366) );
  INVX1 U2074 ( .A(n366), .Y(n367) );
  AND2X2 U2075 ( .A(n1698), .B(n1699), .Y(n368) );
  INVX1 U2076 ( .A(n368), .Y(n369) );
  AND2X2 U2077 ( .A(n1790), .B(n1789), .Y(n370) );
  INVX1 U2078 ( .A(n370), .Y(n371) );
  AND2X2 U2079 ( .A(n2344), .B(n2343), .Y(n372) );
  INVX1 U2080 ( .A(n372), .Y(n373) );
  AND2X2 U2081 ( .A(n2394), .B(n2393), .Y(n374) );
  INVX1 U2082 ( .A(n374), .Y(n375) );
  AND2X2 U2083 ( .A(n2434), .B(n2433), .Y(n376) );
  INVX1 U2084 ( .A(n376), .Y(n377) );
  AND2X2 U2085 ( .A(n2439), .B(n2438), .Y(n378) );
  INVX1 U2086 ( .A(n378), .Y(n379) );
  AND2X2 U2087 ( .A(n2443), .B(n2442), .Y(n380) );
  INVX1 U2088 ( .A(n380), .Y(n381) );
  AND2X2 U2089 ( .A(n2482), .B(n2481), .Y(n382) );
  INVX1 U2090 ( .A(n382), .Y(n383) );
  AND2X2 U2091 ( .A(n100), .B(n1172), .Y(n384) );
  INVX1 U2092 ( .A(n384), .Y(n385) );
  AND2X2 U2093 ( .A(n236), .B(n2916), .Y(n386) );
  INVX1 U2094 ( .A(n386), .Y(n387) );
  AND2X2 U2095 ( .A(n283), .B(n315), .Y(n388) );
  INVX1 U2096 ( .A(n388), .Y(n389) );
  AND2X2 U2097 ( .A(n241), .B(n1172), .Y(n390) );
  INVX1 U2098 ( .A(n390), .Y(n391) );
  BUFX2 U2099 ( .A(n1690), .Y(n392) );
  BUFX2 U2100 ( .A(n1788), .Y(n393) );
  AND2X2 U2101 ( .A(n1636), .B(n130), .Y(n394) );
  INVX1 U2102 ( .A(n394), .Y(n395) );
  AND2X2 U2103 ( .A(n1480), .B(n78), .Y(n396) );
  INVX1 U2104 ( .A(n396), .Y(n397) );
  AND2X2 U2105 ( .A(n1613), .B(n1612), .Y(n398) );
  INVX1 U2106 ( .A(n398), .Y(n399) );
  AND2X2 U2107 ( .A(n12), .B(n17), .Y(n400) );
  AND2X2 U2108 ( .A(n293), .B(n251), .Y(n401) );
  INVX1 U2109 ( .A(n401), .Y(n402) );
  AND2X2 U2110 ( .A(n1675), .B(n1674), .Y(n403) );
  INVX1 U2111 ( .A(n403), .Y(n404) );
  AND2X2 U2112 ( .A(n295), .B(n253), .Y(n405) );
  AND2X2 U2113 ( .A(n2335), .B(n2334), .Y(n406) );
  INVX1 U2114 ( .A(n406), .Y(n407) );
  AND2X2 U2115 ( .A(n2472), .B(n2471), .Y(n408) );
  INVX1 U2116 ( .A(n408), .Y(n409) );
  AND2X2 U2117 ( .A(n819), .B(n1691), .Y(n410) );
  INVX1 U2118 ( .A(n410), .Y(n411) );
  AND2X2 U2119 ( .A(n1614), .B(n1615), .Y(n412) );
  INVX1 U2120 ( .A(n412), .Y(n413) );
  AND2X2 U2121 ( .A(N181), .B(n1634), .Y(n415) );
  AND2X2 U2122 ( .A(n1637), .B(n1638), .Y(n416) );
  INVX1 U2123 ( .A(n416), .Y(n417) );
  AND2X2 U2124 ( .A(n1672), .B(n1673), .Y(n418) );
  INVX1 U2125 ( .A(n418), .Y(n419) );
  AND2X2 U2126 ( .A(n1689), .B(n1688), .Y(n420) );
  INVX1 U2127 ( .A(n420), .Y(n421) );
  AND2X2 U2128 ( .A(n2337), .B(n2336), .Y(n422) );
  INVX1 U2129 ( .A(n422), .Y(n423) );
  INVX1 U2130 ( .A(n424), .Y(n425) );
  AND2X2 U2131 ( .A(n2459), .B(n2458), .Y(n426) );
  INVX1 U2132 ( .A(n426), .Y(n427) );
  AND2X2 U2133 ( .A(n2474), .B(n2473), .Y(n428) );
  INVX1 U2134 ( .A(n428), .Y(n429) );
  INVX1 U2135 ( .A(n430), .Y(n431) );
  BUFX2 U2136 ( .A(n2918), .Y(n432) );
  AND2X2 U2137 ( .A(n1660), .B(n752), .Y(n433) );
  INVX1 U2138 ( .A(n433), .Y(n434) );
  AND2X2 U2139 ( .A(n1594), .B(n1593), .Y(n435) );
  INVX1 U2140 ( .A(n435), .Y(n436) );
  AND2X2 U2141 ( .A(n1599), .B(n1598), .Y(n437) );
  INVX1 U2142 ( .A(n437), .Y(n438) );
  AND2X2 U2143 ( .A(n1646), .B(n1647), .Y(n439) );
  AND2X2 U2144 ( .A(n1656), .B(n1657), .Y(n440) );
  AND2X2 U2145 ( .A(n1666), .B(n1665), .Y(n441) );
  INVX1 U2146 ( .A(n441), .Y(n442) );
  AND2X2 U2147 ( .A(n1692), .B(n1693), .Y(n443) );
  INVX1 U2148 ( .A(n443), .Y(n444) );
  AND2X2 U2149 ( .A(n1697), .B(n1696), .Y(n445) );
  INVX1 U2150 ( .A(n445), .Y(n446) );
  AND2X2 U2151 ( .A(n1707), .B(n1706), .Y(n447) );
  INVX1 U2152 ( .A(n447), .Y(n448) );
  AND2X2 U2153 ( .A(n1742), .B(n1741), .Y(n449) );
  INVX1 U2154 ( .A(n449), .Y(n450) );
  AND2X2 U2155 ( .A(n1787), .B(n1786), .Y(n451) );
  INVX1 U2156 ( .A(n451), .Y(n452) );
  AND2X2 U2157 ( .A(n1796), .B(n1795), .Y(n453) );
  INVX1 U2158 ( .A(n453), .Y(n454) );
  AND2X2 U2159 ( .A(n263), .B(n303), .Y(n455) );
  INVX1 U2160 ( .A(n455), .Y(n456) );
  AND2X2 U2161 ( .A(n1812), .B(n1811), .Y(n457) );
  INVX1 U2162 ( .A(n457), .Y(n458) );
  AND2X2 U2163 ( .A(n2346), .B(n2345), .Y(n459) );
  INVX1 U2164 ( .A(n459), .Y(n460) );
  AND2X2 U2165 ( .A(n2355), .B(n2354), .Y(n461) );
  INVX1 U2166 ( .A(n461), .Y(n462) );
  INVX1 U2167 ( .A(n463), .Y(n464) );
  AND2X2 U2168 ( .A(n2400), .B(n2399), .Y(n465) );
  INVX1 U2169 ( .A(n465), .Y(n466) );
  AND2X2 U2170 ( .A(n2436), .B(n2435), .Y(n467) );
  INVX1 U2171 ( .A(n467), .Y(n468) );
  AND2X2 U2172 ( .A(n2445), .B(n2444), .Y(n469) );
  INVX1 U2173 ( .A(n469), .Y(n470) );
  AND2X2 U2174 ( .A(n2484), .B(n2483), .Y(n471) );
  INVX1 U2175 ( .A(n471), .Y(n472) );
  AND2X2 U2176 ( .A(n1575), .B(n767), .Y(n473) );
  INVX1 U2177 ( .A(n473), .Y(n474) );
  AND2X2 U2178 ( .A(n279), .B(n311), .Y(n475) );
  INVX1 U2179 ( .A(n475), .Y(n476) );
  AND2X2 U2180 ( .A(n240), .B(n286), .Y(n477) );
  INVX1 U2181 ( .A(n477), .Y(n478) );
  AND2X2 U2182 ( .A(n102), .B(n104), .Y(n479) );
  INVX1 U2183 ( .A(n479), .Y(n480) );
  INVX1 U2184 ( .A(n724), .Y(n481) );
  INVX1 U2185 ( .A(n2826), .Y(n482) );
  INVX1 U2186 ( .A(n2953), .Y(n483) );
  INVX1 U2187 ( .A(n2952), .Y(n484) );
  OR2X2 U2188 ( .A(n1633), .B(n1632), .Y(n486) );
  OR2X2 U2189 ( .A(n1671), .B(n1670), .Y(n487) );
  OR2X2 U2190 ( .A(n1686), .B(n1685), .Y(n488) );
  AND2X2 U2191 ( .A(\mem<30><1> ), .B(n1523), .Y(n489) );
  INVX1 U2192 ( .A(n489), .Y(n490) );
  OR2X2 U2193 ( .A(n1725), .B(n1724), .Y(n491) );
  INVX1 U2194 ( .A(n491), .Y(n492) );
  OR2X2 U2195 ( .A(n1061), .B(n1059), .Y(n493) );
  INVX1 U2196 ( .A(n493), .Y(n494) );
  INVX1 U2197 ( .A(n495), .Y(n496) );
  INVX1 U2198 ( .A(n497), .Y(n498) );
  INVX1 U2199 ( .A(n499), .Y(n500) );
  OR2X2 U2200 ( .A(n1079), .B(n1077), .Y(n501) );
  INVX1 U2201 ( .A(n501), .Y(n502) );
  OR2X1 U2202 ( .A(n2418), .B(n2417), .Y(n503) );
  INVX1 U2203 ( .A(n503), .Y(n504) );
  OR2X2 U2204 ( .A(n2465), .B(n2464), .Y(n505) );
  INVX1 U2205 ( .A(n505), .Y(n506) );
  AND2X2 U2206 ( .A(n2844), .B(n1571), .Y(n507) );
  INVX1 U2207 ( .A(n507), .Y(n508) );
  AND2X2 U2208 ( .A(n1571), .B(n2851), .Y(n509) );
  INVX1 U2209 ( .A(n509), .Y(n510) );
  BUFX2 U2210 ( .A(n1586), .Y(n511) );
  INVX1 U2211 ( .A(n511), .Y(n512) );
  INVX1 U2212 ( .A(n511), .Y(n513) );
  BUFX2 U2213 ( .A(n1590), .Y(n514) );
  INVX1 U2214 ( .A(n514), .Y(n515) );
  INVX1 U2215 ( .A(n514), .Y(n516) );
  INVX1 U2216 ( .A(n514), .Y(n517) );
  BUFX2 U2217 ( .A(n1592), .Y(n518) );
  INVX1 U2218 ( .A(n518), .Y(n519) );
  INVX1 U2219 ( .A(n518), .Y(n520) );
  INVX1 U2220 ( .A(n518), .Y(n521) );
  AND2X2 U2221 ( .A(n512), .B(n1616), .Y(n522) );
  OR2X2 U2222 ( .A(n1007), .B(n1053), .Y(n523) );
  INVX1 U2223 ( .A(n523), .Y(n524) );
  OR2X2 U2224 ( .A(n393), .B(n1065), .Y(n525) );
  INVX1 U2225 ( .A(n525), .Y(n526) );
  OR2X2 U2226 ( .A(n1009), .B(n425), .Y(n527) );
  INVX1 U2227 ( .A(n527), .Y(n528) );
  OR2X2 U2228 ( .A(n1011), .B(n431), .Y(n529) );
  INVX1 U2229 ( .A(n529), .Y(n530) );
  OR2X2 U2230 ( .A(n402), .B(n1682), .Y(n531) );
  INVX1 U2231 ( .A(n531), .Y(n532) );
  OR2X2 U2232 ( .A(n1015), .B(n1035), .Y(n533) );
  INVX1 U2233 ( .A(n533), .Y(n534) );
  OR2X2 U2234 ( .A(n1019), .B(n1037), .Y(n535) );
  INVX1 U2235 ( .A(n535), .Y(n536) );
  OR2X2 U2236 ( .A(n751), .B(n1039), .Y(n537) );
  INVX1 U2237 ( .A(n537), .Y(n538) );
  OR2X2 U2238 ( .A(n196), .B(n1041), .Y(n539) );
  INVX1 U2239 ( .A(n539), .Y(n540) );
  OR2X2 U2240 ( .A(n214), .B(n857), .Y(n541) );
  INVX1 U2241 ( .A(n541), .Y(n542) );
  BUFX2 U2242 ( .A(n2887), .Y(n543) );
  INVX1 U2243 ( .A(n2819), .Y(n544) );
  INVX1 U2244 ( .A(n723), .Y(n545) );
  INVX1 U2245 ( .A(n2945), .Y(n546) );
  INVX1 U2246 ( .A(n2944), .Y(n547) );
  OR2X2 U2247 ( .A(n399), .B(n413), .Y(n548) );
  OR2X2 U2248 ( .A(n395), .B(n417), .Y(n549) );
  OR2X2 U2249 ( .A(n1681), .B(n1680), .Y(n550) );
  OR2X2 U2250 ( .A(n392), .B(n421), .Y(n551) );
  AND2X2 U2251 ( .A(n2937), .B(n1575), .Y(n552) );
  INVX1 U2252 ( .A(n552), .Y(n553) );
  AND2X2 U2253 ( .A(n2961), .B(n1575), .Y(n554) );
  INVX1 U2254 ( .A(n554), .Y(n555) );
  BUFX2 U2255 ( .A(n2886), .Y(n556) );
  OR2X2 U2256 ( .A(n419), .B(n404), .Y(n558) );
  OR2X2 U2257 ( .A(n1623), .B(n1622), .Y(n559) );
  OR2X2 U2258 ( .A(n397), .B(n411), .Y(n561) );
  OR2X2 U2259 ( .A(n1049), .B(n1047), .Y(n562) );
  INVX1 U2260 ( .A(n562), .Y(n563) );
  OR2X2 U2261 ( .A(n407), .B(n423), .Y(n564) );
  INVX1 U2262 ( .A(n564), .Y(n565) );
  OR2X2 U2263 ( .A(n1071), .B(n1069), .Y(n566) );
  INVX1 U2264 ( .A(n566), .Y(n567) );
  OR2X2 U2265 ( .A(n220), .B(n427), .Y(n568) );
  INVX1 U2266 ( .A(n568), .Y(n569) );
  OR2X2 U2267 ( .A(n409), .B(n429), .Y(n570) );
  INVX1 U2268 ( .A(n570), .Y(n571) );
  AND2X2 U2269 ( .A(n1423), .B(n136), .Y(n572) );
  INVX1 U2270 ( .A(n572), .Y(n573) );
  AND2X2 U2271 ( .A(n2958), .B(n1423), .Y(n574) );
  INVX1 U2272 ( .A(n574), .Y(n575) );
  AND2X2 U2273 ( .A(n2738), .B(n2737), .Y(n576) );
  INVX1 U2274 ( .A(n576), .Y(n577) );
  AND2X2 U2275 ( .A(n2722), .B(n2721), .Y(n578) );
  INVX1 U2276 ( .A(n578), .Y(n579) );
  AND2X2 U2277 ( .A(n277), .B(n309), .Y(n580) );
  INVX1 U2278 ( .A(n580), .Y(n581) );
  OR2X2 U2279 ( .A(n2794), .B(n2793), .Y(n582) );
  INVX1 U2280 ( .A(n582), .Y(n583) );
  AND2X2 U2281 ( .A(n1443), .B(n1611), .Y(n584) );
  INVX1 U2282 ( .A(n584), .Y(n585) );
  INVX1 U2283 ( .A(n584), .Y(n586) );
  AND2X2 U2284 ( .A(n83), .B(n87), .Y(n587) );
  INVX1 U2285 ( .A(n587), .Y(n588) );
  INVX1 U2286 ( .A(n587), .Y(n589) );
  AND2X2 U2287 ( .A(n861), .B(n1606), .Y(n590) );
  INVX1 U2288 ( .A(n590), .Y(n591) );
  INVX1 U2289 ( .A(n590), .Y(n592) );
  AND2X2 U2290 ( .A(n4), .B(n774), .Y(n593) );
  INVX1 U2291 ( .A(n593), .Y(n594) );
  INVX1 U2292 ( .A(n593), .Y(n595) );
  AND2X2 U2293 ( .A(n712), .B(n1093), .Y(n596) );
  INVX1 U2294 ( .A(n596), .Y(n597) );
  INVX1 U2295 ( .A(n596), .Y(n598) );
  AND2X2 U2296 ( .A(n1508), .B(n774), .Y(n600) );
  INVX1 U2297 ( .A(n600), .Y(n601) );
  AND2X2 U2298 ( .A(n1649), .B(n34), .Y(n609) );
  INVX1 U2299 ( .A(n609), .Y(n610) );
  INVX1 U2300 ( .A(n609), .Y(n611) );
  AND2X2 U2301 ( .A(n521), .B(n15), .Y(n612) );
  INVX1 U2302 ( .A(n612), .Y(n613) );
  INVX1 U2303 ( .A(n612), .Y(n614) );
  INVX1 U2304 ( .A(n2704), .Y(n615) );
  INVX1 U2305 ( .A(n2703), .Y(n616) );
  INVX1 U2306 ( .A(n2705), .Y(n617) );
  INVX1 U2307 ( .A(n2798), .Y(n618) );
  INVX1 U2308 ( .A(n2800), .Y(n619) );
  INVX1 U2309 ( .A(n2799), .Y(n620) );
  OR2X2 U2310 ( .A(n717), .B(n1013), .Y(n621) );
  INVX1 U2311 ( .A(n621), .Y(n622) );
  INVX1 U2312 ( .A(n621), .Y(n623) );
  AND2X2 U2313 ( .A(n628), .B(n631), .Y(n624) );
  INVX1 U2314 ( .A(n624), .Y(n626) );
  OR2X2 U2315 ( .A(n718), .B(n1635), .Y(n627) );
  INVX1 U2316 ( .A(n627), .Y(n628) );
  INVX1 U2317 ( .A(n627), .Y(n629) );
  OR2X2 U2318 ( .A(n22), .B(N181), .Y(n630) );
  INVX1 U2319 ( .A(n630), .Y(n631) );
  INVX1 U2320 ( .A(n630), .Y(n632) );
  AND2X2 U2321 ( .A(n1438), .B(n1619), .Y(n633) );
  AND2X2 U2322 ( .A(n60), .B(n249), .Y(n635) );
  INVX1 U2323 ( .A(n635), .Y(n636) );
  INVX1 U2324 ( .A(n635), .Y(n637) );
  AND2X2 U2325 ( .A(n1595), .B(n49), .Y(n638) );
  INVX1 U2326 ( .A(n638), .Y(n640) );
  AND2X2 U2327 ( .A(n517), .B(n24), .Y(n641) );
  INVX1 U2328 ( .A(n641), .Y(n642) );
  INVX1 U2329 ( .A(n641), .Y(n643) );
  AND2X2 U2330 ( .A(n1651), .B(n519), .Y(n644) );
  INVX1 U2331 ( .A(n644), .Y(n645) );
  INVX1 U2332 ( .A(n644), .Y(n646) );
  AND2X2 U2333 ( .A(n36), .B(n517), .Y(n647) );
  INVX1 U2334 ( .A(n647), .Y(n648) );
  AND2X2 U2335 ( .A(n1649), .B(n15), .Y(n649) );
  INVX1 U2336 ( .A(n649), .Y(n650) );
  AND2X2 U2337 ( .A(n80), .B(n79), .Y(n651) );
  INVX1 U2338 ( .A(n651), .Y(n652) );
  INVX1 U2339 ( .A(n651), .Y(n653) );
  AND2X2 U2340 ( .A(n1093), .B(n1595), .Y(n654) );
  INVX1 U2341 ( .A(n654), .Y(n655) );
  AND2X2 U2342 ( .A(n519), .B(n789), .Y(n656) );
  INVX1 U2343 ( .A(n656), .Y(n657) );
  AND2X2 U2344 ( .A(n516), .B(n1611), .Y(n658) );
  INVX1 U2345 ( .A(n658), .Y(n659) );
  INVX1 U2346 ( .A(n658), .Y(n660) );
  AND2X2 U2347 ( .A(n37), .B(n520), .Y(n661) );
  AND2X2 U2348 ( .A(n519), .B(n1616), .Y(n662) );
  AND2X2 U2349 ( .A(n1651), .B(n1093), .Y(n663) );
  INVX1 U2350 ( .A(n663), .Y(n664) );
  AND2X2 U2351 ( .A(n1650), .B(n52), .Y(n665) );
  INVX1 U2352 ( .A(n665), .Y(n666) );
  AND2X2 U2353 ( .A(n516), .B(n53), .Y(n667) );
  INVX1 U2354 ( .A(n667), .Y(n668) );
  INVX1 U2355 ( .A(n667), .Y(n669) );
  AND2X2 U2356 ( .A(n512), .B(n15), .Y(n670) );
  INVX1 U2357 ( .A(n670), .Y(n671) );
  INVX1 U2358 ( .A(n670), .Y(n672) );
  AND2X2 U2359 ( .A(n36), .B(n1655), .Y(n673) );
  INVX1 U2360 ( .A(n673), .Y(n674) );
  AND2X2 U2361 ( .A(n36), .B(n513), .Y(n675) );
  INVX1 U2362 ( .A(n675), .Y(n676) );
  AND2X2 U2363 ( .A(n1650), .B(n1508), .Y(n677) );
  INVX1 U2364 ( .A(n677), .Y(n678) );
  AND2X2 U2365 ( .A(n1508), .B(n1518), .Y(n679) );
  INVX1 U2366 ( .A(n679), .Y(n680) );
  INVX1 U2367 ( .A(n679), .Y(n681) );
  AND2X2 U2368 ( .A(n1655), .B(n635), .Y(n682) );
  INVX1 U2369 ( .A(n682), .Y(n683) );
  INVX1 U2370 ( .A(n682), .Y(n684) );
  AND2X2 U2371 ( .A(n861), .B(n1515), .Y(n685) );
  INVX1 U2372 ( .A(n685), .Y(n686) );
  AND2X2 U2373 ( .A(n512), .B(n1648), .Y(n687) );
  AND2X2 U2374 ( .A(n520), .B(n23), .Y(n689) );
  AND2X2 U2375 ( .A(n1650), .B(n587), .Y(n691) );
  AND2X2 U2376 ( .A(n513), .B(n2), .Y(n694) );
  AND2X2 U2377 ( .A(n37), .B(n1093), .Y(n695) );
  AND2X2 U2378 ( .A(n712), .B(n512), .Y(n696) );
  AND2X2 U2379 ( .A(n766), .B(n520), .Y(n698) );
  AND2X2 U2380 ( .A(n1443), .B(n1508), .Y(n699) );
  AND2X2 U2381 ( .A(n1093), .B(n52), .Y(n700) );
  AND2X2 U2382 ( .A(n24), .B(n49), .Y(n701) );
  INVX1 U2383 ( .A(n701), .Y(n702) );
  INVX1 U2384 ( .A(n701), .Y(n703) );
  AND2X2 U2385 ( .A(n766), .B(n49), .Y(n704) );
  INVX1 U2386 ( .A(n704), .Y(n705) );
  INVX1 U2387 ( .A(n704), .Y(n706) );
  AND2X2 U2388 ( .A(n766), .B(n1443), .Y(n707) );
  INVX1 U2389 ( .A(n707), .Y(n708) );
  INVX1 U2390 ( .A(n707), .Y(n709) );
  AND2X2 U2391 ( .A(n1581), .B(n1582), .Y(n710) );
  INVX1 U2392 ( .A(n710), .Y(n711) );
  AND2X2 U2393 ( .A(n1603), .B(n623), .Y(n712) );
  INVX1 U2394 ( .A(n766), .Y(n713) );
  AND2X2 U2395 ( .A(n1581), .B(n1426), .Y(n714) );
  AND2X2 U2396 ( .A(n1473), .B(n1514), .Y(n715) );
  AND2X2 U2397 ( .A(n1473), .B(n1583), .Y(n716) );
  INVX1 U2398 ( .A(n716), .Y(n717) );
  INVX1 U2399 ( .A(n716), .Y(n718) );
  AND2X2 U2400 ( .A(n1649), .B(n53), .Y(n719) );
  AND2X2 U2401 ( .A(n513), .B(n1651), .Y(n720) );
  AND2X2 U2402 ( .A(n1578), .B(n227), .Y(n721) );
  AND2X2 U2403 ( .A(n1578), .B(n765), .Y(n723) );
  AND2X2 U2404 ( .A(n1579), .B(n765), .Y(n724) );
  AND2X2 U2405 ( .A(n1428), .B(n2767), .Y(n725) );
  AND2X2 U2406 ( .A(\mem<54><0> ), .B(n14), .Y(n726) );
  INVX1 U2407 ( .A(n726), .Y(n727) );
  AND2X2 U2408 ( .A(\mem<24><1> ), .B(n600), .Y(n728) );
  INVX1 U2409 ( .A(n728), .Y(n729) );
  AND2X2 U2410 ( .A(\mem<29><2> ), .B(n798), .Y(n730) );
  INVX1 U2411 ( .A(n730), .Y(n731) );
  AND2X2 U2412 ( .A(\mem<29><3> ), .B(n799), .Y(n732) );
  INVX1 U2413 ( .A(n732), .Y(n733) );
  AND2X2 U2414 ( .A(\mem<29><4> ), .B(n799), .Y(n734) );
  INVX1 U2415 ( .A(n734), .Y(n735) );
  AND2X2 U2416 ( .A(\mem<29><5> ), .B(n799), .Y(n736) );
  INVX1 U2417 ( .A(n736), .Y(n737) );
  AND2X2 U2418 ( .A(\mem<29><6> ), .B(n798), .Y(n738) );
  INVX1 U2419 ( .A(n738), .Y(n739) );
  AND2X2 U2420 ( .A(\mem<17><0> ), .B(n677), .Y(n740) );
  INVX1 U2421 ( .A(n740), .Y(n741) );
  INVX1 U2422 ( .A(n2392), .Y(n742) );
  INVX1 U2423 ( .A(n742), .Y(n743) );
  AND2X2 U2424 ( .A(n1740), .B(n1739), .Y(n744) );
  INVX1 U2425 ( .A(n744), .Y(n745) );
  AND2X2 U2426 ( .A(n1745), .B(n1744), .Y(n746) );
  INVX1 U2427 ( .A(n746), .Y(n747) );
  AND2X2 U2428 ( .A(n2349), .B(n2348), .Y(n748) );
  INVX1 U2429 ( .A(n748), .Y(n749) );
  AND2X2 U2430 ( .A(n269), .B(n305), .Y(n750) );
  INVX1 U2431 ( .A(n750), .Y(n751) );
  INVX1 U2432 ( .A(n125), .Y(n752) );
  AND2X2 U2433 ( .A(n1782), .B(n1781), .Y(n753) );
  INVX1 U2434 ( .A(n753), .Y(n754) );
  AND2X2 U2435 ( .A(n2386), .B(n2385), .Y(n755) );
  INVX1 U2436 ( .A(n755), .Y(n756) );
  AND2X2 U2437 ( .A(n2391), .B(n2390), .Y(n757) );
  INVX1 U2438 ( .A(n757), .Y(n758) );
  OR2X2 U2439 ( .A(n2475), .B(n4560), .Y(n759) );
  INVX1 U2440 ( .A(n759), .Y(n760) );
  AND2X2 U2441 ( .A(\mem<2><3> ), .B(n786), .Y(n761) );
  INVX1 U2442 ( .A(n761), .Y(n762) );
  AND2X2 U2443 ( .A(\mem<2><5> ), .B(n787), .Y(n763) );
  INVX1 U2444 ( .A(n763), .Y(n764) );
  AND2X2 U2445 ( .A(N181), .B(n1634), .Y(n765) );
  AND2X2 U2446 ( .A(n1603), .B(n622), .Y(n766) );
  AND2X2 U2447 ( .A(n1428), .B(n1429), .Y(n767) );
  AND2X2 U2448 ( .A(n1578), .B(n1429), .Y(n768) );
  AND2X2 U2449 ( .A(\mem<17><1> ), .B(n677), .Y(n769) );
  INVX1 U2450 ( .A(n769), .Y(n770) );
  INVX1 U2451 ( .A(n597), .Y(n3167) );
  AND2X2 U2452 ( .A(n766), .B(n1650), .Y(n771) );
  INVX1 U2453 ( .A(n771), .Y(n772) );
  INVX1 U2454 ( .A(n771), .Y(n773) );
  INVX1 U2455 ( .A(n2975), .Y(n774) );
  INVX2 U2456 ( .A(n2975), .Y(n1649) );
  INVX1 U2457 ( .A(n674), .Y(n775) );
  INVX1 U2458 ( .A(n674), .Y(n776) );
  INVX1 U2459 ( .A(n1264), .Y(n777) );
  INVX1 U2460 ( .A(n676), .Y(n778) );
  INVX1 U2461 ( .A(n676), .Y(n3669) );
  INVX1 U2462 ( .A(n640), .Y(n779) );
  INVX1 U2463 ( .A(n678), .Y(n780) );
  INVX1 U2464 ( .A(n678), .Y(n781) );
  INVX1 U2465 ( .A(n646), .Y(n782) );
  INVX1 U2466 ( .A(n681), .Y(n784) );
  INVX1 U2467 ( .A(n680), .Y(n785) );
  INVX1 U2468 ( .A(n681), .Y(n1467) );
  INVX1 U2469 ( .A(n684), .Y(n786) );
  INVX1 U2470 ( .A(n683), .Y(n787) );
  INVX1 U2471 ( .A(n683), .Y(n1503) );
  INVX2 U2472 ( .A(n650), .Y(n788) );
  INVX1 U2473 ( .A(n653), .Y(n789) );
  INVX1 U2474 ( .A(n589), .Y(n792) );
  INVX1 U2475 ( .A(n588), .Y(n1611) );
  INVX1 U2476 ( .A(n594), .Y(n793) );
  INVX1 U2477 ( .A(n595), .Y(n3166) );
  BUFX2 U2478 ( .A(n522), .Y(n794) );
  INVX1 U2479 ( .A(n773), .Y(n795) );
  INVX1 U2480 ( .A(n773), .Y(n796) );
  INVX1 U2481 ( .A(n772), .Y(n3324) );
  INVX1 U2482 ( .A(n613), .Y(n798) );
  INVX1 U2483 ( .A(n614), .Y(n799) );
  INVX1 U2484 ( .A(n688), .Y(n800) );
  INVX1 U2485 ( .A(n688), .Y(n4471) );
  INVX2 U2486 ( .A(n669), .Y(n801) );
  INVX1 U2487 ( .A(n668), .Y(n4199) );
  INVX1 U2488 ( .A(n128), .Y(n802) );
  INVX1 U2489 ( .A(n1283), .Y(n804) );
  INVX1 U2490 ( .A(\addr<10> ), .Y(n805) );
  INVX1 U2491 ( .A(n805), .Y(n806) );
  INVX2 U2492 ( .A(n703), .Y(n816) );
  INVX1 U2493 ( .A(n666), .Y(n807) );
  INVX1 U2494 ( .A(n809), .Y(n808) );
  INVX1 U2495 ( .A(n665), .Y(n809) );
  AND2X2 U2496 ( .A(n516), .B(n1619), .Y(n810) );
  INVX8 U2497 ( .A(n810), .Y(n2980) );
  INVX1 U2498 ( .A(n3141), .Y(n3114) );
  MUX2X1 U2499 ( .B(\mem<9><4> ), .A(\mem<8><4> ), .S(n1549), .Y(n2769) );
  INVX1 U2500 ( .A(n1534), .Y(n1474) );
  MUX2X1 U2501 ( .B(\mem<33><4> ), .A(\mem<32><4> ), .S(n1550), .Y(n2754) );
  INVX1 U2502 ( .A(n2980), .Y(n3006) );
  MUX2X1 U2503 ( .B(n2753), .A(n2754), .S(n1439), .Y(n2758) );
  INVX1 U2504 ( .A(n672), .Y(n811) );
  INVX1 U2505 ( .A(n671), .Y(n3899) );
  INVX8 U2506 ( .A(n814), .Y(n3087) );
  MUX2X1 U2507 ( .B(\mem<47><5> ), .A(\mem<46><5> ), .S(n1550), .Y(n2849) );
  MUX2X1 U2508 ( .B(n2843), .A(n2842), .S(n1556), .Y(n2844) );
  MUX2X1 U2509 ( .B(n2772), .A(n2773), .S(n812), .Y(n2774) );
  MUX2X1 U2510 ( .B(\mem<39><4> ), .A(\mem<38><4> ), .S(n1549), .Y(n2755) );
  OR2X2 U2511 ( .A(n1424), .B(N182), .Y(n1635) );
  AND2X2 U2512 ( .A(n1655), .B(n1619), .Y(n814) );
  NAND2X1 U2513 ( .A(n2784), .B(n1430), .Y(n815) );
  AND2X2 U2514 ( .A(n1785), .B(n1784), .Y(n1022) );
  MUX2X1 U2515 ( .B(n2734), .A(n2735), .S(n812), .Y(n2736) );
  INVX1 U2516 ( .A(n3087), .Y(n3113) );
  NAND2X1 U2517 ( .A(n817), .B(n818), .Y(n819) );
  INVX1 U2518 ( .A(n1285), .Y(n817) );
  INVX1 U2519 ( .A(n4783), .Y(n818) );
  INVX1 U2520 ( .A(n796), .Y(n820) );
  INVX1 U2521 ( .A(n820), .Y(n821) );
  NAND2X1 U2522 ( .A(n661), .B(\mem<45><1> ), .Y(n1470) );
  INVX2 U2523 ( .A(n643), .Y(n823) );
  INVX1 U2524 ( .A(n642), .Y(n4396) );
  MUX2X1 U2525 ( .B(\mem<59><6> ), .A(\mem<58><6> ), .S(n826), .Y(n2864) );
  INVX1 U2526 ( .A(n1522), .Y(n824) );
  AND2X2 U2527 ( .A(n1443), .B(n15), .Y(n825) );
  OR2X2 U2528 ( .A(n1092), .B(n592), .Y(n2977) );
  INVX1 U2529 ( .A(n1419), .Y(n827) );
  INVX1 U2530 ( .A(n1556), .Y(n1439) );
  MUX2X1 U2531 ( .B(\mem<1><6> ), .A(\mem<0><6> ), .S(n841), .Y(n2859) );
  BUFX2 U2532 ( .A(N181), .Y(n830) );
  INVX2 U2533 ( .A(n660), .Y(n832) );
  INVX1 U2534 ( .A(n659), .Y(n1502) );
  MUX2X1 U2535 ( .B(\mem<19><6> ), .A(\mem<18><6> ), .S(n1493), .Y(n2878) );
  INVX1 U2536 ( .A(n1468), .Y(n1465) );
  NAND2X1 U2537 ( .A(\mem<59><1> ), .B(n522), .Y(n834) );
  INVX1 U2538 ( .A(n824), .Y(n835) );
  INVX1 U2539 ( .A(n1522), .Y(n1499) );
  INVX1 U2540 ( .A(n1499), .Y(n1500) );
  INVX1 U2541 ( .A(n671), .Y(n836) );
  MUX2X1 U2542 ( .B(n2972), .A(n2971), .S(n1559), .Y(n2973) );
  NAND2X1 U2543 ( .A(\mem<45><0> ), .B(n661), .Y(n837) );
  AND2X2 U2544 ( .A(n837), .B(n244), .Y(n1598) );
  MUX2X1 U2545 ( .B(\mem<25><4> ), .A(\mem<24><4> ), .S(n40), .Y(n2740) );
  INVX1 U2546 ( .A(n1414), .Y(n838) );
  INVX1 U2547 ( .A(n709), .Y(n839) );
  INVX1 U2548 ( .A(n709), .Y(n840) );
  INVX1 U2549 ( .A(n1534), .Y(n841) );
  AND2X2 U2550 ( .A(n1438), .B(n54), .Y(n842) );
  MUX2X1 U2551 ( .B(\mem<19><4> ), .A(\mem<18><4> ), .S(n1551), .Y(n2746) );
  INVX1 U2552 ( .A(\addr<9> ), .Y(n843) );
  INVX1 U2553 ( .A(n843), .Y(n844) );
  INVX1 U2554 ( .A(n1469), .Y(n845) );
  INVX1 U2555 ( .A(n845), .Y(n846) );
  INVX2 U2556 ( .A(n845), .Y(n847) );
  INVX2 U2557 ( .A(n1549), .Y(n1454) );
  NAND2X1 U2558 ( .A(\mem<20><0> ), .B(n1467), .Y(n848) );
  AND2X2 U2559 ( .A(n72), .B(n848), .Y(n1638) );
  INVX1 U2560 ( .A(n680), .Y(n852) );
  INVX1 U2561 ( .A(n1457), .Y(n853) );
  INVX2 U2562 ( .A(n3218), .Y(n854) );
  MUX2X1 U2563 ( .B(n2739), .A(n2740), .S(n1519), .Y(n2744) );
  NAND2X1 U2564 ( .A(\mem<55><0> ), .B(n3167), .Y(n855) );
  AND2X2 U2565 ( .A(n855), .B(n727), .Y(n1615) );
  MUX2X1 U2566 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1544), .Y(n2860) );
  MUX2X1 U2567 ( .B(n2865), .A(n2864), .S(n1558), .Y(n2869) );
  INVX1 U2568 ( .A(n2460), .Y(n856) );
  INVX1 U2569 ( .A(n856), .Y(n857) );
  AND2X2 U2570 ( .A(\mem<2><2> ), .B(n787), .Y(n858) );
  INVX1 U2571 ( .A(n858), .Y(n859) );
  INVX4 U2572 ( .A(n586), .Y(n860) );
  INVX1 U2573 ( .A(rst), .Y(n1580) );
  AND2X2 U2574 ( .A(n1578), .B(N181), .Y(n861) );
  AND2X2 U2575 ( .A(n1268), .B(n3141), .Y(n862) );
  INVX1 U2576 ( .A(n862), .Y(n863) );
  AND2X2 U2577 ( .A(n3218), .B(n1422), .Y(n864) );
  INVX1 U2578 ( .A(n864), .Y(n865) );
  AND2X2 U2579 ( .A(n3218), .B(n1269), .Y(n866) );
  INVX1 U2580 ( .A(n866), .Y(n867) );
  AND2X1 U2581 ( .A(n3375), .B(n820), .Y(n868) );
  INVX1 U2582 ( .A(n868), .Y(n869) );
  AND2X1 U2583 ( .A(n3375), .B(n1267), .Y(n870) );
  INVX1 U2584 ( .A(n870), .Y(n871) );
  AND2X1 U2585 ( .A(n1286), .B(n1267), .Y(n872) );
  INVX1 U2586 ( .A(n872), .Y(n873) );
  AND2X2 U2587 ( .A(n1286), .B(n1289), .Y(n874) );
  INVX1 U2588 ( .A(n874), .Y(n875) );
  AND2X2 U2589 ( .A(n3472), .B(n1289), .Y(n876) );
  INVX1 U2590 ( .A(n876), .Y(n877) );
  AND2X1 U2591 ( .A(n3472), .B(n1266), .Y(n878) );
  INVX1 U2592 ( .A(n878), .Y(n879) );
  AND2X1 U2593 ( .A(n1260), .B(n1266), .Y(n880) );
  INVX1 U2594 ( .A(n880), .Y(n881) );
  AND2X1 U2595 ( .A(n3546), .B(n1260), .Y(n882) );
  INVX1 U2596 ( .A(n882), .Y(n883) );
  AND2X1 U2597 ( .A(n3571), .B(n3546), .Y(n884) );
  INVX1 U2598 ( .A(n884), .Y(n885) );
  AND2X1 U2599 ( .A(n3571), .B(n655), .Y(n886) );
  INVX1 U2600 ( .A(n886), .Y(n887) );
  AND2X1 U2601 ( .A(n3620), .B(n655), .Y(n888) );
  INVX1 U2602 ( .A(n888), .Y(n889) );
  AND2X1 U2603 ( .A(n3620), .B(n657), .Y(n890) );
  INVX1 U2604 ( .A(n890), .Y(n891) );
  AND2X1 U2605 ( .A(n640), .B(n657), .Y(n892) );
  INVX1 U2606 ( .A(n892), .Y(n893) );
  AND2X1 U2607 ( .A(n640), .B(n1264), .Y(n894) );
  INVX1 U2608 ( .A(n894), .Y(n895) );
  AND2X1 U2609 ( .A(n1263), .B(n1264), .Y(n896) );
  INVX1 U2610 ( .A(n896), .Y(n897) );
  AND2X2 U2611 ( .A(n1263), .B(n81), .Y(n898) );
  INVX1 U2612 ( .A(n898), .Y(n899) );
  AND2X2 U2613 ( .A(n1287), .B(n1265), .Y(n900) );
  INVX1 U2614 ( .A(n900), .Y(n901) );
  AND2X2 U2615 ( .A(n1271), .B(n803), .Y(n902) );
  INVX1 U2616 ( .A(n902), .Y(n903) );
  AND2X1 U2617 ( .A(n1272), .B(n1271), .Y(n904) );
  INVX1 U2618 ( .A(n904), .Y(n905) );
  AND2X1 U2619 ( .A(n4025), .B(n1272), .Y(n906) );
  INVX1 U2620 ( .A(n906), .Y(n907) );
  AND2X1 U2621 ( .A(n4025), .B(n4050), .Y(n908) );
  INVX1 U2622 ( .A(n908), .Y(n909) );
  AND2X1 U2623 ( .A(n4075), .B(n4050), .Y(n910) );
  INVX1 U2624 ( .A(n910), .Y(n911) );
  AND2X1 U2625 ( .A(n4075), .B(n1436), .Y(n912) );
  INVX1 U2626 ( .A(n912), .Y(n913) );
  AND2X1 U2627 ( .A(n1436), .B(n1273), .Y(n914) );
  INVX1 U2628 ( .A(n914), .Y(n915) );
  AND2X1 U2629 ( .A(n1273), .B(n4148), .Y(n916) );
  INVX1 U2630 ( .A(n916), .Y(n917) );
  AND2X1 U2631 ( .A(n1506), .B(n4148), .Y(n918) );
  INVX1 U2632 ( .A(n918), .Y(n919) );
  AND2X1 U2633 ( .A(n4198), .B(n1506), .Y(n920) );
  INVX1 U2634 ( .A(n920), .Y(n921) );
  AND2X1 U2635 ( .A(n4198), .B(n1275), .Y(n922) );
  INVX1 U2636 ( .A(n922), .Y(n923) );
  INVX1 U2637 ( .A(n924), .Y(n925) );
  INVX1 U2638 ( .A(n926), .Y(n927) );
  AND2X1 U2639 ( .A(n4272), .B(n4297), .Y(n928) );
  INVX1 U2640 ( .A(n928), .Y(n929) );
  AND2X1 U2641 ( .A(n1277), .B(n4297), .Y(n930) );
  INVX1 U2642 ( .A(n930), .Y(n931) );
  AND2X1 U2643 ( .A(n4346), .B(n1277), .Y(n932) );
  INVX1 U2644 ( .A(n932), .Y(n933) );
  AND2X1 U2645 ( .A(n4371), .B(n4346), .Y(n934) );
  INVX1 U2646 ( .A(n934), .Y(n935) );
  AND2X1 U2647 ( .A(n1276), .B(n4371), .Y(n936) );
  INVX1 U2648 ( .A(n936), .Y(n937) );
  AND2X1 U2649 ( .A(n1445), .B(n1276), .Y(n938) );
  INVX1 U2650 ( .A(n938), .Y(n939) );
  AND2X1 U2651 ( .A(n1445), .B(n4445), .Y(n940) );
  INVX1 U2652 ( .A(n940), .Y(n941) );
  AND2X1 U2653 ( .A(n4470), .B(n4445), .Y(n942) );
  INVX1 U2654 ( .A(n942), .Y(n943) );
  AND2X1 U2655 ( .A(n4470), .B(n1274), .Y(n944) );
  INVX1 U2656 ( .A(n944), .Y(n945) );
  AND2X1 U2657 ( .A(n4521), .B(n1274), .Y(n946) );
  INVX1 U2658 ( .A(n946), .Y(n947) );
  BUFX2 U2659 ( .A(n608), .Y(n948) );
  BUFX2 U2660 ( .A(n607), .Y(n949) );
  BUFX2 U2661 ( .A(n606), .Y(n950) );
  BUFX2 U2662 ( .A(n605), .Y(n951) );
  BUFX2 U2663 ( .A(n604), .Y(n952) );
  BUFX2 U2664 ( .A(n603), .Y(n953) );
  BUFX2 U2665 ( .A(n602), .Y(n954) );
  BUFX2 U2666 ( .A(n599), .Y(n955) );
  BUFX2 U2667 ( .A(n4523), .Y(n956) );
  BUFX2 U2668 ( .A(n4526), .Y(n957) );
  BUFX2 U2669 ( .A(n4529), .Y(n958) );
  BUFX2 U2670 ( .A(n4532), .Y(n959) );
  BUFX2 U2671 ( .A(n4535), .Y(n960) );
  BUFX2 U2672 ( .A(n4538), .Y(n961) );
  BUFX2 U2673 ( .A(n4541), .Y(n962) );
  BUFX2 U2674 ( .A(n4545), .Y(n963) );
  AND2X2 U2675 ( .A(\mem<0><0> ), .B(n1496), .Y(n964) );
  INVX1 U2676 ( .A(n964), .Y(n965) );
  AND2X2 U2677 ( .A(\mem<24><0> ), .B(n600), .Y(n966) );
  INVX1 U2678 ( .A(n966), .Y(n967) );
  AND2X2 U2679 ( .A(\mem<0><1> ), .B(n1496), .Y(n968) );
  INVX1 U2680 ( .A(n968), .Y(n969) );
  AND2X2 U2681 ( .A(\mem<61><2> ), .B(n662), .Y(n970) );
  INVX1 U2682 ( .A(n970), .Y(n971) );
  AND2X2 U2683 ( .A(\mem<63><2> ), .B(n2978), .Y(n972) );
  INVX1 U2684 ( .A(n972), .Y(n973) );
  AND2X2 U2685 ( .A(\mem<59><2> ), .B(n522), .Y(n974) );
  INVX1 U2686 ( .A(n974), .Y(n975) );
  AND2X2 U2687 ( .A(\mem<24><2> ), .B(n797), .Y(n976) );
  INVX1 U2688 ( .A(n976), .Y(n977) );
  AND2X2 U2689 ( .A(\mem<61><3> ), .B(n662), .Y(n978) );
  INVX1 U2690 ( .A(n978), .Y(n979) );
  AND2X2 U2691 ( .A(\mem<63><3> ), .B(n2978), .Y(n980) );
  INVX1 U2692 ( .A(n980), .Y(n981) );
  AND2X2 U2693 ( .A(\mem<59><3> ), .B(n522), .Y(n982) );
  INVX1 U2694 ( .A(n982), .Y(n983) );
  AND2X2 U2695 ( .A(\mem<24><3> ), .B(n797), .Y(n984) );
  INVX1 U2696 ( .A(n984), .Y(n985) );
  AND2X2 U2697 ( .A(\mem<24><4> ), .B(n797), .Y(n986) );
  INVX1 U2698 ( .A(n986), .Y(n987) );
  AND2X2 U2699 ( .A(\mem<61><5> ), .B(n662), .Y(n988) );
  INVX1 U2700 ( .A(n988), .Y(n989) );
  AND2X2 U2701 ( .A(\mem<63><5> ), .B(n2978), .Y(n990) );
  INVX1 U2702 ( .A(n990), .Y(n991) );
  AND2X2 U2703 ( .A(\mem<59><5> ), .B(n522), .Y(n992) );
  INVX1 U2704 ( .A(n992), .Y(n993) );
  AND2X2 U2705 ( .A(\mem<24><5> ), .B(n797), .Y(n994) );
  INVX1 U2706 ( .A(n994), .Y(n995) );
  AND2X2 U2707 ( .A(\mem<61><6> ), .B(n662), .Y(n996) );
  INVX1 U2708 ( .A(n996), .Y(n997) );
  AND2X2 U2709 ( .A(\mem<63><6> ), .B(n2978), .Y(n998) );
  INVX1 U2710 ( .A(n998), .Y(n999) );
  AND2X2 U2711 ( .A(\mem<59><6> ), .B(n522), .Y(n1000) );
  INVX1 U2712 ( .A(n1000), .Y(n1001) );
  AND2X2 U2713 ( .A(\mem<24><6> ), .B(n797), .Y(n1002) );
  INVX1 U2714 ( .A(n1002), .Y(n1003) );
  AND2X2 U2715 ( .A(\mem<24><7> ), .B(n797), .Y(n1004) );
  INVX1 U2716 ( .A(n1004), .Y(n1005) );
  INVX1 U2717 ( .A(n1743), .Y(n1006) );
  INVX1 U2718 ( .A(n1006), .Y(n1007) );
  INVX1 U2719 ( .A(n2347), .Y(n1008) );
  INVX1 U2720 ( .A(n1008), .Y(n1009) );
  INVX1 U2721 ( .A(n2485), .Y(n1010) );
  INVX1 U2722 ( .A(n1010), .Y(n1011) );
  AND2X2 U2723 ( .A(N181), .B(N182), .Y(n1012) );
  INVX1 U2724 ( .A(n1012), .Y(n1013) );
  AND2X2 U2725 ( .A(n255), .B(n146), .Y(n1014) );
  INVX1 U2726 ( .A(n1014), .Y(n1015) );
  AND2X2 U2727 ( .A(n1731), .B(n1730), .Y(n1016) );
  INVX1 U2728 ( .A(n1016), .Y(n1017) );
  AND2X2 U2729 ( .A(n259), .B(n299), .Y(n1018) );
  INVX1 U2730 ( .A(n1018), .Y(n1019) );
  AND2X2 U2731 ( .A(n1776), .B(n1775), .Y(n1020) );
  INVX1 U2732 ( .A(n1020), .Y(n1021) );
  INVX1 U2733 ( .A(n1022), .Y(n1023) );
  AND2X2 U2734 ( .A(n2353), .B(n2352), .Y(n1024) );
  INVX1 U2735 ( .A(n1024), .Y(n1025) );
  AND2X2 U2736 ( .A(n2381), .B(n2380), .Y(n1026) );
  INVX1 U2737 ( .A(n1026), .Y(n1027) );
  AND2X2 U2738 ( .A(n2389), .B(n2388), .Y(n1028) );
  INVX1 U2739 ( .A(n1028), .Y(n1029) );
  AND2X2 U2740 ( .A(n2398), .B(n2397), .Y(n1030) );
  INVX1 U2741 ( .A(n1030), .Y(n1031) );
  AND2X2 U2742 ( .A(n2425), .B(n2424), .Y(n1032) );
  INVX1 U2743 ( .A(n1032), .Y(n1033) );
  INVX1 U2744 ( .A(n1720), .Y(n1034) );
  INVX1 U2745 ( .A(n1034), .Y(n1035) );
  INVX1 U2746 ( .A(n1765), .Y(n1036) );
  INVX1 U2747 ( .A(n1036), .Y(n1037) );
  INVX1 U2748 ( .A(n2369), .Y(n1038) );
  INVX1 U2749 ( .A(n1038), .Y(n1039) );
  INVX1 U2750 ( .A(n2413), .Y(n1040) );
  INVX1 U2751 ( .A(n1040), .Y(n1041) );
  AND2X2 U2752 ( .A(n1579), .B(N182), .Y(n1042) );
  AND2X2 U2753 ( .A(n1578), .B(N182), .Y(n1043) );
  AND2X2 U2754 ( .A(n1703), .B(n1702), .Y(n1044) );
  INVX1 U2755 ( .A(n1044), .Y(n1045) );
  AND2X2 U2756 ( .A(n1717), .B(n1716), .Y(n1046) );
  INVX1 U2757 ( .A(n1046), .Y(n1047) );
  AND2X2 U2758 ( .A(n1719), .B(n1718), .Y(n1048) );
  INVX1 U2759 ( .A(n1048), .Y(n1049) );
  AND2X2 U2760 ( .A(n1733), .B(n1732), .Y(n1050) );
  INVX1 U2761 ( .A(n1050), .Y(n1051) );
  INVX1 U2762 ( .A(n1052), .Y(n1053) );
  AND2X2 U2763 ( .A(n1747), .B(n1746), .Y(n1054) );
  INVX1 U2764 ( .A(n1054), .Y(n1055) );
  AND2X2 U2765 ( .A(n1751), .B(n1750), .Y(n1056) );
  INVX1 U2766 ( .A(n1056), .Y(n1057) );
  AND2X2 U2767 ( .A(n1761), .B(n1762), .Y(n1058) );
  INVX1 U2768 ( .A(n1058), .Y(n1059) );
  AND2X2 U2769 ( .A(n1764), .B(n1763), .Y(n1060) );
  INVX1 U2770 ( .A(n1060), .Y(n1061) );
  AND2X2 U2771 ( .A(n1778), .B(n1777), .Y(n1062) );
  INVX1 U2772 ( .A(n1062), .Y(n1063) );
  INVX1 U2773 ( .A(n1064), .Y(n1065) );
  AND2X2 U2774 ( .A(n2351), .B(n2350), .Y(n1066) );
  INVX1 U2775 ( .A(n1066), .Y(n1067) );
  AND2X2 U2776 ( .A(n2366), .B(n2365), .Y(n1068) );
  INVX1 U2777 ( .A(n1068), .Y(n1069) );
  AND2X2 U2778 ( .A(n2368), .B(n2367), .Y(n1070) );
  INVX1 U2779 ( .A(n1070), .Y(n1071) );
  AND2X2 U2780 ( .A(n2383), .B(n2382), .Y(n1072) );
  INVX1 U2781 ( .A(n1072), .Y(n1073) );
  AND2X2 U2782 ( .A(n2396), .B(n2395), .Y(n1074) );
  INVX1 U2783 ( .A(n1074), .Y(n1075) );
  AND2X2 U2784 ( .A(n2410), .B(n2409), .Y(n1076) );
  INVX1 U2785 ( .A(n1076), .Y(n1077) );
  AND2X2 U2786 ( .A(n2412), .B(n2411), .Y(n1078) );
  INVX1 U2787 ( .A(n1078), .Y(n1079) );
  AND2X2 U2788 ( .A(n2427), .B(n2426), .Y(n1080) );
  INVX1 U2789 ( .A(n1080), .Y(n1081) );
  INVX1 U2790 ( .A(n1082), .Y(n1083) );
  AND2X2 U2791 ( .A(n1570), .B(n768), .Y(n1084) );
  INVX1 U2792 ( .A(n1084), .Y(n1085) );
  AND2X2 U2793 ( .A(\mem<2><4> ), .B(n786), .Y(n1086) );
  INVX1 U2794 ( .A(n1086), .Y(n1087) );
  AND2X2 U2795 ( .A(\mem<2><6> ), .B(n786), .Y(n1088) );
  INVX1 U2796 ( .A(n1088), .Y(n1089) );
  AND2X2 U2797 ( .A(\mem<2><7> ), .B(n787), .Y(n1090) );
  INVX1 U2798 ( .A(n1090), .Y(n1091) );
  INVX1 U2799 ( .A(n1654), .Y(n1092) );
  INVX2 U2800 ( .A(n1092), .Y(n1093) );
  INVX1 U2801 ( .A(n1591), .Y(n1654) );
  AND2X1 U2802 ( .A(n719), .B(n1230), .Y(n1382) );
  AND2X1 U2803 ( .A(n4555), .B(n1270), .Y(n1094) );
  AND2X2 U2804 ( .A(n2978), .B(n4555), .Y(n1095) );
  AND2X2 U2805 ( .A(n2980), .B(n2979), .Y(n1096) );
  AND2X1 U2806 ( .A(n1419), .B(n3007), .Y(n1097) );
  AND2X2 U2807 ( .A(n634), .B(n3033), .Y(n1098) );
  AND2X1 U2808 ( .A(n1425), .B(n3060), .Y(n1099) );
  AND2X2 U2809 ( .A(n3087), .B(n3086), .Y(n1100) );
  AND2X2 U2810 ( .A(n3141), .B(n3115), .Y(n1101) );
  AND2X1 U2811 ( .A(n1174), .B(n1268), .Y(n1102) );
  AND2X1 U2812 ( .A(n1422), .B(n3168), .Y(n1103) );
  AND2X2 U2813 ( .A(n3218), .B(n1176), .Y(n1104) );
  AND2X1 U2814 ( .A(n1178), .B(n1269), .Y(n1105) );
  AND2X1 U2815 ( .A(n1477), .B(n3243), .Y(n1106) );
  AND2X1 U2816 ( .A(n3270), .B(n697), .Y(n1107) );
  AND2X1 U2817 ( .A(n1476), .B(n3297), .Y(n1108) );
  AND2X1 U2818 ( .A(n3325), .B(n820), .Y(n1109) );
  AND2X1 U2819 ( .A(n3375), .B(n1180), .Y(n1110) );
  AND2X1 U2820 ( .A(n1182), .B(n1267), .Y(n1111) );
  AND2X1 U2821 ( .A(n1286), .B(n1184), .Y(n1112) );
  AND2X2 U2822 ( .A(n1289), .B(n1186), .Y(n1113) );
  AND2X1 U2823 ( .A(n3472), .B(n1188), .Y(n1114) );
  AND2X1 U2824 ( .A(n1190), .B(n1266), .Y(n1115) );
  AND2X1 U2825 ( .A(n1260), .B(n1192), .Y(n1116) );
  AND2X1 U2826 ( .A(n3546), .B(n1194), .Y(n1117) );
  AND2X1 U2827 ( .A(n3571), .B(n1196), .Y(n1118) );
  AND2X1 U2828 ( .A(n655), .B(n1198), .Y(n1119) );
  AND2X1 U2829 ( .A(n3620), .B(n1200), .Y(n1120) );
  AND2X1 U2830 ( .A(n1202), .B(n657), .Y(n1121) );
  AND2X1 U2831 ( .A(n640), .B(n1204), .Y(n1122) );
  AND2X1 U2832 ( .A(n1206), .B(n1264), .Y(n1123) );
  AND2X1 U2833 ( .A(n1263), .B(n1208), .Y(n1124) );
  AND2X2 U2834 ( .A(n1288), .B(n1210), .Y(n1125) );
  AND2X1 U2835 ( .A(n1212), .B(n1265), .Y(n1126) );
  AND2X2 U2836 ( .A(n1284), .B(n3767), .Y(n1127) );
  AND2X2 U2837 ( .A(n3795), .B(n3794), .Y(n1128) );
  AND2X2 U2838 ( .A(n3821), .B(n1283), .Y(n1129) );
  AND2X2 U2839 ( .A(n1482), .B(n3847), .Y(n1130) );
  AND2X2 U2840 ( .A(n3873), .B(n671), .Y(n1131) );
  AND2X2 U2841 ( .A(n849), .B(n3900), .Y(n1132) );
  AND2X2 U2842 ( .A(n802), .B(n3927), .Y(n1133) );
  AND2X1 U2843 ( .A(n1214), .B(n1271), .Y(n1134) );
  AND2X1 U2844 ( .A(n1272), .B(n1216), .Y(n1135) );
  AND2X1 U2845 ( .A(n4025), .B(n1218), .Y(n1136) );
  AND2X1 U2846 ( .A(n4050), .B(n1220), .Y(n1137) );
  AND2X1 U2847 ( .A(n4075), .B(n1222), .Y(n1138) );
  AND2X1 U2848 ( .A(n1436), .B(n1224), .Y(n1139) );
  AND2X1 U2849 ( .A(n1273), .B(n1226), .Y(n1140) );
  AND2X1 U2850 ( .A(n4148), .B(n1228), .Y(n1141) );
  AND2X1 U2851 ( .A(n1506), .B(n1230), .Y(n1142) );
  AND2X1 U2852 ( .A(n4198), .B(n1232), .Y(n1143) );
  AND2X1 U2853 ( .A(n1275), .B(n1234), .Y(n1144) );
  AND2X1 U2854 ( .A(n4272), .B(n1238), .Y(n1146) );
  AND2X1 U2855 ( .A(n4297), .B(n1240), .Y(n1147) );
  AND2X1 U2856 ( .A(n1277), .B(n1242), .Y(n1148) );
  AND2X1 U2857 ( .A(n4346), .B(n1244), .Y(n1149) );
  AND2X1 U2858 ( .A(n4371), .B(n1246), .Y(n1150) );
  AND2X1 U2859 ( .A(n1276), .B(n1248), .Y(n1151) );
  AND2X1 U2860 ( .A(n1445), .B(n1250), .Y(n1152) );
  AND2X1 U2861 ( .A(n4445), .B(n1252), .Y(n1153) );
  AND2X1 U2862 ( .A(n4470), .B(n1254), .Y(n1154) );
  AND2X1 U2863 ( .A(n1256), .B(n1274), .Y(n1155) );
  AND2X1 U2864 ( .A(n4521), .B(n1258), .Y(n1156) );
  AND2X1 U2865 ( .A(n4543), .B(n1278), .Y(n1157) );
  AND2X2 U2866 ( .A(\mem<3><2> ), .B(n800), .Y(n1158) );
  INVX1 U2867 ( .A(n1158), .Y(n1159) );
  AND2X2 U2868 ( .A(\mem<3><3> ), .B(n4471), .Y(n1160) );
  INVX1 U2869 ( .A(n1160), .Y(n1161) );
  AND2X2 U2870 ( .A(\mem<3><4> ), .B(n19), .Y(n1162) );
  INVX1 U2871 ( .A(n1162), .Y(n1163) );
  AND2X2 U2872 ( .A(\mem<3><5> ), .B(n19), .Y(n1164) );
  INVX1 U2873 ( .A(n1164), .Y(n1165) );
  AND2X2 U2874 ( .A(\mem<3><6> ), .B(n800), .Y(n1166) );
  INVX1 U2875 ( .A(n1166), .Y(n1167) );
  AND2X2 U2876 ( .A(\mem<3><7> ), .B(n4471), .Y(n1168) );
  INVX1 U2877 ( .A(n1168), .Y(n1169) );
  AND2X2 U2878 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n1170) );
  INVX1 U2879 ( .A(n1170), .Y(n1171) );
  AND2X1 U2880 ( .A(enable), .B(n1658), .Y(n1172) );
  INVX1 U2881 ( .A(n1172), .Y(n1173) );
  INVX1 U2882 ( .A(n1174), .Y(n1175) );
  INVX1 U2883 ( .A(n1176), .Y(n1177) );
  INVX1 U2884 ( .A(n1178), .Y(n1179) );
  INVX1 U2885 ( .A(n1180), .Y(n1181) );
  INVX1 U2886 ( .A(n1182), .Y(n1183) );
  INVX1 U2887 ( .A(n1184), .Y(n1185) );
  INVX1 U2888 ( .A(n1186), .Y(n1187) );
  INVX1 U2889 ( .A(n1188), .Y(n1189) );
  INVX1 U2890 ( .A(n1190), .Y(n1191) );
  INVX1 U2891 ( .A(n1192), .Y(n1193) );
  INVX1 U2892 ( .A(n1194), .Y(n1195) );
  INVX1 U2893 ( .A(n1196), .Y(n1197) );
  INVX1 U2894 ( .A(n1198), .Y(n1199) );
  INVX1 U2895 ( .A(n1200), .Y(n1201) );
  INVX1 U2896 ( .A(n1202), .Y(n1203) );
  INVX1 U2897 ( .A(n1204), .Y(n1205) );
  INVX1 U2898 ( .A(n1206), .Y(n1207) );
  INVX1 U2899 ( .A(n1208), .Y(n1209) );
  INVX1 U2900 ( .A(n1210), .Y(n1211) );
  INVX1 U2901 ( .A(n1212), .Y(n1213) );
  INVX1 U2902 ( .A(n1214), .Y(n1215) );
  INVX1 U2903 ( .A(n1216), .Y(n1217) );
  INVX1 U2904 ( .A(n1218), .Y(n1219) );
  INVX1 U2905 ( .A(n1220), .Y(n1221) );
  INVX1 U2906 ( .A(n1222), .Y(n1223) );
  INVX1 U2907 ( .A(n1224), .Y(n1225) );
  INVX1 U2908 ( .A(n1226), .Y(n1227) );
  INVX1 U2909 ( .A(n1228), .Y(n1229) );
  INVX1 U2910 ( .A(n1230), .Y(n1231) );
  INVX1 U2911 ( .A(n1232), .Y(n1233) );
  INVX1 U2912 ( .A(n1234), .Y(n1235) );
  INVX1 U2913 ( .A(n1236), .Y(n1237) );
  INVX1 U2914 ( .A(n1238), .Y(n1239) );
  INVX1 U2915 ( .A(n1240), .Y(n1241) );
  INVX1 U2916 ( .A(n1242), .Y(n1243) );
  INVX1 U2917 ( .A(n1244), .Y(n1245) );
  INVX1 U2918 ( .A(n1246), .Y(n1247) );
  INVX1 U2919 ( .A(n1248), .Y(n1249) );
  INVX1 U2920 ( .A(n1250), .Y(n1251) );
  INVX1 U2921 ( .A(n1252), .Y(n1253) );
  INVX1 U2922 ( .A(n1254), .Y(n1255) );
  INVX1 U2923 ( .A(n1256), .Y(n1257) );
  INVX1 U2924 ( .A(n1258), .Y(n1259) );
  INVX1 U2925 ( .A(n860), .Y(n1260) );
  AND2X2 U2926 ( .A(n1281), .B(n1444), .Y(n1261) );
  INVX1 U2927 ( .A(n1261), .Y(n1262) );
  INVX1 U2928 ( .A(n592), .Y(n1616) );
  INVX1 U2929 ( .A(n776), .Y(n1263) );
  INVX1 U2930 ( .A(n778), .Y(n1264) );
  INVX1 U2931 ( .A(n788), .Y(n1265) );
  INVX1 U2932 ( .A(n694), .Y(n1266) );
  INVX1 U2933 ( .A(n695), .Y(n1267) );
  INVX1 U2934 ( .A(n3166), .Y(n1268) );
  INVX1 U2935 ( .A(n1420), .Y(n1269) );
  INVX1 U2936 ( .A(n2978), .Y(n1270) );
  INVX1 U2937 ( .A(n797), .Y(n1271) );
  INVX1 U2938 ( .A(n813), .Y(n1272) );
  INVX1 U2939 ( .A(n699), .Y(n1273) );
  INVX1 U2940 ( .A(n18), .Y(n1274) );
  INVX1 U2941 ( .A(n801), .Y(n1275) );
  INVX1 U2942 ( .A(n35), .Y(n1276) );
  INVX1 U2943 ( .A(n140), .Y(n1277) );
  INVX1 U2944 ( .A(n591), .Y(n1619) );
  INVX1 U2945 ( .A(n1444), .Y(n1278) );
  INVX1 U2946 ( .A(n1649), .Y(n1279) );
  INVX1 U2947 ( .A(n721), .Y(n1280) );
  INVX1 U2948 ( .A(n1282), .Y(n1281) );
  BUFX2 U2949 ( .A(n625), .Y(n1282) );
  INVX1 U2950 ( .A(n139), .Y(n1284) );
  INVX1 U2951 ( .A(n139), .Y(n1285) );
  INVX1 U2952 ( .A(n832), .Y(n1286) );
  INVX1 U2953 ( .A(n137), .Y(n1287) );
  INVX1 U2954 ( .A(n137), .Y(n1288) );
  AND2X1 U2955 ( .A(n3006), .B(n2979), .Y(n1290) );
  INVX1 U2956 ( .A(n1290), .Y(n1291) );
  INVX1 U2957 ( .A(n1292), .Y(n1293) );
  AND2X1 U2958 ( .A(n3059), .B(n3033), .Y(n1294) );
  INVX1 U2959 ( .A(n1294), .Y(n1295) );
  INVX1 U2960 ( .A(n1296), .Y(n1297) );
  AND2X1 U2961 ( .A(n3113), .B(n3086), .Y(n1298) );
  INVX1 U2962 ( .A(n1298), .Y(n1299) );
  AND2X1 U2963 ( .A(n3114), .B(n3115), .Y(n1300) );
  INVX1 U2964 ( .A(n1300), .Y(n1301) );
  AND2X2 U2965 ( .A(n3166), .B(n1174), .Y(n1302) );
  INVX1 U2966 ( .A(n1302), .Y(n1303) );
  INVX1 U2967 ( .A(n1304), .Y(n1305) );
  AND2X2 U2968 ( .A(n854), .B(n1176), .Y(n1306) );
  INVX1 U2969 ( .A(n1306), .Y(n1307) );
  AND2X1 U2970 ( .A(n1420), .B(n1178), .Y(n1308) );
  INVX1 U2971 ( .A(n1308), .Y(n1309) );
  AND2X1 U2972 ( .A(n833), .B(n3243), .Y(n1310) );
  INVX1 U2973 ( .A(n1310), .Y(n1311) );
  AND2X2 U2974 ( .A(n3296), .B(n3270), .Y(n1312) );
  INVX1 U2975 ( .A(n1312), .Y(n1313) );
  AND2X1 U2976 ( .A(n1442), .B(n3297), .Y(n1314) );
  INVX1 U2977 ( .A(n1314), .Y(n1315) );
  AND2X1 U2978 ( .A(n1416), .B(n3325), .Y(n1316) );
  INVX1 U2979 ( .A(n1316), .Y(n1317) );
  AND2X2 U2980 ( .A(n835), .B(n1180), .Y(n1318) );
  INVX1 U2981 ( .A(n1318), .Y(n1319) );
  AND2X2 U2982 ( .A(n695), .B(n1182), .Y(n1320) );
  INVX1 U2983 ( .A(n1320), .Y(n1321) );
  AND2X2 U2984 ( .A(n832), .B(n1184), .Y(n1322) );
  INVX1 U2985 ( .A(n1322), .Y(n1323) );
  AND2X2 U2986 ( .A(n1459), .B(n1186), .Y(n1324) );
  INVX1 U2987 ( .A(n1324), .Y(n1325) );
  AND2X2 U2988 ( .A(n1466), .B(n1188), .Y(n1326) );
  INVX1 U2989 ( .A(n1326), .Y(n1327) );
  AND2X2 U2990 ( .A(n694), .B(n1190), .Y(n1328) );
  INVX1 U2991 ( .A(n1328), .Y(n1329) );
  AND2X2 U2992 ( .A(n860), .B(n1192), .Y(n1330) );
  INVX1 U2993 ( .A(n1330), .Y(n1331) );
  AND2X2 U2994 ( .A(n42), .B(n1194), .Y(n1332) );
  INVX1 U2995 ( .A(n1332), .Y(n1333) );
  AND2X1 U2996 ( .A(n1464), .B(n1196), .Y(n1334) );
  INVX1 U2997 ( .A(n1334), .Y(n1335) );
  AND2X2 U2998 ( .A(n790), .B(n1198), .Y(n1336) );
  INVX1 U2999 ( .A(n1336), .Y(n1337) );
  AND2X2 U3000 ( .A(n783), .B(n1200), .Y(n1338) );
  INVX1 U3001 ( .A(n1338), .Y(n1339) );
  AND2X2 U3002 ( .A(n791), .B(n1202), .Y(n1340) );
  INVX1 U3003 ( .A(n1340), .Y(n1341) );
  AND2X2 U3004 ( .A(n779), .B(n1204), .Y(n1342) );
  INVX1 U3005 ( .A(n1342), .Y(n1343) );
  AND2X2 U3006 ( .A(n777), .B(n1206), .Y(n1344) );
  INVX1 U3007 ( .A(n1344), .Y(n1345) );
  AND2X2 U3008 ( .A(n775), .B(n1208), .Y(n1346) );
  INVX1 U3009 ( .A(n1346), .Y(n1347) );
  AND2X2 U3010 ( .A(n3718), .B(n1210), .Y(n1348) );
  INVX1 U3011 ( .A(n1348), .Y(n1349) );
  AND2X2 U3012 ( .A(n788), .B(n1212), .Y(n1350) );
  INVX1 U3013 ( .A(n1350), .Y(n1351) );
  AND2X2 U3014 ( .A(n3793), .B(n3767), .Y(n1352) );
  INVX1 U3015 ( .A(n1352), .Y(n1353) );
  AND2X1 U3016 ( .A(n1418), .B(n3794), .Y(n1354) );
  INVX1 U3017 ( .A(n1354), .Y(n1355) );
  INVX1 U3018 ( .A(n1356), .Y(n1357) );
  AND2X1 U3019 ( .A(n1507), .B(n3847), .Y(n1358) );
  INVX1 U3020 ( .A(n1358), .Y(n1359) );
  INVX1 U3021 ( .A(n1360), .Y(n1361) );
  AND2X2 U3022 ( .A(n825), .B(n3900), .Y(n1362) );
  INVX1 U3023 ( .A(n1362), .Y(n1363) );
  AND2X1 U3024 ( .A(n3926), .B(n3927), .Y(n1364) );
  INVX1 U3025 ( .A(n1364), .Y(n1365) );
  AND2X2 U3026 ( .A(n797), .B(n1214), .Y(n1366) );
  INVX1 U3027 ( .A(n1366), .Y(n1367) );
  AND2X2 U3028 ( .A(n813), .B(n1216), .Y(n1368) );
  INVX1 U3029 ( .A(n1368), .Y(n1369) );
  AND2X2 U3030 ( .A(n1435), .B(n1218), .Y(n1370) );
  INVX1 U3031 ( .A(n1370), .Y(n1371) );
  AND2X2 U3032 ( .A(n782), .B(n1220), .Y(n1372) );
  INVX1 U3033 ( .A(n1372), .Y(n1373) );
  AND2X2 U3034 ( .A(n852), .B(n1222), .Y(n1374) );
  INVX1 U3035 ( .A(n1374), .Y(n1375) );
  AND2X2 U3036 ( .A(n13), .B(n1224), .Y(n1376) );
  INVX1 U3037 ( .A(n1376), .Y(n1377) );
  AND2X2 U3038 ( .A(n699), .B(n1226), .Y(n1378) );
  INVX1 U3039 ( .A(n1378), .Y(n1379) );
  AND2X2 U3040 ( .A(n780), .B(n1228), .Y(n1380) );
  INVX1 U3041 ( .A(n1380), .Y(n1381) );
  INVX1 U3042 ( .A(n1382), .Y(n1383) );
  AND2X2 U3043 ( .A(n851), .B(n1232), .Y(n1384) );
  INVX1 U3044 ( .A(n1384), .Y(n1385) );
  AND2X2 U3045 ( .A(n801), .B(n1234), .Y(n1386) );
  INVX1 U3046 ( .A(n1386), .Y(n1387) );
  AND2X2 U3047 ( .A(n26), .B(n1236), .Y(n1388) );
  INVX1 U3048 ( .A(n1388), .Y(n1389) );
  AND2X2 U3049 ( .A(n1458), .B(n1238), .Y(n1390) );
  INVX1 U3050 ( .A(n1390), .Y(n1391) );
  AND2X2 U3051 ( .A(n847), .B(n1240), .Y(n1392) );
  INVX1 U3052 ( .A(n1392), .Y(n1393) );
  AND2X2 U3053 ( .A(n140), .B(n1242), .Y(n1394) );
  INVX1 U3054 ( .A(n1394), .Y(n1395) );
  AND2X1 U3055 ( .A(n1478), .B(n1244), .Y(n1396) );
  INVX1 U3056 ( .A(n1396), .Y(n1397) );
  AND2X2 U3057 ( .A(n10), .B(n1246), .Y(n1398) );
  INVX1 U3058 ( .A(n1398), .Y(n1399) );
  AND2X2 U3059 ( .A(n35), .B(n1248), .Y(n1400) );
  INVX1 U3060 ( .A(n1400), .Y(n1401) );
  AND2X2 U3061 ( .A(n823), .B(n1250), .Y(n1402) );
  INVX1 U3062 ( .A(n1402), .Y(n1403) );
  AND2X2 U3063 ( .A(n1486), .B(n1252), .Y(n1404) );
  INVX1 U3064 ( .A(n1404), .Y(n1405) );
  AND2X2 U3065 ( .A(n816), .B(n1254), .Y(n1406) );
  INVX1 U3066 ( .A(n1406), .Y(n1407) );
  AND2X2 U3067 ( .A(n800), .B(n1256), .Y(n1408) );
  INVX1 U3068 ( .A(n1408), .Y(n1409) );
  AND2X2 U3069 ( .A(n787), .B(n1258), .Y(n1410) );
  INVX1 U3070 ( .A(n1410), .Y(n1411) );
  AND2X2 U3071 ( .A(n1444), .B(n4543), .Y(n1412) );
  INVX1 U3072 ( .A(n1412), .Y(n1413) );
  OAI21X1 U3073 ( .A(n1683), .B(n802), .C(n969), .Y(n1686) );
  INVX1 U3074 ( .A(\mem<25><1> ), .Y(n1683) );
  INVX1 U3075 ( .A(n585), .Y(n3497) );
  NOR2X1 U3076 ( .A(\addr<12> ), .B(\addr<11> ), .Y(n1581) );
  OAI21X1 U3077 ( .A(n1668), .B(n3141), .C(n1667), .Y(n1671) );
  INVX1 U3078 ( .A(\mem<57><1> ), .Y(n1668) );
  INVX4 U3079 ( .A(n1526), .Y(n3141) );
  OAI21X1 U3080 ( .A(n1669), .B(n3087), .C(n834), .Y(n1670) );
  INVX1 U3081 ( .A(\mem<58><1> ), .Y(n1669) );
  INVX1 U3082 ( .A(N182), .Y(n1414) );
  AND2X2 U3083 ( .A(n774), .B(n789), .Y(n1415) );
  BUFX2 U3084 ( .A(n821), .Y(n1416) );
  INVX1 U3085 ( .A(n686), .Y(n1417) );
  INVX1 U3086 ( .A(n3795), .Y(n1418) );
  MUX2X1 U3087 ( .B(\mem<27><6> ), .A(\mem<26><6> ), .S(n1524), .Y(n2908) );
  MUX2X1 U3088 ( .B(\mem<31><6> ), .A(\mem<30><6> ), .S(n1550), .Y(n2910) );
  INVX1 U3089 ( .A(n662), .Y(n1419) );
  BUFX2 U3090 ( .A(n6), .Y(n1420) );
  MUX2X1 U3091 ( .B(n135), .A(n2801), .S(n1421), .Y(n2805) );
  BUFX2 U3092 ( .A(n598), .Y(n1422) );
  MUX2X1 U3093 ( .B(n2899), .A(n2898), .S(n1423), .Y(n2900) );
  INVX8 U3094 ( .A(n1427), .Y(n1423) );
  MUX2X1 U3095 ( .B(\mem<60><6> ), .A(\mem<61><6> ), .S(n1452), .Y(n2867) );
  MUX2X1 U3096 ( .B(\mem<17><6> ), .A(\mem<16><6> ), .S(n1487), .Y(n2879) );
  MUX2X1 U3097 ( .B(\mem<39><7> ), .A(\mem<38><7> ), .S(n1550), .Y(n2933) );
  MUX2X1 U3098 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1542), .Y(n2911) );
  INVX4 U3099 ( .A(N180), .Y(n1424) );
  INVX1 U3100 ( .A(n5), .Y(n1579) );
  INVX1 U3101 ( .A(n794), .Y(n1425) );
  MUX2X1 U3102 ( .B(n2861), .A(n2860), .S(n1558), .Y(n2862) );
  NOR3X1 U3103 ( .A(\addr<14> ), .B(\addr<13> ), .C(\addr<15> ), .Y(n1426) );
  INVX1 U3104 ( .A(n1578), .Y(n1428) );
  AND2X2 U3105 ( .A(N181), .B(N182), .Y(n1429) );
  MUX2X1 U3106 ( .B(\mem<41><6> ), .A(\mem<40><6> ), .S(n1550), .Y(n2889) );
  MUX2X1 U3107 ( .B(\mem<53><5> ), .A(\mem<52><5> ), .S(n1483), .Y(n2843) );
  MUX2X1 U3108 ( .B(n2716), .A(n2717), .S(n1430), .Y(n2718) );
  INVX1 U3109 ( .A(N177), .Y(n1431) );
  INVX1 U3110 ( .A(N177), .Y(n1535) );
  INVX1 U3111 ( .A(n1540), .Y(n1433) );
  MUX2X1 U3112 ( .B(\mem<63><5> ), .A(\mem<62><5> ), .S(n1550), .Y(n2837) );
  MUX2X1 U3113 ( .B(n2931), .A(n2930), .S(n1570), .Y(n2932) );
  INVX1 U3114 ( .A(n1475), .Y(n1434) );
  MUX2X1 U3115 ( .B(\mem<33><5> ), .A(\mem<32><5> ), .S(n1487), .Y(n2831) );
  AND2X2 U3116 ( .A(n517), .B(n1651), .Y(n1435) );
  INVX1 U3117 ( .A(n1435), .Y(n4025) );
  MUX2X1 U3118 ( .B(\mem<43><6> ), .A(\mem<42><6> ), .S(n841), .Y(n2888) );
  MUX2X1 U3119 ( .B(\mem<25><6> ), .A(\mem<24><6> ), .S(n1548), .Y(n2909) );
  INVX1 U3120 ( .A(n720), .Y(n1436) );
  MUX2X1 U3121 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1454), .Y(n2807) );
  MUX2X1 U3122 ( .B(n2892), .A(n2893), .S(n1437), .Y(n2901) );
  INVX1 U3123 ( .A(n1579), .Y(n1577) );
  MUX2X1 U3124 ( .B(\mem<17><5> ), .A(\mem<16><5> ), .S(n38), .Y(n2824) );
  MUX2X1 U3125 ( .B(\mem<21><5> ), .A(\mem<20><5> ), .S(n1551), .Y(n2821) );
  INVX8 U3126 ( .A(n1548), .Y(n1545) );
  MUX2X1 U3127 ( .B(\mem<41><5> ), .A(\mem<40><5> ), .S(n1474), .Y(n2853) );
  MUX2X1 U3128 ( .B(\mem<3><7> ), .A(\mem<2><7> ), .S(n826), .Y(n2919) );
  INVX1 U3129 ( .A(n50), .Y(n1438) );
  MUX2X1 U3130 ( .B(n2862), .A(n2863), .S(n1427), .Y(n2871) );
  MUX2X1 U3131 ( .B(\mem<5><6> ), .A(\mem<4><6> ), .S(n841), .Y(n2861) );
  MUX2X1 U3132 ( .B(\mem<23><5> ), .A(\mem<22><5> ), .S(n1487), .Y(n2820) );
  INVX8 U3133 ( .A(n1489), .Y(n1544) );
  MUX2X1 U3134 ( .B(\mem<7><7> ), .A(\mem<6><7> ), .S(n1487), .Y(n2921) );
  MUX2X1 U3135 ( .B(\mem<1><7> ), .A(\mem<0><7> ), .S(n1550), .Y(n2920) );
  MUX2X1 U3136 ( .B(n2919), .A(n2920), .S(n1439), .Y(n2924) );
  INVX8 U3137 ( .A(n1548), .Y(n1542) );
  MUX2X1 U3138 ( .B(\mem<39><6> ), .A(\mem<38><6> ), .S(n841), .Y(n2904) );
  MUX2X1 U3139 ( .B(\mem<37><6> ), .A(\mem<36><6> ), .S(n1474), .Y(n2905) );
  MUX2X1 U3140 ( .B(\mem<5><7> ), .A(\mem<4><7> ), .S(n1433), .Y(n2922) );
  MUX2X1 U3141 ( .B(\mem<19><7> ), .A(\mem<18><7> ), .S(n38), .Y(n2949) );
  MUX2X1 U3142 ( .B(\mem<15><7> ), .A(\mem<14><7> ), .S(n1474), .Y(n2928) );
  INVX1 U3143 ( .A(n1533), .Y(n1441) );
  INVX8 U3144 ( .A(n1564), .Y(n1563) );
  MUX2X1 U3145 ( .B(\mem<13><7> ), .A(\mem<12><7> ), .S(n1549), .Y(n2929) );
  MUX2X1 U3146 ( .B(n2877), .A(n2876), .S(n1570), .Y(n2885) );
  MUX2X1 U3147 ( .B(\mem<35><7> ), .A(\mem<34><7> ), .S(n40), .Y(n2935) );
  INVX2 U3148 ( .A(n1496), .Y(n2475) );
  INVX1 U3149 ( .A(n1476), .Y(n1442) );
  AND2X2 U3150 ( .A(n1485), .B(n1585), .Y(n1443) );
  INVX1 U3151 ( .A(n666), .Y(n1444) );
  AND2X2 U3152 ( .A(n1524), .B(n30), .Y(n1650) );
  INVX1 U3153 ( .A(n823), .Y(n1445) );
  INVX2 U3154 ( .A(n826), .Y(n1543) );
  INVX1 U3155 ( .A(n783), .Y(n3620) );
  AND2X2 U3156 ( .A(n1438), .B(n53), .Y(n1446) );
  INVX1 U3157 ( .A(n853), .Y(n4272) );
  INVX1 U3158 ( .A(\addr<11> ), .Y(n1448) );
  INVX1 U3159 ( .A(n1448), .Y(n1449) );
  INVX1 U3160 ( .A(n1534), .Y(n1450) );
  AND2X2 U3161 ( .A(n1649), .B(n1648), .Y(n1451) );
  INVX1 U3162 ( .A(n1451), .Y(n4371) );
  MUX2X1 U3163 ( .B(n2906), .A(n2907), .S(n1437), .Y(n2915) );
  MUX2X1 U3164 ( .B(n2858), .A(n2859), .S(n58), .Y(n2863) );
  INVX1 U3165 ( .A(n1550), .Y(n1452) );
  INVX1 U3166 ( .A(n1550), .Y(n1453) );
  INVX1 U3167 ( .A(n1450), .Y(n1540) );
  AND2X2 U3168 ( .A(n1093), .B(n53), .Y(n1455) );
  INVX1 U3169 ( .A(n851), .Y(n4198) );
  AND2X2 U3170 ( .A(n1649), .B(n651), .Y(n1456) );
  INVX1 U3171 ( .A(n1456), .Y(n3571) );
  MUX2X1 U3172 ( .B(\mem<31><7> ), .A(\mem<30><7> ), .S(n1550), .Y(n2938) );
  INVX1 U3173 ( .A(n1446), .Y(n1457) );
  INVX1 U3174 ( .A(n1457), .Y(n1458) );
  MUX2X1 U3175 ( .B(\mem<25><7> ), .A(\mem<24><7> ), .S(n1549), .Y(n2942) );
  MUX2X1 U3176 ( .B(n2869), .A(n2868), .S(n1570), .Y(n2870) );
  INVX1 U3177 ( .A(n1289), .Y(n1459) );
  INVX1 U3178 ( .A(n3571), .Y(n1460) );
  NAND2X1 U3179 ( .A(n2970), .B(n1461), .Y(n1462) );
  NAND2X1 U3180 ( .A(n1555), .B(n2969), .Y(n1463) );
  INVX1 U3181 ( .A(n1555), .Y(n1461) );
  INVX8 U3182 ( .A(n1552), .Y(n1565) );
  BUFX2 U3183 ( .A(n1460), .Y(n1464) );
  INVX1 U3184 ( .A(n852), .Y(n4075) );
  INVX1 U3185 ( .A(n515), .Y(n1481) );
  INVX8 U3186 ( .A(n1553), .Y(n1567) );
  MUX2X1 U3187 ( .B(n2744), .A(n2743), .S(n1570), .Y(n2745) );
  AND2X2 U3188 ( .A(n49), .B(n792), .Y(n1468) );
  INVX1 U3189 ( .A(n1466), .Y(n3472) );
  AND2X2 U3190 ( .A(n513), .B(n53), .Y(n1469) );
  INVX1 U3191 ( .A(n847), .Y(n4297) );
  AND2X2 U3192 ( .A(n1470), .B(n74), .Y(n1665) );
  INVX1 U3193 ( .A(n43), .Y(n3546) );
  AND2X2 U3194 ( .A(n1650), .B(n1505), .Y(n1472) );
  INVX1 U3195 ( .A(n1472), .Y(n4346) );
  NOR2X1 U3196 ( .A(\addr<7> ), .B(\addr<6> ), .Y(n1473) );
  INVX1 U3197 ( .A(n1441), .Y(n1475) );
  INVX1 U3198 ( .A(n839), .Y(n1476) );
  INVX1 U3199 ( .A(N181), .Y(n2688) );
  MUX2X1 U3200 ( .B(\mem<21><4> ), .A(\mem<20><4> ), .S(n1487), .Y(n2749) );
  INVX1 U3201 ( .A(n833), .Y(n1477) );
  INVX8 U3202 ( .A(n1554), .Y(n1552) );
  INVX8 U3203 ( .A(n1552), .Y(n1566) );
  BUFX2 U3204 ( .A(n1472), .Y(n1478) );
  NAND2X1 U3205 ( .A(n799), .B(n1479), .Y(n1480) );
  INVX1 U3206 ( .A(n4774), .Y(n1479) );
  OR2X2 U3207 ( .A(n713), .B(n1481), .Y(n3218) );
  INVX1 U3208 ( .A(n1602), .Y(n1606) );
  MUX2X1 U3209 ( .B(\mem<33><6> ), .A(\mem<32><6> ), .S(n1440), .Y(n2903) );
  INVX1 U3210 ( .A(n842), .Y(n1482) );
  MUX2X1 U3211 ( .B(\mem<51><7> ), .A(\mem<50><7> ), .S(n1550), .Y(n2966) );
  MUX2X1 U3212 ( .B(\mem<57><7> ), .A(\mem<56><7> ), .S(n1549), .Y(n2960) );
  MUX2X1 U3213 ( .B(\mem<13><6> ), .A(\mem<12><6> ), .S(n1548), .Y(n2875) );
  INVX1 U3214 ( .A(n816), .Y(n4470) );
  MUX2X1 U3215 ( .B(\mem<17><7> ), .A(\mem<16><7> ), .S(n1549), .Y(n2950) );
  MUX2X1 U3216 ( .B(\mem<33><7> ), .A(\mem<32><7> ), .S(n1549), .Y(n2936) );
  INVX1 U3217 ( .A(n1486), .Y(n4445) );
  INVX1 U3218 ( .A(n1534), .Y(n1488) );
  MUX2X1 U3219 ( .B(\mem<21><7> ), .A(\mem<20><7> ), .S(n1440), .Y(n2947) );
  INVX1 U3220 ( .A(n781), .Y(n4148) );
  MUX2X1 U3221 ( .B(\mem<11><6> ), .A(\mem<10><6> ), .S(n1450), .Y(n2872) );
  MUX2X1 U3222 ( .B(\mem<9><6> ), .A(\mem<8><6> ), .S(n1474), .Y(n2873) );
  BUFX4 U3223 ( .A(n1535), .Y(n1489) );
  MUX2X1 U3224 ( .B(\mem<41><7> ), .A(\mem<40><7> ), .S(n1550), .Y(n2972) );
  MUX2X1 U3225 ( .B(\mem<27><4> ), .A(\mem<26><4> ), .S(n1434), .Y(n2739) );
  NAND2X1 U3226 ( .A(\mem<10><5> ), .B(n1490), .Y(n1491) );
  NAND2X1 U3227 ( .A(\mem<11><5> ), .B(n1484), .Y(n1492) );
  INVX1 U3228 ( .A(n1485), .Y(n1490) );
  NAND2X1 U3229 ( .A(\mem<34><3> ), .B(n1493), .Y(n1494) );
  NAND2X1 U3230 ( .A(\mem<35><3> ), .B(n1454), .Y(n1495) );
  NOR3X1 U3231 ( .A(n138), .B(n1498), .C(n1497), .Y(n1496) );
  OR2X2 U3232 ( .A(n1626), .B(n1625), .Y(n1498) );
  INVX1 U3233 ( .A(n1288), .Y(n1659) );
  INVX1 U3234 ( .A(n1287), .Y(n1584) );
  MUX2X1 U3235 ( .B(\mem<5><5> ), .A(\mem<4><5> ), .S(n1450), .Y(n2803) );
  BUFX2 U3236 ( .A(\addr<14> ), .Y(n1501) );
  INVX1 U3237 ( .A(n786), .Y(n4521) );
  MUX2X1 U3238 ( .B(\mem<7><5> ), .A(\mem<6><5> ), .S(n1551), .Y(n2802) );
  INVX1 U3239 ( .A(n611), .Y(n1504) );
  AND2X2 U3240 ( .A(n629), .B(n632), .Y(n1505) );
  INVX1 U3241 ( .A(n90), .Y(n1506) );
  INVX1 U3242 ( .A(n610), .Y(n4149) );
  AND2X2 U3243 ( .A(n246), .B(n289), .Y(n2916) );
  BUFX2 U3244 ( .A(n842), .Y(n1507) );
  INVX8 U3245 ( .A(n1548), .Y(n1546) );
  MUX2X1 U3246 ( .B(\mem<1><5> ), .A(\mem<0><5> ), .S(n1550), .Y(n2801) );
  AND2X2 U3247 ( .A(n822), .B(n93), .Y(n1508) );
  INVX4 U3248 ( .A(N178), .Y(n1554) );
  MUX2X1 U3249 ( .B(\mem<3><6> ), .A(\mem<2><6> ), .S(n1548), .Y(n2858) );
  NAND2X1 U3250 ( .A(\mem<2><5> ), .B(n1509), .Y(n1510) );
  NAND2X1 U3251 ( .A(\mem<3><5> ), .B(n1484), .Y(n1511) );
  INVX1 U3252 ( .A(n1540), .Y(n1509) );
  NAND2X1 U3253 ( .A(\mem<40><0> ), .B(n1415), .Y(n1512) );
  AND2X2 U3254 ( .A(n1512), .B(n1513), .Y(n1596) );
  NOR3X1 U3255 ( .A(\addr<9> ), .B(\addr<10> ), .C(\addr<8> ), .Y(n1514) );
  INVX1 U3256 ( .A(n1568), .Y(n1575) );
  INVX1 U3257 ( .A(N179), .Y(n1569) );
  NOR3X1 U3258 ( .A(N182), .B(n717), .C(n711), .Y(n1515) );
  INVX1 U3259 ( .A(n718), .Y(n1601) );
  INVX1 U3260 ( .A(n45), .Y(n1600) );
  INVX1 U3261 ( .A(N182), .Y(n1634) );
  INVX1 U3262 ( .A(n1553), .Y(n1525) );
  MUX2X1 U3263 ( .B(\mem<61><7> ), .A(\mem<60><7> ), .S(n1548), .Y(n2957) );
  NAND3X1 U3264 ( .A(n1574), .B(n1552), .C(n39), .Y(n1516) );
  INVX1 U3265 ( .A(n782), .Y(n4050) );
  INVX1 U3266 ( .A(n803), .Y(n3926) );
  INVX1 U3267 ( .A(n1569), .Y(n1568) );
  INVX1 U3268 ( .A(n1568), .Y(n1576) );
  NAND2X1 U3269 ( .A(n1519), .B(n2934), .Y(n1520) );
  NAND2X1 U3270 ( .A(n2933), .B(n1555), .Y(n1521) );
  INVX1 U3271 ( .A(n1555), .Y(n1519) );
  AND2X2 U3272 ( .A(n1649), .B(n1611), .Y(n1522) );
  INVX1 U3273 ( .A(n835), .Y(n3375) );
  INVX1 U3274 ( .A(n1541), .Y(n1524) );
  AND2X2 U3275 ( .A(n515), .B(n685), .Y(n1523) );
  AND2X2 U3276 ( .A(n1616), .B(n1650), .Y(n1526) );
  INVX4 U3277 ( .A(n2977), .Y(n2978) );
  INVX4 U3278 ( .A(n1284), .Y(n3793) );
  INVX8 U3279 ( .A(n47), .Y(n1550) );
  INVX8 U3280 ( .A(n1567), .Y(n1555) );
  INVX8 U3281 ( .A(n1567), .Y(n1556) );
  INVX8 U3282 ( .A(n1566), .Y(n1557) );
  INVX8 U3283 ( .A(n1566), .Y(n1559) );
  INVX8 U3284 ( .A(n1565), .Y(n1560) );
  INVX8 U3285 ( .A(n1565), .Y(n1561) );
  INVX8 U3286 ( .A(n1565), .Y(n1562) );
  NAND3X1 U3287 ( .A(n1572), .B(n1553), .C(n1475), .Y(n2975) );
  NOR3X1 U3288 ( .A(\addr<9> ), .B(\addr<10> ), .C(\addr<8> ), .Y(n1583) );
  NOR3X1 U3289 ( .A(\addr<14> ), .B(\addr<13> ), .C(\addr<15> ), .Y(n1582) );
  NAND2X1 U3290 ( .A(\mem<32><0> ), .B(n649), .Y(n1589) );
  NAND2X1 U3291 ( .A(\mem<33><0> ), .B(n1584), .Y(n1588) );
  NOR2X1 U3292 ( .A(n1552), .B(n1571), .Y(n1585) );
  AND2X2 U3293 ( .A(n1485), .B(n95), .Y(n1655) );
  NAND3X1 U3294 ( .A(n1573), .B(n1553), .C(n1483), .Y(n1586) );
  AOI22X1 U3295 ( .A(\mem<34><0> ), .B(n673), .C(\mem<35><0> ), .D(n3669), .Y(
        n1587) );
  NAND3X1 U3296 ( .A(n1572), .B(n1564), .C(n32), .Y(n1590) );
  NAND3X1 U3297 ( .A(n1572), .B(n1552), .C(n38), .Y(n1591) );
  AOI22X1 U3298 ( .A(\mem<38><0> ), .B(n647), .C(\mem<39><0> ), .D(n654), .Y(
        n1594) );
  NAND3X1 U3299 ( .A(n1572), .B(n1565), .C(n1549), .Y(n1592) );
  AOI22X1 U3300 ( .A(\mem<36><0> ), .B(n638), .C(\mem<37><0> ), .D(n656), .Y(
        n1593) );
  AOI22X1 U3301 ( .A(\mem<42><0> ), .B(n3497), .C(\mem<43><0> ), .D(n694), .Y(
        n1597) );
  AOI22X1 U3302 ( .A(\mem<46><0> ), .B(n1502), .C(\mem<47><0> ), .D(n695), .Y(
        n1599) );
  NAND3X1 U3303 ( .A(n1601), .B(n1600), .C(N182), .Y(n1602) );
  NOR2X1 U3304 ( .A(n711), .B(n1578), .Y(n1603) );
  NAND2X1 U3305 ( .A(\mem<56><0> ), .B(n793), .Y(n1604) );
  OAI21X1 U3306 ( .A(n3141), .B(n1605), .C(n1604), .Y(n1610) );
  NAND2X1 U3307 ( .A(\mem<59><0> ), .B(n522), .Y(n1607) );
  OAI21X1 U3308 ( .A(n3087), .B(n1608), .C(n1607), .Y(n1609) );
  AOI22X1 U3309 ( .A(\mem<50><0> ), .B(n3323), .C(\mem<51><0> ), .D(n3296), 
        .Y(n1613) );
  AOI22X1 U3310 ( .A(\mem<48><0> ), .B(n1500), .C(\mem<49><0> ), .D(n3324), 
        .Y(n1612) );
  AOI22X1 U3311 ( .A(\mem<52><0> ), .B(n3269), .C(\mem<53><0> ), .D(n698), .Y(
        n1614) );
  NAND2X1 U3312 ( .A(\mem<61><0> ), .B(n662), .Y(n1617) );
  OAI21X1 U3313 ( .A(n634), .B(n1618), .C(n1617), .Y(n1623) );
  NAND2X1 U3314 ( .A(\mem<63><0> ), .B(n2978), .Y(n1620) );
  OAI21X1 U3315 ( .A(n2980), .B(n1621), .C(n1620), .Y(n1622) );
  NAND2X1 U3316 ( .A(n1501), .B(\addr<15> ), .Y(n1624) );
  NAND2X1 U3317 ( .A(\addr<8> ), .B(n844), .Y(n1626) );
  NAND2X1 U3318 ( .A(n1449), .B(n806), .Y(n1625) );
  NAND3X1 U3319 ( .A(n1485), .B(n1570), .C(n1563), .Y(n1628) );
  NAND3X1 U3320 ( .A(N181), .B(N182), .C(n1578), .Y(n1627) );
  NOR3X1 U3321 ( .A(n1171), .B(n1627), .C(n1628), .Y(n1629) );
  OAI21X1 U3322 ( .A(n803), .B(n1630), .C(n965), .Y(n1633) );
  AND2X2 U3323 ( .A(n822), .B(n93), .Y(n1651) );
  OAI21X1 U3324 ( .A(n671), .B(n1631), .C(n967), .Y(n1632) );
  AOI22X1 U3325 ( .A(\mem<19><0> ), .B(n720), .C(\mem<16><0> ), .D(n90), .Y(
        n1636) );
  AOI22X1 U3326 ( .A(\mem<21><0> ), .B(n1517), .C(\mem<18><0> ), .D(n699), .Y(
        n1637) );
  OAI21X1 U3327 ( .A(n1283), .B(n1639), .C(n319), .Y(n1643) );
  NAND2X1 U3328 ( .A(\mem<28><0> ), .B(n842), .Y(n1640) );
  OAI21X1 U3329 ( .A(n1285), .B(n1641), .C(n1640), .Y(n1642) );
  AOI22X1 U3330 ( .A(\mem<2><0> ), .B(n1503), .C(\mem<3><0> ), .D(n4471), .Y(
        n1645) );
  AOI22X1 U3331 ( .A(\mem<1><0> ), .B(n665), .C(\mem<14><0> ), .D(n4199), .Y(
        n1644) );
  AOI22X1 U3332 ( .A(\mem<6><0> ), .B(n16), .C(\mem<7><0> ), .D(n55), .Y(n1647) );
  AOI22X1 U3333 ( .A(\mem<4><0> ), .B(n21), .C(\mem<5><0> ), .D(n689), .Y(
        n1646) );
  AOI22X1 U3334 ( .A(\mem<11><0> ), .B(n846), .C(\mem<8><0> ), .D(n20), .Y(
        n1653) );
  AOI22X1 U3335 ( .A(\mem<9><0> ), .B(n1472), .C(\mem<22><0> ), .D(n1435), .Y(
        n1652) );
  AOI22X1 U3336 ( .A(\mem<15><0> ), .B(n1455), .C(\mem<12><0> ), .D(n1446), 
        .Y(n1657) );
  AOI22X1 U3337 ( .A(\mem<13><0> ), .B(n56), .C(\mem<10><0> ), .D(n140), .Y(
        n1656) );
  AOI21X1 U3338 ( .A(n59), .B(n11), .C(n1173), .Y(\data_out<0> ) );
  AOI22X1 U3339 ( .A(\mem<34><1> ), .B(n673), .C(\mem<35><1> ), .D(n3669), .Y(
        n1660) );
  AOI22X1 U3340 ( .A(\mem<38><1> ), .B(n647), .C(\mem<39><1> ), .D(n654), .Y(
        n1662) );
  AOI22X1 U3341 ( .A(\mem<36><1> ), .B(n638), .C(\mem<37><1> ), .D(n656), .Y(
        n1661) );
  AOI22X1 U3342 ( .A(\mem<42><1> ), .B(n3), .C(\mem<43><1> ), .D(n694), .Y(
        n1664) );
  AOI22X1 U3343 ( .A(\mem<40><1> ), .B(n1456), .C(\mem<41><1> ), .D(n1471), 
        .Y(n1663) );
  AOI22X1 U3344 ( .A(\mem<46><1> ), .B(n1502), .C(\mem<47><1> ), .D(n695), .Y(
        n1666) );
  NAND2X1 U3345 ( .A(\mem<56><1> ), .B(n51), .Y(n1667) );
  AOI22X1 U3346 ( .A(\mem<50><1> ), .B(n3323), .C(\mem<51><1> ), .D(n3296), 
        .Y(n1673) );
  AOI22X1 U3347 ( .A(\mem<48><1> ), .B(n1522), .C(\mem<49><1> ), .D(n3324), 
        .Y(n1672) );
  AOI22X1 U3348 ( .A(\mem<54><1> ), .B(n14), .C(\mem<55><1> ), .D(n3167), .Y(
        n1675) );
  AOI22X1 U3349 ( .A(\mem<52><1> ), .B(n3269), .C(\mem<53><1> ), .D(n698), .Y(
        n1674) );
  NAND2X1 U3350 ( .A(\mem<61><1> ), .B(n662), .Y(n1676) );
  OAI21X1 U3351 ( .A(n634), .B(n1677), .C(n1676), .Y(n1681) );
  NAND2X1 U3352 ( .A(\mem<63><1> ), .B(n2978), .Y(n1678) );
  OAI21X1 U3353 ( .A(n2980), .B(n1679), .C(n1678), .Y(n1680) );
  OAI21X1 U3354 ( .A(n1684), .B(n672), .C(n729), .Y(n1685) );
  AOI22X1 U3355 ( .A(\mem<19><1> ), .B(n13), .C(\mem<16><1> ), .D(n4149), .Y(
        n1687) );
  NAND3X1 U3356 ( .A(n490), .B(n770), .C(n1687), .Y(n1690) );
  AOI22X1 U3357 ( .A(\mem<23><1> ), .B(n813), .C(\mem<20><1> ), .D(n785), .Y(
        n1689) );
  AOI22X1 U3358 ( .A(\mem<21><1> ), .B(n1517), .C(\mem<18><1> ), .D(n699), .Y(
        n1688) );
  NAND2X1 U3359 ( .A(\mem<28><1> ), .B(n842), .Y(n1691) );
  AOI22X1 U3360 ( .A(\mem<2><1> ), .B(n1503), .C(\mem<3><1> ), .D(n18), .Y(
        n1693) );
  AOI22X1 U3361 ( .A(\mem<1><1> ), .B(n665), .C(\mem<14><1> ), .D(n4199), .Y(
        n1692) );
  AOI22X1 U3362 ( .A(\mem<6><1> ), .B(n4396), .C(\mem<7><1> ), .D(n55), .Y(
        n1695) );
  AOI22X1 U3363 ( .A(\mem<4><1> ), .B(n1447), .C(\mem<5><1> ), .D(n689), .Y(
        n1694) );
  AOI22X1 U3364 ( .A(\mem<11><1> ), .B(n846), .C(\mem<8><1> ), .D(n57), .Y(
        n1697) );
  AOI22X1 U3365 ( .A(\mem<9><1> ), .B(n1472), .C(\mem<22><1> ), .D(n1435), .Y(
        n1696) );
  AOI22X1 U3366 ( .A(\mem<15><1> ), .B(n1455), .C(\mem<12><1> ), .D(n1446), 
        .Y(n1699) );
  AOI22X1 U3367 ( .A(\mem<13><1> ), .B(n56), .C(\mem<10><1> ), .D(n140), .Y(
        n1698) );
  AOI21X1 U3368 ( .A(n27), .B(n532), .C(n1173), .Y(\data_out<1> ) );
  AOI22X1 U3369 ( .A(\mem<35><2> ), .B(n777), .C(\mem<34><2> ), .D(n775), .Y(
        n1701) );
  INVX2 U3370 ( .A(n81), .Y(n3718) );
  AOI22X1 U3371 ( .A(\mem<33><2> ), .B(n3718), .C(\mem<32><2> ), .D(n788), .Y(
        n1700) );
  AOI22X1 U3372 ( .A(\mem<39><2> ), .B(n790), .C(\mem<38><2> ), .D(n783), .Y(
        n1703) );
  AOI22X1 U3373 ( .A(\mem<37><2> ), .B(n791), .C(\mem<36><2> ), .D(n85), .Y(
        n1702) );
  AOI22X1 U3374 ( .A(\mem<43><2> ), .B(n694), .C(\mem<42><2> ), .D(n860), .Y(
        n1705) );
  AOI22X1 U3375 ( .A(\mem<41><2> ), .B(n43), .C(\mem<40><2> ), .D(n1415), .Y(
        n1704) );
  AOI22X1 U3376 ( .A(\mem<47><2> ), .B(n695), .C(\mem<46><2> ), .D(n832), .Y(
        n1707) );
  AOI22X1 U3377 ( .A(\mem<45><2> ), .B(n8), .C(\mem<44><2> ), .D(n1466), .Y(
        n1706) );
  OAI21X1 U3378 ( .A(n634), .B(n1708), .C(n971), .Y(n1711) );
  OAI21X1 U3379 ( .A(n2980), .B(n1709), .C(n973), .Y(n1710) );
  OAI21X1 U3380 ( .A(n3141), .B(n1712), .C(n321), .Y(n1715) );
  OAI21X1 U3381 ( .A(n3087), .B(n1713), .C(n975), .Y(n1714) );
  AOI22X1 U3382 ( .A(\mem<51><2> ), .B(n3296), .C(\mem<50><2> ), .D(n840), .Y(
        n1717) );
  AOI22X1 U3383 ( .A(\mem<49><2> ), .B(n796), .C(\mem<48><2> ), .D(n1500), .Y(
        n1716) );
  AOI22X1 U3384 ( .A(\mem<55><2> ), .B(n831), .C(\mem<54><2> ), .D(n854), .Y(
        n1719) );
  AOI22X1 U3385 ( .A(\mem<53><2> ), .B(n698), .C(\mem<52><2> ), .D(n833), .Y(
        n1718) );
  NAND3X1 U3386 ( .A(n148), .B(n150), .C(n563), .Y(n1720) );
  OAI21X1 U3387 ( .A(n1482), .B(n1721), .C(n731), .Y(n1725) );
  NAND2X1 U3388 ( .A(\mem<31><2> ), .B(n3793), .Y(n1722) );
  OAI21X1 U3389 ( .A(n3795), .B(n1723), .C(n1722), .Y(n1724) );
  OAI21X1 U3390 ( .A(n802), .B(n1726), .C(n977), .Y(n1729) );
  OAI21X1 U3391 ( .A(n849), .B(n1727), .C(n323), .Y(n1728) );
  AOI22X1 U3392 ( .A(\mem<19><2> ), .B(n13), .C(\mem<18><2> ), .D(n699), .Y(
        n1731) );
  AOI22X1 U3393 ( .A(\mem<17><2> ), .B(n780), .C(\mem<16><2> ), .D(n1504), .Y(
        n1730) );
  AOI22X1 U3394 ( .A(\mem<23><2> ), .B(n813), .C(\mem<22><2> ), .D(n1435), .Y(
        n1733) );
  AOI22X1 U3395 ( .A(\mem<21><2> ), .B(n1517), .C(\mem<20><2> ), .D(n785), .Y(
        n1732) );
  NAND3X1 U3396 ( .A(n492), .B(n152), .C(n154), .Y(n1743) );
  NOR2X1 U3397 ( .A(n2475), .B(n4563), .Y(n1734) );
  AOI21X1 U3398 ( .A(\mem<1><2> ), .B(n807), .C(n1734), .Y(n1735) );
  NAND3X1 U3399 ( .A(n1735), .B(n1159), .C(n859), .Y(n1738) );
  AOI22X1 U3400 ( .A(\mem<7><2> ), .B(n35), .C(\mem<6><2> ), .D(n823), .Y(
        n1737) );
  AOI22X1 U3401 ( .A(\mem<5><2> ), .B(n689), .C(\mem<4><2> ), .D(n816), .Y(
        n1736) );
  AOI22X1 U3402 ( .A(\mem<11><2> ), .B(n847), .C(\mem<10><2> ), .D(n140), .Y(
        n1740) );
  AOI22X1 U3403 ( .A(\mem<9><2> ), .B(n1472), .C(\mem<8><2> ), .D(n57), .Y(
        n1739) );
  AOI22X1 U3404 ( .A(\mem<15><2> ), .B(n851), .C(\mem<14><2> ), .D(n801), .Y(
        n1742) );
  AOI22X1 U3405 ( .A(\mem<13><2> ), .B(n56), .C(\mem<12><2> ), .D(n1446), .Y(
        n1741) );
  AOI21X1 U3406 ( .A(n534), .B(n524), .C(n1173), .Y(\data_out<2> ) );
  AOI22X1 U3407 ( .A(\mem<35><3> ), .B(n777), .C(\mem<34><3> ), .D(n775), .Y(
        n1745) );
  AOI22X1 U3408 ( .A(\mem<33><3> ), .B(n3718), .C(\mem<32><3> ), .D(n788), .Y(
        n1744) );
  AOI22X1 U3409 ( .A(\mem<39><3> ), .B(n790), .C(\mem<38><3> ), .D(n783), .Y(
        n1747) );
  AOI22X1 U3410 ( .A(\mem<37><3> ), .B(n791), .C(\mem<36><3> ), .D(n84), .Y(
        n1746) );
  AOI22X1 U3411 ( .A(\mem<43><3> ), .B(n694), .C(\mem<42><3> ), .D(n860), .Y(
        n1749) );
  AOI22X1 U3412 ( .A(\mem<41><3> ), .B(n43), .C(\mem<40><3> ), .D(n1456), .Y(
        n1748) );
  AOI22X1 U3413 ( .A(\mem<47><3> ), .B(n695), .C(\mem<46><3> ), .D(n832), .Y(
        n1751) );
  AOI22X1 U3414 ( .A(\mem<45><3> ), .B(n8), .C(\mem<44><3> ), .D(n1466), .Y(
        n1750) );
  OAI21X1 U3415 ( .A(n634), .B(n1752), .C(n979), .Y(n1755) );
  OAI21X1 U3416 ( .A(n2980), .B(n1753), .C(n981), .Y(n1754) );
  NAND2X1 U3417 ( .A(\mem<56><3> ), .B(n3166), .Y(n1756) );
  OAI21X1 U3418 ( .A(n3141), .B(n1757), .C(n1756), .Y(n1760) );
  OAI21X1 U3419 ( .A(n3087), .B(n1758), .C(n983), .Y(n1759) );
  AOI22X1 U3420 ( .A(\mem<51><3> ), .B(n3296), .C(\mem<50><3> ), .D(n839), .Y(
        n1762) );
  AOI22X1 U3421 ( .A(\mem<49><3> ), .B(n795), .C(\mem<48><3> ), .D(n1500), .Y(
        n1761) );
  AOI22X1 U3422 ( .A(\mem<55><3> ), .B(n3167), .C(\mem<54><3> ), .D(n854), .Y(
        n1764) );
  AOI22X1 U3423 ( .A(\mem<53><3> ), .B(n698), .C(\mem<52><3> ), .D(n833), .Y(
        n1763) );
  NAND3X1 U3424 ( .A(n494), .B(n162), .C(n160), .Y(n1765) );
  OAI21X1 U3425 ( .A(n1482), .B(n1766), .C(n733), .Y(n1770) );
  NAND2X1 U3426 ( .A(\mem<31><3> ), .B(n3793), .Y(n1767) );
  OAI21X1 U3427 ( .A(n3795), .B(n1768), .C(n1767), .Y(n1769) );
  OAI21X1 U3428 ( .A(n802), .B(n1771), .C(n985), .Y(n1774) );
  OAI21X1 U3429 ( .A(n849), .B(n1772), .C(n325), .Y(n1773) );
  AOI22X1 U3430 ( .A(\mem<19><3> ), .B(n720), .C(\mem<18><3> ), .D(n699), .Y(
        n1776) );
  AOI22X1 U3431 ( .A(\mem<17><3> ), .B(n781), .C(\mem<16><3> ), .D(n1504), .Y(
        n1775) );
  AOI22X1 U3432 ( .A(\mem<23><3> ), .B(n813), .C(\mem<22><3> ), .D(n1435), .Y(
        n1778) );
  AOI22X1 U3433 ( .A(\mem<21><3> ), .B(n1517), .C(\mem<20><3> ), .D(n785), .Y(
        n1777) );
  NAND3X1 U3434 ( .A(n496), .B(n164), .C(n166), .Y(n1788) );
  NOR2X1 U3435 ( .A(n2475), .B(n4562), .Y(n1779) );
  AOI21X1 U3436 ( .A(\mem<1><3> ), .B(n808), .C(n1779), .Y(n1780) );
  NAND3X1 U3437 ( .A(n762), .B(n1161), .C(n1780), .Y(n1783) );
  AOI22X1 U3438 ( .A(\mem<7><3> ), .B(n35), .C(\mem<6><3> ), .D(n823), .Y(
        n1782) );
  AOI22X1 U3439 ( .A(\mem<5><3> ), .B(n689), .C(\mem<4><3> ), .D(n816), .Y(
        n1781) );
  AOI22X1 U3440 ( .A(\mem<11><3> ), .B(n847), .C(\mem<10><3> ), .D(n140), .Y(
        n1785) );
  AOI22X1 U3441 ( .A(\mem<9><3> ), .B(n1472), .C(\mem<8><3> ), .D(n829), .Y(
        n1784) );
  AOI22X1 U3442 ( .A(\mem<15><3> ), .B(n851), .C(\mem<14><3> ), .D(n801), .Y(
        n1787) );
  AOI22X1 U3443 ( .A(\mem<13><3> ), .B(n56), .C(\mem<12><3> ), .D(n1446), .Y(
        n1786) );
  AOI21X1 U3444 ( .A(n536), .B(n526), .C(n1173), .Y(\data_out<3> ) );
  AOI22X1 U3445 ( .A(\mem<35><4> ), .B(n778), .C(\mem<34><4> ), .D(n776), .Y(
        n1790) );
  AOI22X1 U3446 ( .A(\mem<33><4> ), .B(n3718), .C(\mem<32><4> ), .D(n788), .Y(
        n1789) );
  AOI22X1 U3447 ( .A(\mem<39><4> ), .B(n654), .C(\mem<38><4> ), .D(n783), .Y(
        n1792) );
  AOI22X1 U3448 ( .A(\mem<37><4> ), .B(n656), .C(\mem<36><4> ), .D(n85), .Y(
        n1791) );
  AOI22X1 U3449 ( .A(\mem<43><4> ), .B(n694), .C(\mem<42><4> ), .D(n860), .Y(
        n1794) );
  AOI22X1 U3450 ( .A(\mem<41><4> ), .B(n42), .C(\mem<40><4> ), .D(n1456), .Y(
        n1793) );
  AOI22X1 U3451 ( .A(\mem<47><4> ), .B(n695), .C(\mem<46><4> ), .D(n832), .Y(
        n1796) );
  AOI22X1 U3452 ( .A(\mem<45><4> ), .B(n661), .C(\mem<44><4> ), .D(n1466), .Y(
        n1795) );
  NAND2X1 U3453 ( .A(\mem<61><4> ), .B(n662), .Y(n1797) );
  OAI21X1 U3454 ( .A(n634), .B(n1798), .C(n1797), .Y(n1802) );
  NAND2X1 U3455 ( .A(\mem<63><4> ), .B(n2978), .Y(n1799) );
  OAI21X1 U3456 ( .A(n2980), .B(n1800), .C(n1799), .Y(n1801) );
  NAND2X1 U3457 ( .A(\mem<56><4> ), .B(n3166), .Y(n1803) );
  OAI21X1 U3458 ( .A(n3141), .B(n1804), .C(n1803), .Y(n1808) );
  NAND2X1 U3459 ( .A(\mem<59><4> ), .B(n522), .Y(n1805) );
  OAI21X1 U3460 ( .A(n3087), .B(n1806), .C(n1805), .Y(n1807) );
  AOI22X1 U3461 ( .A(\mem<51><4> ), .B(n3296), .C(\mem<50><4> ), .D(n839), .Y(
        n1810) );
  AOI22X1 U3462 ( .A(\mem<49><4> ), .B(n796), .C(\mem<48><4> ), .D(n835), .Y(
        n1809) );
  AOI22X1 U3463 ( .A(\mem<55><4> ), .B(n831), .C(\mem<54><4> ), .D(n854), .Y(
        n1812) );
  AOI22X1 U3464 ( .A(\mem<53><4> ), .B(n698), .C(\mem<52><4> ), .D(n833), .Y(
        n1811) );
  OAI21X1 U3465 ( .A(n1482), .B(n1813), .C(n735), .Y(n2329) );
  NAND2X1 U3466 ( .A(\mem<31><4> ), .B(n3793), .Y(n1814) );
  OAI21X1 U3467 ( .A(n3795), .B(n1815), .C(n1814), .Y(n2328) );
  OAI21X1 U3468 ( .A(n802), .B(n2330), .C(n987), .Y(n2333) );
  OAI21X1 U3469 ( .A(n849), .B(n2331), .C(n327), .Y(n2332) );
  AOI22X1 U3470 ( .A(\mem<19><4> ), .B(n720), .C(\mem<18><4> ), .D(n699), .Y(
        n2335) );
  AOI22X1 U3471 ( .A(\mem<17><4> ), .B(n781), .C(\mem<16><4> ), .D(n719), .Y(
        n2334) );
  AOI22X1 U3472 ( .A(\mem<23><4> ), .B(n813), .C(\mem<22><4> ), .D(n1435), .Y(
        n2337) );
  AOI22X1 U3473 ( .A(\mem<21><4> ), .B(n1517), .C(\mem<20><4> ), .D(n784), .Y(
        n2336) );
  NAND3X1 U3474 ( .A(n498), .B(n176), .C(n565), .Y(n2347) );
  NOR2X1 U3475 ( .A(n2475), .B(n4561), .Y(n2338) );
  AOI21X1 U3476 ( .A(\mem<1><4> ), .B(n808), .C(n2338), .Y(n2339) );
  NAND3X1 U3477 ( .A(n1087), .B(n1163), .C(n2339), .Y(n2342) );
  AOI22X1 U3478 ( .A(\mem<7><4> ), .B(n35), .C(\mem<6><4> ), .D(n823), .Y(
        n2341) );
  AOI22X1 U3479 ( .A(\mem<5><4> ), .B(n689), .C(\mem<4><4> ), .D(n816), .Y(
        n2340) );
  AOI22X1 U3480 ( .A(\mem<11><4> ), .B(n847), .C(\mem<10><4> ), .D(n140), .Y(
        n2344) );
  AOI22X1 U3481 ( .A(\mem<9><4> ), .B(n1472), .C(\mem<8><4> ), .D(n57), .Y(
        n2343) );
  AOI22X1 U3482 ( .A(\mem<15><4> ), .B(n851), .C(\mem<14><4> ), .D(n801), .Y(
        n2346) );
  AOI22X1 U3483 ( .A(\mem<13><4> ), .B(n56), .C(\mem<12><4> ), .D(n1446), .Y(
        n2345) );
  AOI21X1 U3484 ( .A(n174), .B(n528), .C(n1173), .Y(\data_out<4> ) );
  AOI22X1 U3485 ( .A(\mem<35><5> ), .B(n777), .C(\mem<34><5> ), .D(n775), .Y(
        n2349) );
  AOI22X1 U3486 ( .A(\mem<33><5> ), .B(n3718), .C(\mem<32><5> ), .D(n788), .Y(
        n2348) );
  AOI22X1 U3487 ( .A(\mem<39><5> ), .B(n790), .C(\mem<38><5> ), .D(n783), .Y(
        n2351) );
  AOI22X1 U3488 ( .A(\mem<37><5> ), .B(n791), .C(\mem<36><5> ), .D(n779), .Y(
        n2350) );
  AOI22X1 U3489 ( .A(\mem<43><5> ), .B(n694), .C(\mem<42><5> ), .D(n860), .Y(
        n2353) );
  AOI22X1 U3490 ( .A(\mem<41><5> ), .B(n42), .C(\mem<40><5> ), .D(n1456), .Y(
        n2352) );
  AOI22X1 U3491 ( .A(\mem<47><5> ), .B(n695), .C(\mem<46><5> ), .D(n832), .Y(
        n2355) );
  AOI22X1 U3492 ( .A(\mem<45><5> ), .B(n1459), .C(\mem<44><5> ), .D(n1466), 
        .Y(n2354) );
  OAI21X1 U3493 ( .A(n634), .B(n2356), .C(n989), .Y(n2359) );
  OAI21X1 U3494 ( .A(n2980), .B(n2357), .C(n991), .Y(n2358) );
  NAND2X1 U3495 ( .A(\mem<56><5> ), .B(n3166), .Y(n2360) );
  OAI21X1 U3496 ( .A(n3141), .B(n2361), .C(n2360), .Y(n2364) );
  OAI21X1 U3497 ( .A(n3087), .B(n2362), .C(n993), .Y(n2363) );
  AOI22X1 U3498 ( .A(\mem<51><5> ), .B(n3296), .C(\mem<50><5> ), .D(n840), .Y(
        n2366) );
  AOI22X1 U3499 ( .A(\mem<49><5> ), .B(n795), .C(\mem<48><5> ), .D(n835), .Y(
        n2365) );
  AOI22X1 U3500 ( .A(\mem<55><5> ), .B(n831), .C(\mem<54><5> ), .D(n854), .Y(
        n2368) );
  AOI22X1 U3501 ( .A(\mem<53><5> ), .B(n6), .C(\mem<52><5> ), .D(n833), .Y(
        n2367) );
  NAND3X1 U3502 ( .A(n182), .B(n184), .C(n567), .Y(n2369) );
  OAI21X1 U3503 ( .A(n1482), .B(n2370), .C(n737), .Y(n2374) );
  NAND2X1 U3504 ( .A(\mem<31><5> ), .B(n3793), .Y(n2371) );
  OAI21X1 U3505 ( .A(n3795), .B(n2372), .C(n2371), .Y(n2373) );
  OAI21X1 U3506 ( .A(n802), .B(n2375), .C(n995), .Y(n2379) );
  NAND2X1 U3507 ( .A(\mem<27><5> ), .B(n811), .Y(n2376) );
  OAI21X1 U3508 ( .A(n849), .B(n2377), .C(n2376), .Y(n2378) );
  AOI22X1 U3509 ( .A(\mem<19><5> ), .B(n13), .C(\mem<18><5> ), .D(n699), .Y(
        n2381) );
  AOI22X1 U3510 ( .A(\mem<17><5> ), .B(n780), .C(\mem<16><5> ), .D(n719), .Y(
        n2380) );
  AOI22X1 U3511 ( .A(\mem<23><5> ), .B(n813), .C(\mem<22><5> ), .D(n1435), .Y(
        n2383) );
  AOI22X1 U3512 ( .A(\mem<21><5> ), .B(n782), .C(\mem<20><5> ), .D(n784), .Y(
        n2382) );
  NAND3X1 U3513 ( .A(n500), .B(n186), .C(n188), .Y(n2392) );
  AOI21X1 U3514 ( .A(\mem<1><5> ), .B(n807), .C(n760), .Y(n2384) );
  NAND3X1 U3515 ( .A(n2384), .B(n1165), .C(n764), .Y(n2387) );
  AOI22X1 U3516 ( .A(\mem<7><5> ), .B(n35), .C(\mem<6><5> ), .D(n823), .Y(
        n2386) );
  AOI22X1 U3517 ( .A(\mem<5><5> ), .B(n689), .C(\mem<4><5> ), .D(n816), .Y(
        n2385) );
  AOI22X1 U3518 ( .A(\mem<11><5> ), .B(n847), .C(\mem<10><5> ), .D(n140), .Y(
        n2389) );
  AOI22X1 U3519 ( .A(\mem<9><5> ), .B(n1472), .C(\mem<8><5> ), .D(n57), .Y(
        n2388) );
  AOI22X1 U3520 ( .A(\mem<15><5> ), .B(n851), .C(\mem<14><5> ), .D(n801), .Y(
        n2391) );
  AOI22X1 U3521 ( .A(\mem<13><5> ), .B(n56), .C(\mem<12><5> ), .D(n1458), .Y(
        n2390) );
  AOI21X1 U3522 ( .A(n538), .B(n190), .C(n1173), .Y(\data_out<5> ) );
  AOI22X1 U3523 ( .A(\mem<35><6> ), .B(n778), .C(\mem<34><6> ), .D(n776), .Y(
        n2394) );
  AOI22X1 U3524 ( .A(\mem<33><6> ), .B(n3718), .C(\mem<32><6> ), .D(n788), .Y(
        n2393) );
  AOI22X1 U3525 ( .A(\mem<39><6> ), .B(n790), .C(\mem<38><6> ), .D(n783), .Y(
        n2396) );
  AOI22X1 U3526 ( .A(\mem<37><6> ), .B(n791), .C(\mem<36><6> ), .D(n779), .Y(
        n2395) );
  AOI22X1 U3527 ( .A(\mem<43><6> ), .B(n694), .C(\mem<42><6> ), .D(n860), .Y(
        n2398) );
  AOI22X1 U3528 ( .A(\mem<41><6> ), .B(n43), .C(\mem<40><6> ), .D(n1460), .Y(
        n2397) );
  AOI22X1 U3529 ( .A(\mem<47><6> ), .B(n695), .C(\mem<46><6> ), .D(n832), .Y(
        n2400) );
  AOI22X1 U3530 ( .A(\mem<45><6> ), .B(n1459), .C(\mem<44><6> ), .D(n1466), 
        .Y(n2399) );
  OAI21X1 U3531 ( .A(n634), .B(n2401), .C(n997), .Y(n2404) );
  OAI21X1 U3532 ( .A(n2980), .B(n2402), .C(n999), .Y(n2403) );
  OAI21X1 U3533 ( .A(n3141), .B(n2405), .C(n329), .Y(n2408) );
  OAI21X1 U3534 ( .A(n3087), .B(n2406), .C(n1001), .Y(n2407) );
  AOI22X1 U3535 ( .A(\mem<51><6> ), .B(n3296), .C(\mem<50><6> ), .D(n840), .Y(
        n2410) );
  AOI22X1 U3536 ( .A(\mem<49><6> ), .B(n821), .C(\mem<48><6> ), .D(n835), .Y(
        n2409) );
  AOI22X1 U3537 ( .A(\mem<55><6> ), .B(n831), .C(\mem<54><6> ), .D(n854), .Y(
        n2412) );
  AOI22X1 U3538 ( .A(\mem<53><6> ), .B(n6), .C(\mem<52><6> ), .D(n833), .Y(
        n2411) );
  NAND3X1 U3539 ( .A(n502), .B(n200), .C(n198), .Y(n2413) );
  OAI21X1 U3540 ( .A(n1482), .B(n2414), .C(n739), .Y(n2418) );
  NAND2X1 U3541 ( .A(\mem<31><6> ), .B(n3793), .Y(n2415) );
  OAI21X1 U3542 ( .A(n3795), .B(n2416), .C(n2415), .Y(n2417) );
  OAI21X1 U3543 ( .A(n802), .B(n2419), .C(n1003), .Y(n2423) );
  NAND2X1 U3544 ( .A(\mem<27><6> ), .B(n811), .Y(n2420) );
  OAI21X1 U3545 ( .A(n849), .B(n2421), .C(n2420), .Y(n2422) );
  AOI22X1 U3546 ( .A(\mem<19><6> ), .B(n13), .C(\mem<18><6> ), .D(n699), .Y(
        n2425) );
  AOI22X1 U3547 ( .A(\mem<17><6> ), .B(n781), .C(\mem<16><6> ), .D(n1504), .Y(
        n2424) );
  AOI22X1 U3548 ( .A(\mem<23><6> ), .B(n813), .C(\mem<22><6> ), .D(n1435), .Y(
        n2427) );
  AOI22X1 U3549 ( .A(\mem<21><6> ), .B(n782), .C(\mem<20><6> ), .D(n852), .Y(
        n2426) );
  NAND3X1 U3550 ( .A(n504), .B(n202), .C(n204), .Y(n2437) );
  NOR2X1 U3551 ( .A(n2475), .B(n4559), .Y(n2428) );
  AOI21X1 U3552 ( .A(\mem<1><6> ), .B(n1444), .C(n2428), .Y(n2429) );
  NAND3X1 U3553 ( .A(n2429), .B(n1167), .C(n1089), .Y(n2432) );
  AOI22X1 U3554 ( .A(\mem<7><6> ), .B(n35), .C(\mem<6><6> ), .D(n823), .Y(
        n2431) );
  AOI22X1 U3555 ( .A(\mem<5><6> ), .B(n1486), .C(\mem<4><6> ), .D(n816), .Y(
        n2430) );
  AOI22X1 U3556 ( .A(\mem<11><6> ), .B(n847), .C(\mem<10><6> ), .D(n140), .Y(
        n2434) );
  AOI22X1 U3557 ( .A(\mem<9><6> ), .B(n1472), .C(\mem<8><6> ), .D(n10), .Y(
        n2433) );
  AOI22X1 U3558 ( .A(\mem<15><6> ), .B(n851), .C(\mem<14><6> ), .D(n801), .Y(
        n2436) );
  AOI22X1 U3559 ( .A(\mem<13><6> ), .B(n26), .C(\mem<12><6> ), .D(n853), .Y(
        n2435) );
  AOI21X1 U3560 ( .A(n540), .B(n208), .C(n1173), .Y(\data_out<6> ) );
  AOI22X1 U3561 ( .A(\mem<35><7> ), .B(n778), .C(\mem<34><7> ), .D(n776), .Y(
        n2439) );
  AOI22X1 U3562 ( .A(\mem<33><7> ), .B(n3718), .C(\mem<32><7> ), .D(n788), .Y(
        n2438) );
  AOI22X1 U3563 ( .A(\mem<39><7> ), .B(n654), .C(\mem<38><7> ), .D(n783), .Y(
        n2441) );
  AOI22X1 U3564 ( .A(\mem<37><7> ), .B(n656), .C(\mem<36><7> ), .D(n84), .Y(
        n2440) );
  AOI22X1 U3565 ( .A(\mem<43><7> ), .B(n694), .C(\mem<42><7> ), .D(n860), .Y(
        n2443) );
  AOI22X1 U3566 ( .A(\mem<41><7> ), .B(n42), .C(\mem<40><7> ), .D(n1415), .Y(
        n2442) );
  AOI22X1 U3567 ( .A(\mem<47><7> ), .B(n695), .C(\mem<46><7> ), .D(n832), .Y(
        n2445) );
  AOI22X1 U3568 ( .A(\mem<45><7> ), .B(n8), .C(\mem<44><7> ), .D(n1466), .Y(
        n2444) );
  OAI21X1 U3569 ( .A(n634), .B(n2446), .C(n331), .Y(n2450) );
  NAND2X1 U3570 ( .A(\mem<63><7> ), .B(n2978), .Y(n2447) );
  OAI21X1 U3571 ( .A(n2980), .B(n2448), .C(n2447), .Y(n2449) );
  OAI21X1 U3572 ( .A(n3141), .B(n2451), .C(n333), .Y(n2455) );
  NAND2X1 U3573 ( .A(\mem<59><7> ), .B(n522), .Y(n2452) );
  OAI21X1 U3574 ( .A(n3087), .B(n2453), .C(n2452), .Y(n2454) );
  AOI22X1 U3575 ( .A(\mem<51><7> ), .B(n3296), .C(\mem<50><7> ), .D(n839), .Y(
        n2457) );
  AOI22X1 U3576 ( .A(\mem<49><7> ), .B(n795), .C(\mem<48><7> ), .D(n835), .Y(
        n2456) );
  AOI22X1 U3577 ( .A(\mem<55><7> ), .B(n831), .C(\mem<54><7> ), .D(n854), .Y(
        n2459) );
  AOI22X1 U3578 ( .A(\mem<53><7> ), .B(n6), .C(\mem<52><7> ), .D(n833), .Y(
        n2458) );
  NAND3X1 U3579 ( .A(n216), .B(n218), .C(n569), .Y(n2460) );
  OAI21X1 U3580 ( .A(n1482), .B(n2461), .C(n335), .Y(n2465) );
  NAND2X1 U3581 ( .A(\mem<31><7> ), .B(n3793), .Y(n2462) );
  OAI21X1 U3582 ( .A(n3795), .B(n2463), .C(n2462), .Y(n2464) );
  OAI21X1 U3583 ( .A(n803), .B(n2466), .C(n1005), .Y(n2470) );
  NAND2X1 U3584 ( .A(\mem<27><7> ), .B(n811), .Y(n2467) );
  OAI21X1 U3585 ( .A(n849), .B(n2468), .C(n2467), .Y(n2469) );
  AOI22X1 U3586 ( .A(\mem<19><7> ), .B(n720), .C(\mem<18><7> ), .D(n699), .Y(
        n2472) );
  AOI22X1 U3587 ( .A(\mem<17><7> ), .B(n780), .C(\mem<16><7> ), .D(n719), .Y(
        n2471) );
  AOI22X1 U3588 ( .A(\mem<23><7> ), .B(n813), .C(\mem<22><7> ), .D(n1435), .Y(
        n2474) );
  AOI22X1 U3589 ( .A(\mem<21><7> ), .B(n1517), .C(\mem<20><7> ), .D(n784), .Y(
        n2473) );
  NAND3X1 U3590 ( .A(n506), .B(n222), .C(n571), .Y(n2485) );
  NOR2X1 U3591 ( .A(n2475), .B(n4558), .Y(n2476) );
  AOI21X1 U3592 ( .A(\mem<1><7> ), .B(n808), .C(n2476), .Y(n2477) );
  NAND3X1 U3593 ( .A(n2477), .B(n1169), .C(n1091), .Y(n2480) );
  AOI22X1 U3594 ( .A(\mem<7><7> ), .B(n35), .C(\mem<6><7> ), .D(n823), .Y(
        n2479) );
  AOI22X1 U3595 ( .A(\mem<5><7> ), .B(n689), .C(\mem<4><7> ), .D(n816), .Y(
        n2478) );
  AOI22X1 U3596 ( .A(\mem<11><7> ), .B(n847), .C(\mem<10><7> ), .D(n140), .Y(
        n2482) );
  AOI22X1 U3597 ( .A(\mem<9><7> ), .B(n1472), .C(\mem<8><7> ), .D(n57), .Y(
        n2481) );
  AOI22X1 U3598 ( .A(\mem<15><7> ), .B(n851), .C(\mem<14><7> ), .D(n801), .Y(
        n2484) );
  AOI22X1 U3599 ( .A(\mem<13><7> ), .B(n56), .C(\mem<12><7> ), .D(n1446), .Y(
        n2483) );
  AOI21X1 U3600 ( .A(n542), .B(n530), .C(n1173), .Y(\data_out<7> ) );
  MUX2X1 U3601 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1542), .Y(n2487) );
  MUX2X1 U3602 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n33), .Y(n2486) );
  MUX2X1 U3603 ( .B(n2487), .A(n2486), .S(n1562), .Y(n2491) );
  MUX2X1 U3604 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1542), .Y(n2489) );
  MUX2X1 U3605 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n33), .Y(n2488) );
  MUX2X1 U3606 ( .B(n2489), .A(n2488), .S(n1561), .Y(n2490) );
  MUX2X1 U3607 ( .B(n2491), .A(n2490), .S(n1423), .Y(n2499) );
  MUX2X1 U3608 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n33), .Y(n2493) );
  MUX2X1 U3609 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n33), .Y(n2492) );
  MUX2X1 U3610 ( .B(n2493), .A(n2492), .S(n1562), .Y(n2497) );
  MUX2X1 U3611 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n33), .Y(n2495) );
  MUX2X1 U3612 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n33), .Y(n2494) );
  MUX2X1 U3613 ( .B(n2495), .A(n2494), .S(n1561), .Y(n2496) );
  MUX2X1 U3614 ( .B(n2497), .A(n2496), .S(n1423), .Y(n2498) );
  MUX2X1 U3615 ( .B(n2499), .A(n2498), .S(n1577), .Y(n2515) );
  MUX2X1 U3616 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1542), .Y(n2501) );
  MUX2X1 U3617 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n33), .Y(n2500) );
  MUX2X1 U3618 ( .B(n2501), .A(n2500), .S(n1561), .Y(n2505) );
  MUX2X1 U3619 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1543), .Y(n2503) );
  MUX2X1 U3620 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n33), .Y(n2502) );
  MUX2X1 U3621 ( .B(n2503), .A(n2502), .S(n1561), .Y(n2504) );
  MUX2X1 U3622 ( .B(n2505), .A(n2504), .S(n1571), .Y(n2513) );
  MUX2X1 U3623 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n33), .Y(n2507) );
  MUX2X1 U3624 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n33), .Y(n2506) );
  MUX2X1 U3625 ( .B(n2507), .A(n2506), .S(n1562), .Y(n2511) );
  MUX2X1 U3626 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1542), .Y(n2509) );
  MUX2X1 U3627 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1545), .Y(n2508) );
  MUX2X1 U3628 ( .B(n2509), .A(n2508), .S(n1561), .Y(n2510) );
  MUX2X1 U3629 ( .B(n2511), .A(n2510), .S(n1423), .Y(n2512) );
  MUX2X1 U3630 ( .B(n2513), .A(n2512), .S(n1577), .Y(n2514) );
  MUX2X1 U3631 ( .B(n2515), .A(n2514), .S(n830), .Y(n2547) );
  MUX2X1 U3632 ( .B(\mem<32><0> ), .A(\mem<33><0> ), .S(n33), .Y(n2517) );
  MUX2X1 U3633 ( .B(\mem<34><0> ), .A(\mem<35><0> ), .S(n1545), .Y(n2516) );
  MUX2X1 U3634 ( .B(n2517), .A(n2516), .S(n1563), .Y(n2521) );
  MUX2X1 U3635 ( .B(\mem<36><0> ), .A(\mem<37><0> ), .S(n33), .Y(n2519) );
  MUX2X1 U3636 ( .B(\mem<38><0> ), .A(\mem<39><0> ), .S(n33), .Y(n2518) );
  MUX2X1 U3637 ( .B(n2519), .A(n2518), .S(n1563), .Y(n2520) );
  MUX2X1 U3638 ( .B(n2521), .A(n2520), .S(n1571), .Y(n2529) );
  MUX2X1 U3639 ( .B(\mem<40><0> ), .A(\mem<41><0> ), .S(n1545), .Y(n2523) );
  MUX2X1 U3640 ( .B(\mem<42><0> ), .A(\mem<43><0> ), .S(n33), .Y(n2522) );
  MUX2X1 U3641 ( .B(n2523), .A(n2522), .S(n1563), .Y(n2527) );
  MUX2X1 U3642 ( .B(\mem<44><0> ), .A(\mem<45><0> ), .S(n1545), .Y(n2525) );
  MUX2X1 U3643 ( .B(\mem<46><0> ), .A(\mem<47><0> ), .S(n33), .Y(n2524) );
  MUX2X1 U3644 ( .B(n2525), .A(n2524), .S(n1563), .Y(n2526) );
  MUX2X1 U3645 ( .B(n2527), .A(n2526), .S(n1423), .Y(n2528) );
  MUX2X1 U3646 ( .B(n2529), .A(n2528), .S(n1577), .Y(n2545) );
  MUX2X1 U3647 ( .B(\mem<48><0> ), .A(\mem<49><0> ), .S(n33), .Y(n2531) );
  MUX2X1 U3648 ( .B(\mem<50><0> ), .A(\mem<51><0> ), .S(n1), .Y(n2530) );
  MUX2X1 U3649 ( .B(n2531), .A(n2530), .S(n1563), .Y(n2535) );
  MUX2X1 U3650 ( .B(\mem<52><0> ), .A(\mem<53><0> ), .S(n1543), .Y(n2533) );
  MUX2X1 U3651 ( .B(\mem<54><0> ), .A(\mem<55><0> ), .S(n1543), .Y(n2532) );
  MUX2X1 U3652 ( .B(n2533), .A(n2532), .S(n1563), .Y(n2534) );
  MUX2X1 U3653 ( .B(n2535), .A(n2534), .S(n1571), .Y(n2543) );
  MUX2X1 U3654 ( .B(\mem<56><0> ), .A(\mem<57><0> ), .S(n1), .Y(n2537) );
  MUX2X1 U3655 ( .B(\mem<58><0> ), .A(\mem<59><0> ), .S(n1), .Y(n2536) );
  MUX2X1 U3656 ( .B(n2537), .A(n2536), .S(n1563), .Y(n2541) );
  MUX2X1 U3657 ( .B(\mem<60><0> ), .A(\mem<61><0> ), .S(n1), .Y(n2539) );
  MUX2X1 U3658 ( .B(\mem<62><0> ), .A(\mem<63><0> ), .S(n1), .Y(n2538) );
  MUX2X1 U3659 ( .B(n2539), .A(n2538), .S(n1563), .Y(n2540) );
  MUX2X1 U3660 ( .B(n2541), .A(n2540), .S(n1571), .Y(n2542) );
  MUX2X1 U3661 ( .B(n2543), .A(n2542), .S(n1577), .Y(n2544) );
  MUX2X1 U3662 ( .B(n2545), .A(n2544), .S(n830), .Y(n2546) );
  MUX2X1 U3663 ( .B(n2547), .A(n2546), .S(n838), .Y(n2548) );
  AND2X2 U3664 ( .A(n1172), .B(n2548), .Y(\data_out<8> ) );
  MUX2X1 U3665 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1544), .Y(n2550) );
  MUX2X1 U3666 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1544), .Y(n2549) );
  MUX2X1 U3667 ( .B(n2550), .A(n2549), .S(n1563), .Y(n2554) );
  MUX2X1 U3668 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1544), .Y(n2552) );
  MUX2X1 U3669 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1544), .Y(n2551) );
  MUX2X1 U3670 ( .B(n2552), .A(n2551), .S(n1563), .Y(n2553) );
  MUX2X1 U3671 ( .B(n2554), .A(n2553), .S(n1571), .Y(n2562) );
  MUX2X1 U3672 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1544), .Y(n2556) );
  MUX2X1 U3673 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1484), .Y(n2555) );
  MUX2X1 U3674 ( .B(n2556), .A(n2555), .S(n1563), .Y(n2560) );
  MUX2X1 U3675 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1), .Y(n2558) );
  MUX2X1 U3676 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1), .Y(n2557) );
  MUX2X1 U3677 ( .B(n2558), .A(n2557), .S(n1563), .Y(n2559) );
  MUX2X1 U3678 ( .B(n2560), .A(n2559), .S(n1423), .Y(n2561) );
  MUX2X1 U3679 ( .B(n2562), .A(n2561), .S(n1577), .Y(n2578) );
  MUX2X1 U3680 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1484), .Y(n2564) );
  MUX2X1 U3681 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1), .Y(n2563) );
  MUX2X1 U3682 ( .B(n2564), .A(n2563), .S(n1562), .Y(n2568) );
  MUX2X1 U3683 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1544), .Y(n2566) );
  MUX2X1 U3684 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1544), .Y(n2565) );
  MUX2X1 U3685 ( .B(n2566), .A(n2565), .S(n1562), .Y(n2567) );
  MUX2X1 U3686 ( .B(n2568), .A(n2567), .S(n1423), .Y(n2576) );
  MUX2X1 U3687 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1), .Y(n2570) );
  MUX2X1 U3688 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1), .Y(n2569) );
  MUX2X1 U3689 ( .B(n2570), .A(n2569), .S(n1562), .Y(n2574) );
  MUX2X1 U3690 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1544), .Y(n2572) );
  MUX2X1 U3691 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1), .Y(n2571) );
  MUX2X1 U3692 ( .B(n2572), .A(n2571), .S(n1562), .Y(n2573) );
  MUX2X1 U3693 ( .B(n2574), .A(n2573), .S(n1423), .Y(n2575) );
  MUX2X1 U3694 ( .B(n2576), .A(n2575), .S(n1577), .Y(n2577) );
  MUX2X1 U3695 ( .B(n2578), .A(n2577), .S(n830), .Y(n2610) );
  MUX2X1 U3696 ( .B(\mem<32><1> ), .A(\mem<33><1> ), .S(n1), .Y(n2580) );
  MUX2X1 U3697 ( .B(\mem<34><1> ), .A(\mem<35><1> ), .S(n1), .Y(n2579) );
  MUX2X1 U3698 ( .B(n2580), .A(n2579), .S(n1562), .Y(n2584) );
  MUX2X1 U3699 ( .B(\mem<36><1> ), .A(\mem<37><1> ), .S(n1545), .Y(n2582) );
  MUX2X1 U3700 ( .B(\mem<38><1> ), .A(\mem<39><1> ), .S(n1545), .Y(n2581) );
  MUX2X1 U3701 ( .B(n2582), .A(n2581), .S(n1562), .Y(n2583) );
  MUX2X1 U3702 ( .B(n2584), .A(n2583), .S(n1571), .Y(n2592) );
  MUX2X1 U3703 ( .B(\mem<40><1> ), .A(\mem<41><1> ), .S(n1545), .Y(n2586) );
  MUX2X1 U3704 ( .B(\mem<42><1> ), .A(\mem<43><1> ), .S(n1545), .Y(n2585) );
  MUX2X1 U3705 ( .B(n2586), .A(n2585), .S(n1562), .Y(n2590) );
  MUX2X1 U3706 ( .B(\mem<44><1> ), .A(\mem<45><1> ), .S(n1545), .Y(n2588) );
  MUX2X1 U3707 ( .B(\mem<46><1> ), .A(\mem<47><1> ), .S(n1545), .Y(n2587) );
  MUX2X1 U3708 ( .B(n2588), .A(n2587), .S(n1562), .Y(n2589) );
  MUX2X1 U3709 ( .B(n2590), .A(n2589), .S(n1423), .Y(n2591) );
  MUX2X1 U3710 ( .B(n2592), .A(n2591), .S(n1577), .Y(n2608) );
  MUX2X1 U3711 ( .B(\mem<48><1> ), .A(\mem<49><1> ), .S(n1545), .Y(n2594) );
  MUX2X1 U3712 ( .B(\mem<50><1> ), .A(\mem<51><1> ), .S(n1545), .Y(n2593) );
  MUX2X1 U3713 ( .B(n2594), .A(n2593), .S(n1562), .Y(n2598) );
  MUX2X1 U3714 ( .B(\mem<52><1> ), .A(\mem<53><1> ), .S(n1545), .Y(n2596) );
  MUX2X1 U3715 ( .B(\mem<54><1> ), .A(\mem<55><1> ), .S(n1545), .Y(n2595) );
  MUX2X1 U3716 ( .B(n2596), .A(n2595), .S(n1562), .Y(n2597) );
  MUX2X1 U3717 ( .B(n2598), .A(n2597), .S(n1423), .Y(n2606) );
  MUX2X1 U3718 ( .B(\mem<56><1> ), .A(\mem<57><1> ), .S(n1545), .Y(n2600) );
  MUX2X1 U3719 ( .B(\mem<58><1> ), .A(\mem<59><1> ), .S(n1545), .Y(n2599) );
  MUX2X1 U3720 ( .B(n2600), .A(n2599), .S(n1562), .Y(n2604) );
  MUX2X1 U3721 ( .B(\mem<60><1> ), .A(\mem<61><1> ), .S(n33), .Y(n2602) );
  MUX2X1 U3722 ( .B(\mem<62><1> ), .A(\mem<63><1> ), .S(n1545), .Y(n2601) );
  MUX2X1 U3723 ( .B(n2602), .A(n2601), .S(n1562), .Y(n2603) );
  MUX2X1 U3724 ( .B(n2604), .A(n2603), .S(n1423), .Y(n2605) );
  MUX2X1 U3725 ( .B(n2606), .A(n2605), .S(n1577), .Y(n2607) );
  MUX2X1 U3726 ( .B(n2608), .A(n2607), .S(n830), .Y(n2609) );
  MUX2X1 U3727 ( .B(n2610), .A(n2609), .S(n838), .Y(n2611) );
  AND2X2 U3728 ( .A(n1172), .B(n2611), .Y(\data_out<9> ) );
  MUX2X1 U3729 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1542), .Y(n2613) );
  MUX2X1 U3730 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n33), .Y(n2612) );
  MUX2X1 U3731 ( .B(n2613), .A(n2612), .S(n1561), .Y(n2617) );
  MUX2X1 U3732 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1542), .Y(n2615) );
  MUX2X1 U3733 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1542), .Y(n2614) );
  MUX2X1 U3734 ( .B(n2615), .A(n2614), .S(n1561), .Y(n2616) );
  MUX2X1 U3735 ( .B(n2617), .A(n2616), .S(n1423), .Y(n2625) );
  MUX2X1 U3736 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n33), .Y(n2619) );
  MUX2X1 U3737 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n33), .Y(n2618) );
  MUX2X1 U3738 ( .B(n2619), .A(n2618), .S(n1561), .Y(n2623) );
  MUX2X1 U3739 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1542), .Y(n2621) );
  MUX2X1 U3740 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n33), .Y(n2620) );
  MUX2X1 U3741 ( .B(n2621), .A(n2620), .S(n1561), .Y(n2622) );
  MUX2X1 U3742 ( .B(n2623), .A(n2622), .S(n1423), .Y(n2624) );
  MUX2X1 U3743 ( .B(n2625), .A(n2624), .S(n1577), .Y(n2641) );
  MUX2X1 U3744 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1542), .Y(n2627) );
  MUX2X1 U3745 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1542), .Y(n2626) );
  MUX2X1 U3746 ( .B(n2627), .A(n2626), .S(n1561), .Y(n2631) );
  MUX2X1 U3747 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1542), .Y(n2629) );
  MUX2X1 U3748 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1542), .Y(n2628) );
  MUX2X1 U3749 ( .B(n2629), .A(n2628), .S(n1561), .Y(n2630) );
  MUX2X1 U3750 ( .B(n2631), .A(n2630), .S(n1423), .Y(n2639) );
  MUX2X1 U3751 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1542), .Y(n2633) );
  MUX2X1 U3752 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1542), .Y(n2632) );
  MUX2X1 U3753 ( .B(n2633), .A(n2632), .S(n1561), .Y(n2637) );
  MUX2X1 U3754 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1542), .Y(n2635) );
  MUX2X1 U3755 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1542), .Y(n2634) );
  MUX2X1 U3756 ( .B(n2635), .A(n2634), .S(n1561), .Y(n2636) );
  MUX2X1 U3757 ( .B(n2637), .A(n2636), .S(n1423), .Y(n2638) );
  MUX2X1 U3758 ( .B(n2639), .A(n2638), .S(n1577), .Y(n2640) );
  MUX2X1 U3759 ( .B(n2641), .A(n2640), .S(n830), .Y(n2673) );
  MUX2X1 U3760 ( .B(\mem<32><2> ), .A(\mem<33><2> ), .S(n1542), .Y(n2643) );
  MUX2X1 U3761 ( .B(\mem<34><2> ), .A(\mem<35><2> ), .S(n1542), .Y(n2642) );
  MUX2X1 U3762 ( .B(n2643), .A(n2642), .S(n1561), .Y(n2647) );
  MUX2X1 U3763 ( .B(\mem<36><2> ), .A(\mem<37><2> ), .S(n1542), .Y(n2645) );
  MUX2X1 U3764 ( .B(\mem<38><2> ), .A(\mem<39><2> ), .S(n1542), .Y(n2644) );
  MUX2X1 U3765 ( .B(n2645), .A(n2644), .S(n1561), .Y(n2646) );
  MUX2X1 U3766 ( .B(n2647), .A(n2646), .S(n1423), .Y(n2655) );
  MUX2X1 U3767 ( .B(\mem<40><2> ), .A(\mem<41><2> ), .S(n1542), .Y(n2649) );
  MUX2X1 U3768 ( .B(\mem<42><2> ), .A(\mem<43><2> ), .S(n1546), .Y(n2648) );
  MUX2X1 U3769 ( .B(n2649), .A(n2648), .S(n1561), .Y(n2653) );
  MUX2X1 U3770 ( .B(\mem<44><2> ), .A(\mem<45><2> ), .S(n1546), .Y(n2651) );
  MUX2X1 U3771 ( .B(\mem<46><2> ), .A(\mem<47><2> ), .S(n1546), .Y(n2650) );
  MUX2X1 U3772 ( .B(n2651), .A(n2650), .S(n1561), .Y(n2652) );
  MUX2X1 U3773 ( .B(n2653), .A(n2652), .S(n1423), .Y(n2654) );
  MUX2X1 U3774 ( .B(n2655), .A(n2654), .S(n1577), .Y(n2671) );
  MUX2X1 U3775 ( .B(\mem<48><2> ), .A(\mem<49><2> ), .S(n1546), .Y(n2657) );
  MUX2X1 U3776 ( .B(\mem<50><2> ), .A(\mem<51><2> ), .S(n1546), .Y(n2656) );
  MUX2X1 U3777 ( .B(n2657), .A(n2656), .S(n1560), .Y(n2661) );
  MUX2X1 U3778 ( .B(\mem<52><2> ), .A(\mem<53><2> ), .S(n1546), .Y(n2659) );
  MUX2X1 U3779 ( .B(\mem<54><2> ), .A(\mem<55><2> ), .S(n1546), .Y(n2658) );
  MUX2X1 U3780 ( .B(n2659), .A(n2658), .S(n1560), .Y(n2660) );
  MUX2X1 U3781 ( .B(n2661), .A(n2660), .S(n1423), .Y(n2669) );
  MUX2X1 U3782 ( .B(\mem<56><2> ), .A(\mem<57><2> ), .S(n1546), .Y(n2663) );
  MUX2X1 U3783 ( .B(\mem<58><2> ), .A(\mem<59><2> ), .S(n1546), .Y(n2662) );
  MUX2X1 U3784 ( .B(n2663), .A(n2662), .S(n1560), .Y(n2667) );
  MUX2X1 U3785 ( .B(\mem<60><2> ), .A(\mem<61><2> ), .S(n1546), .Y(n2665) );
  MUX2X1 U3786 ( .B(\mem<62><2> ), .A(\mem<63><2> ), .S(n1546), .Y(n2664) );
  MUX2X1 U3787 ( .B(n2665), .A(n2664), .S(n1560), .Y(n2666) );
  MUX2X1 U3788 ( .B(n2667), .A(n2666), .S(n1423), .Y(n2668) );
  MUX2X1 U3789 ( .B(n2669), .A(n2668), .S(n1577), .Y(n2670) );
  MUX2X1 U3790 ( .B(n2671), .A(n2670), .S(n830), .Y(n2672) );
  MUX2X1 U3791 ( .B(n2673), .A(n2672), .S(n838), .Y(n2674) );
  AND2X2 U3792 ( .A(n1172), .B(n2674), .Y(\data_out<10> ) );
  MUX2X1 U3793 ( .B(\mem<56><3> ), .A(\mem<57><3> ), .S(n1546), .Y(n2676) );
  MUX2X1 U3794 ( .B(\mem<58><3> ), .A(\mem<59><3> ), .S(n44), .Y(n2675) );
  MUX2X1 U3795 ( .B(n2676), .A(n2675), .S(n1560), .Y(n2680) );
  MUX2X1 U3796 ( .B(\mem<60><3> ), .A(\mem<61><3> ), .S(n1537), .Y(n2678) );
  MUX2X1 U3797 ( .B(\mem<62><3> ), .A(\mem<63><3> ), .S(n1537), .Y(n2677) );
  MUX2X1 U3798 ( .B(n2678), .A(n2677), .S(n1560), .Y(n2679) );
  MUX2X1 U3799 ( .B(n2680), .A(n2679), .S(n1423), .Y(n2681) );
  NAND3X1 U3800 ( .A(n2681), .B(n1429), .C(n1578), .Y(n2705) );
  MUX2X1 U3801 ( .B(\mem<48><3> ), .A(\mem<49><3> ), .S(n1537), .Y(n2683) );
  MUX2X1 U3802 ( .B(\mem<50><3> ), .A(\mem<51><3> ), .S(n48), .Y(n2682) );
  MUX2X1 U3803 ( .B(n2683), .A(n2682), .S(n1560), .Y(n2687) );
  MUX2X1 U3804 ( .B(\mem<52><3> ), .A(\mem<53><3> ), .S(n1544), .Y(n2685) );
  MUX2X1 U3805 ( .B(\mem<54><3> ), .A(\mem<55><3> ), .S(n1485), .Y(n2684) );
  MUX2X1 U3806 ( .B(n2685), .A(n2684), .S(n1560), .Y(n2686) );
  MUX2X1 U3807 ( .B(n2687), .A(n2686), .S(n1570), .Y(n2696) );
  MUX2X1 U3808 ( .B(\mem<40><3> ), .A(\mem<41><3> ), .S(n1546), .Y(n2690) );
  MUX2X1 U3809 ( .B(\mem<42><3> ), .A(\mem<43><3> ), .S(n1546), .Y(n2689) );
  MUX2X1 U3810 ( .B(n2690), .A(n2689), .S(n1560), .Y(n2694) );
  MUX2X1 U3811 ( .B(\mem<44><3> ), .A(\mem<45><3> ), .S(n1545), .Y(n2692) );
  MUX2X1 U3812 ( .B(\mem<46><3> ), .A(\mem<47><3> ), .S(n1453), .Y(n2691) );
  MUX2X1 U3813 ( .B(n2692), .A(n2691), .S(n1560), .Y(n2693) );
  MUX2X1 U3814 ( .B(n2694), .A(n2693), .S(n1570), .Y(n2695) );
  AOI22X1 U3815 ( .A(n767), .B(n2696), .C(n721), .D(n2695), .Y(n2704) );
  MUX2X1 U3816 ( .B(\mem<32><3> ), .A(\mem<33><3> ), .S(n1546), .Y(n2697) );
  MUX2X1 U3817 ( .B(n2697), .A(n133), .S(n1560), .Y(n2701) );
  MUX2X1 U3818 ( .B(\mem<36><3> ), .A(\mem<37><3> ), .S(n1546), .Y(n2699) );
  MUX2X1 U3819 ( .B(\mem<38><3> ), .A(\mem<39><3> ), .S(n1539), .Y(n2698) );
  MUX2X1 U3820 ( .B(n2699), .A(n2698), .S(n1560), .Y(n2700) );
  MUX2X1 U3821 ( .B(n2701), .A(n2700), .S(n1570), .Y(n2702) );
  AOI21X1 U3822 ( .A(n2702), .B(n722), .C(n1173), .Y(n2703) );
  MUX2X1 U3823 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1485), .Y(n2707) );
  MUX2X1 U3824 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n48), .Y(n2706) );
  MUX2X1 U3825 ( .B(n2707), .A(n2706), .S(n1559), .Y(n2711) );
  MUX2X1 U3826 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1543), .Y(n2709) );
  MUX2X1 U3827 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1485), .Y(n2708) );
  MUX2X1 U3828 ( .B(n2709), .A(n2708), .S(n1559), .Y(n2710) );
  MUX2X1 U3829 ( .B(n2711), .A(n2710), .S(n1570), .Y(n2713) );
  OR2X2 U3830 ( .A(N182), .B(N181), .Y(n2712) );
  NAND3X1 U3831 ( .A(n2713), .B(n2767), .C(n1428), .Y(n2722) );
  MUX2X1 U3832 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1544), .Y(n2715) );
  MUX2X1 U3833 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n48), .Y(n2714) );
  MUX2X1 U3834 ( .B(n2715), .A(n2714), .S(n1559), .Y(n2719) );
  MUX2X1 U3835 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1454), .Y(n2717) );
  MUX2X1 U3836 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1544), .Y(n2716) );
  MUX2X1 U3837 ( .B(n2719), .A(n2718), .S(n1570), .Y(n2720) );
  NAND3X1 U3838 ( .A(n2720), .B(n2767), .C(n1578), .Y(n2721) );
  MUX2X1 U3839 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n33), .Y(n2724) );
  MUX2X1 U3840 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1542), .Y(n2723) );
  MUX2X1 U3841 ( .B(n2724), .A(n2723), .S(n1559), .Y(n2728) );
  MUX2X1 U3842 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1485), .Y(n2726) );
  MUX2X1 U3843 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1454), .Y(n2725) );
  MUX2X1 U3844 ( .B(n2726), .A(n2725), .S(n1559), .Y(n2727) );
  MUX2X1 U3845 ( .B(n2728), .A(n2727), .S(n1570), .Y(n2729) );
  NAND3X1 U3846 ( .A(n2729), .B(n765), .C(n1578), .Y(n2738) );
  MUX2X1 U3847 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1542), .Y(n2731) );
  MUX2X1 U3848 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1537), .Y(n2730) );
  MUX2X1 U3849 ( .B(n2731), .A(n2730), .S(n1559), .Y(n2735) );
  MUX2X1 U3850 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1545), .Y(n2733) );
  MUX2X1 U3851 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1544), .Y(n2732) );
  MUX2X1 U3852 ( .B(n2733), .A(n2732), .S(n1559), .Y(n2734) );
  NAND3X1 U3853 ( .A(n1428), .B(n765), .C(n2736), .Y(n2737) );
  NOR3X1 U3854 ( .A(n577), .B(n579), .C(n120), .Y(\data_out<11> ) );
  MUX2X1 U3855 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1536), .Y(n2741) );
  MUX2X1 U3856 ( .B(n2742), .A(n2741), .S(n1559), .Y(n2743) );
  MUX2X1 U3857 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1542), .Y(n2747) );
  MUX2X1 U3858 ( .B(n2747), .A(n2746), .S(n1559), .Y(n2751) );
  MUX2X1 U3859 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1536), .Y(n2748) );
  MUX2X1 U3860 ( .B(n2749), .A(n2748), .S(n1558), .Y(n2750) );
  MUX2X1 U3861 ( .B(n2751), .A(n2750), .S(n1570), .Y(n2752) );
  MUX2X1 U3862 ( .B(\mem<34><4> ), .A(\mem<35><4> ), .S(n1538), .Y(n2753) );
  MUX2X1 U3863 ( .B(\mem<36><4> ), .A(\mem<37><4> ), .S(n1538), .Y(n2756) );
  MUX2X1 U3864 ( .B(n2756), .A(n2755), .S(n1558), .Y(n2757) );
  MUX2X1 U3865 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1537), .Y(n2761) );
  MUX2X1 U3866 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1537), .Y(n2760) );
  MUX2X1 U3867 ( .B(n2761), .A(n2760), .S(n1558), .Y(n2765) );
  MUX2X1 U3868 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1537), .Y(n2763) );
  MUX2X1 U3869 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n44), .Y(n2762) );
  MUX2X1 U3870 ( .B(n2763), .A(n2762), .S(n1558), .Y(n2764) );
  MUX2X1 U3871 ( .B(n2765), .A(n2764), .S(n1570), .Y(n2766) );
  MUX2X1 U3872 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1544), .Y(n2768) );
  MUX2X1 U3873 ( .B(n2769), .A(n2768), .S(n1558), .Y(n2773) );
  MUX2X1 U3874 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1537), .Y(n2771) );
  MUX2X1 U3875 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1545), .Y(n2770) );
  MUX2X1 U3876 ( .B(n2771), .A(n2770), .S(n1558), .Y(n2772) );
  NOR2X1 U3877 ( .A(n1280), .B(n1575), .Y(n2782) );
  MUX2X1 U3878 ( .B(\mem<44><4> ), .A(\mem<45><4> ), .S(n1537), .Y(n2776) );
  MUX2X1 U3879 ( .B(\mem<46><4> ), .A(\mem<47><4> ), .S(n1536), .Y(n2775) );
  MUX2X1 U3880 ( .B(n2776), .A(n2775), .S(n1558), .Y(n2777) );
  AOI21X1 U3881 ( .A(n2782), .B(n2781), .C(n233), .Y(n2800) );
  NOR2X1 U3882 ( .A(n242), .B(n1575), .Y(n2790) );
  MUX2X1 U3883 ( .B(\mem<52><4> ), .A(\mem<53><4> ), .S(n1545), .Y(n2784) );
  MUX2X1 U3884 ( .B(\mem<54><4> ), .A(\mem<55><4> ), .S(n1545), .Y(n2783) );
  NOR2X1 U3885 ( .A(n1280), .B(n1423), .Y(n2789) );
  MUX2X1 U3886 ( .B(\mem<40><4> ), .A(\mem<41><4> ), .S(n48), .Y(n2786) );
  MUX2X1 U3887 ( .B(\mem<42><4> ), .A(\mem<43><4> ), .S(n1546), .Y(n2785) );
  MUX2X1 U3888 ( .B(n2786), .A(n2785), .S(n1558), .Y(n2787) );
  AOI22X1 U3889 ( .A(n2790), .B(n127), .C(n2789), .D(n2788), .Y(n2799) );
  MUX2X1 U3890 ( .B(n2792), .A(n2791), .S(n1558), .Y(n2794) );
  NAND2X1 U3891 ( .A(n1576), .B(n768), .Y(n2793) );
  NOR3X1 U3892 ( .A(n1173), .B(n583), .C(n235), .Y(n2798) );
  NOR3X1 U3893 ( .A(n118), .B(n581), .C(n122), .Y(\data_out<12> ) );
  MUX2X1 U3894 ( .B(n2803), .A(n2802), .S(n1557), .Y(n2804) );
  MUX2X1 U3895 ( .B(n2805), .A(n2804), .S(n1570), .Y(n2806) );
  MUX2X1 U3896 ( .B(n2807), .A(n132), .S(n1557), .Y(n2811) );
  MUX2X1 U3897 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1544), .Y(n2809) );
  MUX2X1 U3898 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1544), .Y(n2808) );
  MUX2X1 U3899 ( .B(n2809), .A(n2808), .S(n1557), .Y(n2810) );
  MUX2X1 U3900 ( .B(n2811), .A(n2810), .S(n1570), .Y(n2812) );
  MUX2X1 U3901 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1541), .Y(n2814) );
  NAND2X1 U3902 ( .A(n1571), .B(n2815), .Y(n2819) );
  MUX2X1 U3903 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1547), .Y(n2817) );
  MUX2X1 U3904 ( .B(n2817), .A(n2816), .S(n1557), .Y(n2818) );
  MUX2X1 U3905 ( .B(n2821), .A(n2820), .S(n1557), .Y(n2822) );
  NAND2X1 U3906 ( .A(n1575), .B(n2825), .Y(n2826) );
  MUX2X1 U3907 ( .B(n2828), .A(n2827), .S(n1557), .Y(n2829) );
  MUX2X1 U3908 ( .B(\mem<34><5> ), .A(\mem<35><5> ), .S(n1539), .Y(n2830) );
  MUX2X1 U3909 ( .B(n2831), .A(n2830), .S(n1557), .Y(n2832) );
  NAND3X1 U3910 ( .A(n106), .B(n111), .C(n116), .Y(n2833) );
  MUX2X1 U3911 ( .B(\mem<58><5> ), .A(\mem<59><5> ), .S(n1539), .Y(n2834) );
  MUX2X1 U3912 ( .B(n2835), .A(n2834), .S(n1557), .Y(n2836) );
  NAND2X1 U3913 ( .A(n2836), .B(n1575), .Y(n2841) );
  MUX2X1 U3914 ( .B(\mem<60><5> ), .A(\mem<61><5> ), .S(n1485), .Y(n2838) );
  MUX2X1 U3915 ( .B(n2838), .A(n2837), .S(n1556), .Y(n2839) );
  NAND2X1 U3916 ( .A(n2839), .B(n1571), .Y(n2840) );
  MUX2X1 U3917 ( .B(\mem<54><5> ), .A(\mem<55><5> ), .S(n1485), .Y(n2842) );
  MUX2X1 U3918 ( .B(\mem<48><5> ), .A(\mem<49><5> ), .S(n44), .Y(n2846) );
  MUX2X1 U3919 ( .B(\mem<50><5> ), .A(\mem<51><5> ), .S(n1544), .Y(n2845) );
  MUX2X1 U3920 ( .B(n2846), .A(n2845), .S(n1561), .Y(n2847) );
  NAND2X1 U3921 ( .A(n1575), .B(n2847), .Y(n2848) );
  NAND3X1 U3922 ( .A(n508), .B(n767), .C(n2848), .Y(n2857) );
  MUX2X1 U3923 ( .B(n2850), .A(n2849), .S(n1560), .Y(n2851) );
  MUX2X1 U3924 ( .B(\mem<42><5> ), .A(\mem<43><5> ), .S(n1539), .Y(n2852) );
  MUX2X1 U3925 ( .B(n2853), .A(n2852), .S(n1561), .Y(n2854) );
  NAND2X1 U3926 ( .A(n1575), .B(n2854), .Y(n2855) );
  NAND3X1 U3927 ( .A(n2855), .B(n510), .C(n721), .Y(n2856) );
  AND2X2 U3928 ( .A(n281), .B(n313), .Y(\data_out<13> ) );
  MUX2X1 U3929 ( .B(\mem<56><6> ), .A(\mem<57><6> ), .S(n1544), .Y(n2865) );
  MUX2X1 U3930 ( .B(\mem<62><6> ), .A(\mem<63><6> ), .S(n44), .Y(n2866) );
  AOI22X1 U3931 ( .A(n725), .B(n2871), .C(n768), .D(n2870), .Y(n2887) );
  MUX2X1 U3932 ( .B(n2873), .A(n2872), .S(n1562), .Y(n2877) );
  MUX2X1 U3933 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1453), .Y(n2874) );
  MUX2X1 U3934 ( .B(n2875), .A(n2874), .S(n1561), .Y(n2876) );
  MUX2X1 U3935 ( .B(n2879), .A(n2878), .S(n1561), .Y(n2883) );
  MUX2X1 U3936 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1536), .Y(n2881) );
  MUX2X1 U3937 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1544), .Y(n2880) );
  MUX2X1 U3938 ( .B(n2881), .A(n2880), .S(n1556), .Y(n2882) );
  MUX2X1 U3939 ( .B(n2883), .A(n2882), .S(n1570), .Y(n2884) );
  AOI22X1 U3940 ( .A(n231), .B(n2885), .C(n724), .D(n2884), .Y(n2886) );
  NAND3X1 U3941 ( .A(n1172), .B(n543), .C(n556), .Y(n2918) );
  MUX2X1 U3942 ( .B(n2889), .A(n2888), .S(n1556), .Y(n2893) );
  MUX2X1 U3943 ( .B(\mem<44><6> ), .A(\mem<45><6> ), .S(n1542), .Y(n2891) );
  MUX2X1 U3944 ( .B(\mem<46><6> ), .A(\mem<47><6> ), .S(n1540), .Y(n2890) );
  MUX2X1 U3945 ( .B(n2891), .A(n2890), .S(n1556), .Y(n2892) );
  MUX2X1 U3946 ( .B(\mem<48><6> ), .A(\mem<49><6> ), .S(n1544), .Y(n2895) );
  MUX2X1 U3947 ( .B(\mem<50><6> ), .A(\mem<51><6> ), .S(n1544), .Y(n2894) );
  MUX2X1 U3948 ( .B(n2895), .A(n2894), .S(n1556), .Y(n2899) );
  MUX2X1 U3949 ( .B(\mem<52><6> ), .A(\mem<53><6> ), .S(n1539), .Y(n2897) );
  MUX2X1 U3950 ( .B(\mem<54><6> ), .A(\mem<55><6> ), .S(n1546), .Y(n2896) );
  MUX2X1 U3951 ( .B(n2897), .A(n2896), .S(n1556), .Y(n2898) );
  AOI22X1 U3952 ( .A(n721), .B(n2901), .C(n767), .D(n2900), .Y(n2917) );
  MUX2X1 U3953 ( .B(\mem<34><6> ), .A(\mem<35><6> ), .S(n1544), .Y(n2902) );
  MUX2X1 U3954 ( .B(n2903), .A(n2902), .S(n1556), .Y(n2907) );
  MUX2X1 U3955 ( .B(n2905), .A(n2904), .S(n1556), .Y(n2906) );
  MUX2X1 U3956 ( .B(n2909), .A(n2908), .S(n1556), .Y(n2913) );
  MUX2X1 U3957 ( .B(n2911), .A(n2910), .S(n1556), .Y(n2912) );
  MUX2X1 U3958 ( .B(n2913), .A(n2912), .S(n1570), .Y(n2914) );
  MUX2X1 U3959 ( .B(n2922), .A(n2921), .S(n1556), .Y(n2923) );
  MUX2X1 U3960 ( .B(n2924), .A(n2923), .S(n1570), .Y(n2925) );
  MUX2X1 U3961 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1454), .Y(n2927) );
  MUX2X1 U3962 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1454), .Y(n2926) );
  MUX2X1 U3963 ( .B(n2927), .A(n2926), .S(n1556), .Y(n2931) );
  MUX2X1 U3964 ( .B(n2929), .A(n2928), .S(n1555), .Y(n2930) );
  MUX2X1 U3965 ( .B(\mem<36><7> ), .A(\mem<37><7> ), .S(n1452), .Y(n2934) );
  MUX2X1 U3966 ( .B(n2936), .A(n2935), .S(n1555), .Y(n2937) );
  NAND3X1 U3967 ( .A(n722), .B(n553), .C(n573), .Y(n2954) );
  MUX2X1 U3968 ( .B(n2939), .A(n2938), .S(n1555), .Y(n2940) );
  NAND2X1 U3969 ( .A(n2940), .B(n1571), .Y(n2945) );
  MUX2X1 U3970 ( .B(n2942), .A(n2941), .S(n1555), .Y(n2943) );
  NAND2X1 U3971 ( .A(n2943), .B(n1575), .Y(n2944) );
  MUX2X1 U3972 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1485), .Y(n2946) );
  MUX2X1 U3973 ( .B(n2947), .A(n2946), .S(n1555), .Y(n2948) );
  NAND2X1 U3974 ( .A(n2948), .B(n1571), .Y(n2953) );
  NAND2X1 U3975 ( .A(n2951), .B(n1575), .Y(n2952) );
  MUX2X1 U3976 ( .B(\mem<62><7> ), .A(\mem<63><7> ), .S(n1537), .Y(n2956) );
  MUX2X1 U3977 ( .B(n2957), .A(n2956), .S(n1555), .Y(n2958) );
  MUX2X1 U3978 ( .B(\mem<58><7> ), .A(\mem<59><7> ), .S(n1538), .Y(n2959) );
  MUX2X1 U3979 ( .B(n2960), .A(n2959), .S(n1555), .Y(n2961) );
  NAND3X1 U3980 ( .A(n768), .B(n555), .C(n575), .Y(n2962) );
  MUX2X1 U3981 ( .B(\mem<54><7> ), .A(\mem<55><7> ), .S(n1539), .Y(n2963) );
  MUX2X1 U3982 ( .B(n2964), .A(n2963), .S(n1555), .Y(n2965) );
  MUX2X1 U3983 ( .B(n2967), .A(n2966), .S(n1555), .Y(n2968) );
  NAND2X1 U3984 ( .A(n1571), .B(n131), .Y(n2974) );
  AND2X2 U3985 ( .A(n285), .B(n317), .Y(\data_out<15> ) );
  OAI21X1 U3986 ( .A(n592), .B(n1279), .C(n1270), .Y(n2976) );
  AOI22X1 U3987 ( .A(\data_in<15> ), .B(n1094), .C(\data_in<7> ), .D(n1095), 
        .Y(n608) );
  AOI22X1 U3988 ( .A(\data_in<14> ), .B(n1094), .C(\data_in<6> ), .D(n1095), 
        .Y(n607) );
  AOI22X1 U3989 ( .A(\data_in<13> ), .B(n1094), .C(\data_in<5> ), .D(n1095), 
        .Y(n606) );
  AOI22X1 U3990 ( .A(\data_in<12> ), .B(n1094), .C(\data_in<4> ), .D(n1095), 
        .Y(n605) );
  AOI22X1 U3991 ( .A(\data_in<11> ), .B(n1094), .C(\data_in<3> ), .D(n1095), 
        .Y(n604) );
  AOI22X1 U3992 ( .A(\data_in<10> ), .B(n1094), .C(\data_in<2> ), .D(n1095), 
        .Y(n603) );
  AOI22X1 U3993 ( .A(\data_in<9> ), .B(n1094), .C(\data_in<1> ), .D(n1095), 
        .Y(n602) );
  AOI22X1 U3994 ( .A(\data_in<8> ), .B(n1094), .C(\data_in<0> ), .D(n1095), 
        .Y(n599) );
  INVX2 U3995 ( .A(n1282), .Y(n4496) );
  OAI21X1 U3996 ( .A(n2978), .B(n3006), .C(n4496), .Y(n3002) );
  AOI22X1 U3997 ( .A(\data_in<8> ), .B(n1096), .C(n2981), .D(n3002), .Y(n2982)
         );
  OAI21X1 U3998 ( .A(n1291), .B(n2983), .C(n2982), .Y(n1824) );
  AOI22X1 U3999 ( .A(\data_in<9> ), .B(n1096), .C(n2984), .D(n3002), .Y(n2985)
         );
  OAI21X1 U4000 ( .A(n1291), .B(n2986), .C(n2985), .Y(n1825) );
  AOI22X1 U4001 ( .A(\data_in<10> ), .B(n1096), .C(n2987), .D(n3002), .Y(n2988) );
  OAI21X1 U4002 ( .A(n1291), .B(n2989), .C(n2988), .Y(n1826) );
  AOI22X1 U4003 ( .A(\data_in<11> ), .B(n1096), .C(n2990), .D(n3002), .Y(n2991) );
  OAI21X1 U4004 ( .A(n1291), .B(n2992), .C(n2991), .Y(n1827) );
  AOI22X1 U4005 ( .A(\data_in<12> ), .B(n1096), .C(n2993), .D(n3002), .Y(n2994) );
  OAI21X1 U4006 ( .A(n1291), .B(n2995), .C(n2994), .Y(n1828) );
  AOI22X1 U4007 ( .A(\data_in<13> ), .B(n1096), .C(n2996), .D(n3002), .Y(n2997) );
  OAI21X1 U4008 ( .A(n1291), .B(n2998), .C(n2997), .Y(n1829) );
  AOI22X1 U4009 ( .A(\data_in<14> ), .B(n1096), .C(n2999), .D(n3002), .Y(n3000) );
  OAI21X1 U4010 ( .A(n1291), .B(n3001), .C(n3000), .Y(n1830) );
  AOI22X1 U4011 ( .A(\data_in<15> ), .B(n1096), .C(n3003), .D(n3002), .Y(n3004) );
  OAI21X1 U4012 ( .A(n1291), .B(n3005), .C(n3004), .Y(n1831) );
  OAI21X1 U4013 ( .A(n827), .B(n3006), .C(n4496), .Y(n3029) );
  AOI22X1 U4014 ( .A(\data_in<8> ), .B(n1097), .C(n3008), .D(n3029), .Y(n3009)
         );
  OAI21X1 U4015 ( .A(n1293), .B(n3010), .C(n3009), .Y(n1832) );
  AOI22X1 U4016 ( .A(\data_in<9> ), .B(n1097), .C(n3011), .D(n3029), .Y(n3012)
         );
  OAI21X1 U4017 ( .A(n1293), .B(n3013), .C(n3012), .Y(n1833) );
  AOI22X1 U4018 ( .A(\data_in<10> ), .B(n1097), .C(n3014), .D(n3029), .Y(n3015) );
  OAI21X1 U4019 ( .A(n1293), .B(n3016), .C(n3015), .Y(n1834) );
  AOI22X1 U4020 ( .A(\data_in<11> ), .B(n1097), .C(n3017), .D(n3029), .Y(n3018) );
  OAI21X1 U4021 ( .A(n1293), .B(n3019), .C(n3018), .Y(n1835) );
  AOI22X1 U4022 ( .A(\data_in<12> ), .B(n1097), .C(n3020), .D(n3029), .Y(n3021) );
  OAI21X1 U4023 ( .A(n1293), .B(n3022), .C(n3021), .Y(n1836) );
  AOI22X1 U4024 ( .A(\data_in<13> ), .B(n1097), .C(n3023), .D(n3029), .Y(n3024) );
  OAI21X1 U4025 ( .A(n1293), .B(n3025), .C(n3024), .Y(n1837) );
  AOI22X1 U4026 ( .A(\data_in<14> ), .B(n1097), .C(n3026), .D(n3029), .Y(n3027) );
  OAI21X1 U4027 ( .A(n1293), .B(n3028), .C(n3027), .Y(n1838) );
  AOI22X1 U4028 ( .A(\data_in<15> ), .B(n1097), .C(n3030), .D(n3029), .Y(n3031) );
  OAI21X1 U4029 ( .A(n1293), .B(n3032), .C(n3031), .Y(n1839) );
  OAI21X1 U4030 ( .A(n827), .B(n3059), .C(n4496), .Y(n3055) );
  AOI22X1 U4031 ( .A(\data_in<8> ), .B(n1098), .C(n3034), .D(n3055), .Y(n3035)
         );
  OAI21X1 U4032 ( .A(n1295), .B(n3036), .C(n3035), .Y(n1840) );
  AOI22X1 U4033 ( .A(\data_in<9> ), .B(n1098), .C(n3037), .D(n3055), .Y(n3038)
         );
  OAI21X1 U4034 ( .A(n1295), .B(n3039), .C(n3038), .Y(n1841) );
  AOI22X1 U4035 ( .A(\data_in<10> ), .B(n1098), .C(n3040), .D(n3055), .Y(n3041) );
  OAI21X1 U4036 ( .A(n1295), .B(n3042), .C(n3041), .Y(n1842) );
  AOI22X1 U4037 ( .A(\data_in<11> ), .B(n1098), .C(n3043), .D(n3055), .Y(n3044) );
  OAI21X1 U4038 ( .A(n1295), .B(n3045), .C(n3044), .Y(n1843) );
  AOI22X1 U4039 ( .A(\data_in<12> ), .B(n1098), .C(n3046), .D(n3055), .Y(n3047) );
  OAI21X1 U4040 ( .A(n1295), .B(n3048), .C(n3047), .Y(n1844) );
  AOI22X1 U4041 ( .A(\data_in<13> ), .B(n1098), .C(n3049), .D(n3055), .Y(n3050) );
  OAI21X1 U4042 ( .A(n1295), .B(n3051), .C(n3050), .Y(n1845) );
  AOI22X1 U4043 ( .A(\data_in<14> ), .B(n1098), .C(n3052), .D(n3055), .Y(n3053) );
  OAI21X1 U4044 ( .A(n1295), .B(n3054), .C(n3053), .Y(n1846) );
  AOI22X1 U4045 ( .A(\data_in<15> ), .B(n1098), .C(n3056), .D(n3055), .Y(n3057) );
  OAI21X1 U4046 ( .A(n1295), .B(n3058), .C(n3057), .Y(n1847) );
  OAI21X1 U4047 ( .A(n794), .B(n3059), .C(n4496), .Y(n3082) );
  AOI22X1 U4048 ( .A(\data_in<8> ), .B(n1099), .C(n3061), .D(n3082), .Y(n3062)
         );
  OAI21X1 U4049 ( .A(n1297), .B(n3063), .C(n3062), .Y(n1848) );
  AOI22X1 U4050 ( .A(\data_in<9> ), .B(n1099), .C(n3064), .D(n3082), .Y(n3065)
         );
  OAI21X1 U4051 ( .A(n1297), .B(n3066), .C(n3065), .Y(n1849) );
  AOI22X1 U4052 ( .A(\data_in<10> ), .B(n1099), .C(n3067), .D(n3082), .Y(n3068) );
  OAI21X1 U4053 ( .A(n1297), .B(n3069), .C(n3068), .Y(n1850) );
  AOI22X1 U4054 ( .A(\data_in<11> ), .B(n1099), .C(n3070), .D(n3082), .Y(n3071) );
  OAI21X1 U4055 ( .A(n1297), .B(n3072), .C(n3071), .Y(n1851) );
  AOI22X1 U4056 ( .A(\data_in<12> ), .B(n1099), .C(n3073), .D(n3082), .Y(n3074) );
  OAI21X1 U4057 ( .A(n1297), .B(n3075), .C(n3074), .Y(n1852) );
  AOI22X1 U4058 ( .A(\data_in<13> ), .B(n1099), .C(n3076), .D(n3082), .Y(n3077) );
  OAI21X1 U4059 ( .A(n1297), .B(n3078), .C(n3077), .Y(n1853) );
  AOI22X1 U4060 ( .A(\data_in<14> ), .B(n1099), .C(n3079), .D(n3082), .Y(n3080) );
  OAI21X1 U4061 ( .A(n1297), .B(n3081), .C(n3080), .Y(n1854) );
  AOI22X1 U4062 ( .A(\data_in<15> ), .B(n1099), .C(n3083), .D(n3082), .Y(n3084) );
  OAI21X1 U4063 ( .A(n1297), .B(n3085), .C(n3084), .Y(n1855) );
  OAI21X1 U4064 ( .A(n794), .B(n3113), .C(n4496), .Y(n3109) );
  AOI22X1 U4065 ( .A(\data_in<8> ), .B(n1100), .C(n3088), .D(n3109), .Y(n3089)
         );
  OAI21X1 U4066 ( .A(n1299), .B(n3090), .C(n3089), .Y(n1856) );
  AOI22X1 U4067 ( .A(\data_in<9> ), .B(n1100), .C(n3091), .D(n3109), .Y(n3092)
         );
  OAI21X1 U4068 ( .A(n1299), .B(n3093), .C(n3092), .Y(n1857) );
  AOI22X1 U4069 ( .A(\data_in<10> ), .B(n1100), .C(n3094), .D(n3109), .Y(n3095) );
  OAI21X1 U4070 ( .A(n1299), .B(n3096), .C(n3095), .Y(n1858) );
  AOI22X1 U4071 ( .A(\data_in<11> ), .B(n1100), .C(n3097), .D(n3109), .Y(n3098) );
  OAI21X1 U4072 ( .A(n1299), .B(n3099), .C(n3098), .Y(n1859) );
  AOI22X1 U4073 ( .A(\data_in<12> ), .B(n1100), .C(n3100), .D(n3109), .Y(n3101) );
  OAI21X1 U4074 ( .A(n1299), .B(n3102), .C(n3101), .Y(n1860) );
  AOI22X1 U4075 ( .A(\data_in<13> ), .B(n1100), .C(n3103), .D(n3109), .Y(n3104) );
  OAI21X1 U4076 ( .A(n1299), .B(n3105), .C(n3104), .Y(n1861) );
  AOI22X1 U4077 ( .A(\data_in<14> ), .B(n1100), .C(n3106), .D(n3109), .Y(n3107) );
  OAI21X1 U4078 ( .A(n1299), .B(n3108), .C(n3107), .Y(n1862) );
  AOI22X1 U4079 ( .A(\data_in<15> ), .B(n1100), .C(n3110), .D(n3109), .Y(n3111) );
  OAI21X1 U4080 ( .A(n1299), .B(n3112), .C(n3111), .Y(n1863) );
  OAI21X1 U4081 ( .A(n3114), .B(n3113), .C(n4496), .Y(n3137) );
  AOI22X1 U4082 ( .A(\data_in<8> ), .B(n1101), .C(n3116), .D(n3137), .Y(n3117)
         );
  OAI21X1 U4083 ( .A(n1301), .B(n3118), .C(n3117), .Y(n1864) );
  AOI22X1 U4084 ( .A(\data_in<9> ), .B(n1101), .C(n3119), .D(n3137), .Y(n3120)
         );
  OAI21X1 U4085 ( .A(n1301), .B(n3121), .C(n3120), .Y(n1865) );
  AOI22X1 U4086 ( .A(\data_in<10> ), .B(n1101), .C(n3122), .D(n3137), .Y(n3123) );
  OAI21X1 U4087 ( .A(n1301), .B(n3124), .C(n3123), .Y(n1866) );
  AOI22X1 U4088 ( .A(\data_in<11> ), .B(n1101), .C(n3125), .D(n3137), .Y(n3126) );
  OAI21X1 U4089 ( .A(n1301), .B(n3127), .C(n3126), .Y(n1867) );
  AOI22X1 U4090 ( .A(\data_in<12> ), .B(n1101), .C(n3128), .D(n3137), .Y(n3129) );
  OAI21X1 U4091 ( .A(n1301), .B(n3130), .C(n3129), .Y(n1868) );
  AOI22X1 U4092 ( .A(\data_in<13> ), .B(n1101), .C(n3131), .D(n3137), .Y(n3132) );
  OAI21X1 U4093 ( .A(n1301), .B(n3133), .C(n3132), .Y(n1869) );
  AOI22X1 U4094 ( .A(\data_in<14> ), .B(n1101), .C(n3134), .D(n3137), .Y(n3135) );
  OAI21X1 U4095 ( .A(n1301), .B(n3136), .C(n3135), .Y(n1870) );
  AOI22X1 U4096 ( .A(\data_in<15> ), .B(n1101), .C(n3138), .D(n3137), .Y(n3139) );
  OAI21X1 U4097 ( .A(n1301), .B(n3140), .C(n3139), .Y(n1871) );
  AOI22X1 U4098 ( .A(\data_in<8> ), .B(n1102), .C(n3142), .D(n1175), .Y(n3143)
         );
  OAI21X1 U4099 ( .A(n1303), .B(n3144), .C(n3143), .Y(n1872) );
  AOI22X1 U4100 ( .A(\data_in<9> ), .B(n1102), .C(n3145), .D(n1175), .Y(n3146)
         );
  OAI21X1 U4101 ( .A(n1303), .B(n3147), .C(n3146), .Y(n1873) );
  AOI22X1 U4102 ( .A(\data_in<10> ), .B(n1102), .C(n3148), .D(n1175), .Y(n3149) );
  OAI21X1 U4103 ( .A(n1303), .B(n3150), .C(n3149), .Y(n1874) );
  AOI22X1 U4104 ( .A(\data_in<11> ), .B(n1102), .C(n3151), .D(n1175), .Y(n3152) );
  OAI21X1 U4105 ( .A(n1303), .B(n3153), .C(n3152), .Y(n1875) );
  AOI22X1 U4106 ( .A(\data_in<12> ), .B(n1102), .C(n3154), .D(n1175), .Y(n3155) );
  OAI21X1 U4107 ( .A(n1303), .B(n3156), .C(n3155), .Y(n1876) );
  AOI22X1 U4108 ( .A(\data_in<13> ), .B(n1102), .C(n3157), .D(n1175), .Y(n3158) );
  OAI21X1 U4109 ( .A(n1303), .B(n3159), .C(n3158), .Y(n1877) );
  AOI22X1 U4110 ( .A(\data_in<14> ), .B(n1102), .C(n3160), .D(n1175), .Y(n3161) );
  OAI21X1 U4111 ( .A(n1303), .B(n3162), .C(n3161), .Y(n1878) );
  AOI22X1 U4112 ( .A(\data_in<15> ), .B(n1102), .C(n3163), .D(n1175), .Y(n3164) );
  OAI21X1 U4113 ( .A(n1303), .B(n3165), .C(n3164), .Y(n1879) );
  OAI21X1 U4114 ( .A(n793), .B(n831), .C(n4496), .Y(n3190) );
  AOI22X1 U4115 ( .A(\data_in<8> ), .B(n1103), .C(n3169), .D(n1527), .Y(n3170)
         );
  OAI21X1 U4116 ( .A(n1305), .B(n3171), .C(n3170), .Y(n1880) );
  AOI22X1 U4117 ( .A(\data_in<9> ), .B(n1103), .C(n3172), .D(n1527), .Y(n3173)
         );
  OAI21X1 U4118 ( .A(n1305), .B(n3174), .C(n3173), .Y(n1881) );
  AOI22X1 U4119 ( .A(\data_in<10> ), .B(n1103), .C(n3175), .D(n1527), .Y(n3176) );
  OAI21X1 U4120 ( .A(n1305), .B(n3177), .C(n3176), .Y(n1882) );
  AOI22X1 U4121 ( .A(\data_in<11> ), .B(n1103), .C(n3178), .D(n1527), .Y(n3179) );
  OAI21X1 U4122 ( .A(n1305), .B(n3180), .C(n3179), .Y(n1883) );
  AOI22X1 U4123 ( .A(\data_in<12> ), .B(n1103), .C(n3181), .D(n1527), .Y(n3182) );
  OAI21X1 U4124 ( .A(n1305), .B(n3183), .C(n3182), .Y(n1884) );
  AOI22X1 U4125 ( .A(\data_in<13> ), .B(n1103), .C(n3184), .D(n1527), .Y(n3185) );
  OAI21X1 U4126 ( .A(n1305), .B(n3186), .C(n3185), .Y(n1885) );
  AOI22X1 U4127 ( .A(\data_in<14> ), .B(n1103), .C(n3187), .D(n1527), .Y(n3188) );
  OAI21X1 U4128 ( .A(n1305), .B(n3189), .C(n3188), .Y(n1886) );
  AOI22X1 U4129 ( .A(\data_in<15> ), .B(n1103), .C(n3191), .D(n1527), .Y(n3192) );
  OAI21X1 U4130 ( .A(n1305), .B(n3193), .C(n3192), .Y(n1887) );
  AOI22X1 U4131 ( .A(\data_in<8> ), .B(n1104), .C(n3194), .D(n1177), .Y(n3195)
         );
  OAI21X1 U4132 ( .A(n1307), .B(n3196), .C(n3195), .Y(n1888) );
  AOI22X1 U4133 ( .A(\data_in<9> ), .B(n1104), .C(n3197), .D(n1177), .Y(n3198)
         );
  OAI21X1 U4134 ( .A(n1307), .B(n3199), .C(n3198), .Y(n1889) );
  AOI22X1 U4135 ( .A(\data_in<10> ), .B(n1104), .C(n3200), .D(n1177), .Y(n3201) );
  OAI21X1 U4136 ( .A(n1307), .B(n3202), .C(n3201), .Y(n1890) );
  AOI22X1 U4137 ( .A(\data_in<11> ), .B(n1104), .C(n3203), .D(n1177), .Y(n3204) );
  OAI21X1 U4138 ( .A(n1307), .B(n3205), .C(n3204), .Y(n1891) );
  AOI22X1 U4139 ( .A(\data_in<12> ), .B(n1104), .C(n3206), .D(n1177), .Y(n3207) );
  OAI21X1 U4140 ( .A(n1307), .B(n3208), .C(n3207), .Y(n1892) );
  AOI22X1 U4141 ( .A(\data_in<13> ), .B(n1104), .C(n3209), .D(n1177), .Y(n3210) );
  OAI21X1 U4142 ( .A(n1307), .B(n3211), .C(n3210), .Y(n1893) );
  AOI22X1 U4143 ( .A(\data_in<14> ), .B(n1104), .C(n3212), .D(n1177), .Y(n3213) );
  OAI21X1 U4144 ( .A(n1307), .B(n3214), .C(n3213), .Y(n1894) );
  AOI22X1 U4145 ( .A(\data_in<15> ), .B(n1104), .C(n3215), .D(n1177), .Y(n3216) );
  OAI21X1 U4146 ( .A(n1307), .B(n3217), .C(n3216), .Y(n1895) );
  AOI22X1 U4147 ( .A(\data_in<8> ), .B(n1105), .C(n3219), .D(n1179), .Y(n3220)
         );
  OAI21X1 U4148 ( .A(n1309), .B(n3221), .C(n3220), .Y(n1896) );
  AOI22X1 U4149 ( .A(\data_in<9> ), .B(n1105), .C(n3222), .D(n1179), .Y(n3223)
         );
  OAI21X1 U4150 ( .A(n1309), .B(n3224), .C(n3223), .Y(n1897) );
  AOI22X1 U4151 ( .A(\data_in<10> ), .B(n1105), .C(n3225), .D(n1179), .Y(n3226) );
  OAI21X1 U4152 ( .A(n1309), .B(n3227), .C(n3226), .Y(n1898) );
  AOI22X1 U4153 ( .A(\data_in<11> ), .B(n1105), .C(n3228), .D(n1179), .Y(n3229) );
  OAI21X1 U4154 ( .A(n1309), .B(n3230), .C(n3229), .Y(n1899) );
  AOI22X1 U4155 ( .A(\data_in<12> ), .B(n1105), .C(n3231), .D(n1179), .Y(n3232) );
  OAI21X1 U4156 ( .A(n1309), .B(n3233), .C(n3232), .Y(n1900) );
  AOI22X1 U4157 ( .A(\data_in<13> ), .B(n1105), .C(n3234), .D(n1179), .Y(n3235) );
  OAI21X1 U4158 ( .A(n1309), .B(n3236), .C(n3235), .Y(n1901) );
  AOI22X1 U4159 ( .A(\data_in<14> ), .B(n1105), .C(n3237), .D(n1179), .Y(n3238) );
  OAI21X1 U4160 ( .A(n1309), .B(n3239), .C(n3238), .Y(n1902) );
  AOI22X1 U4161 ( .A(\data_in<15> ), .B(n1105), .C(n3240), .D(n1179), .Y(n3241) );
  OAI21X1 U4162 ( .A(n1309), .B(n3242), .C(n3241), .Y(n1903) );
  OAI21X1 U4163 ( .A(n1420), .B(n833), .C(n4496), .Y(n3265) );
  AOI22X1 U4164 ( .A(\data_in<8> ), .B(n1106), .C(n3244), .D(n3265), .Y(n3245)
         );
  OAI21X1 U4165 ( .A(n1311), .B(n3246), .C(n3245), .Y(n1904) );
  AOI22X1 U4166 ( .A(\data_in<9> ), .B(n1106), .C(n3247), .D(n3265), .Y(n3248)
         );
  OAI21X1 U4167 ( .A(n1311), .B(n3249), .C(n3248), .Y(n1905) );
  AOI22X1 U4168 ( .A(\data_in<10> ), .B(n1106), .C(n3250), .D(n3265), .Y(n3251) );
  OAI21X1 U4169 ( .A(n1311), .B(n3252), .C(n3251), .Y(n1906) );
  AOI22X1 U4170 ( .A(\data_in<11> ), .B(n1106), .C(n3253), .D(n3265), .Y(n3254) );
  OAI21X1 U4171 ( .A(n1311), .B(n3255), .C(n3254), .Y(n1907) );
  AOI22X1 U4172 ( .A(\data_in<12> ), .B(n1106), .C(n3256), .D(n3265), .Y(n3257) );
  OAI21X1 U4173 ( .A(n1311), .B(n3258), .C(n3257), .Y(n1908) );
  AOI22X1 U4174 ( .A(\data_in<13> ), .B(n1106), .C(n3259), .D(n3265), .Y(n3260) );
  OAI21X1 U4175 ( .A(n1311), .B(n3261), .C(n3260), .Y(n1909) );
  AOI22X1 U4176 ( .A(\data_in<14> ), .B(n1106), .C(n3262), .D(n3265), .Y(n3263) );
  OAI21X1 U4177 ( .A(n1311), .B(n3264), .C(n3263), .Y(n1910) );
  AOI22X1 U4178 ( .A(\data_in<15> ), .B(n1106), .C(n3266), .D(n3265), .Y(n3267) );
  OAI21X1 U4179 ( .A(n1311), .B(n3268), .C(n3267), .Y(n1911) );
  OAI21X1 U4180 ( .A(n3296), .B(n833), .C(n4496), .Y(n3292) );
  AOI22X1 U4181 ( .A(\data_in<8> ), .B(n1107), .C(n3271), .D(n3292), .Y(n3272)
         );
  OAI21X1 U4182 ( .A(n1313), .B(n3273), .C(n3272), .Y(n1912) );
  AOI22X1 U4183 ( .A(\data_in<9> ), .B(n1107), .C(n3274), .D(n3292), .Y(n3275)
         );
  OAI21X1 U4184 ( .A(n1313), .B(n3276), .C(n3275), .Y(n1913) );
  AOI22X1 U4185 ( .A(\data_in<10> ), .B(n1107), .C(n3277), .D(n3292), .Y(n3278) );
  OAI21X1 U4186 ( .A(n1313), .B(n3279), .C(n3278), .Y(n1914) );
  AOI22X1 U4187 ( .A(\data_in<11> ), .B(n1107), .C(n3280), .D(n3292), .Y(n3281) );
  OAI21X1 U4188 ( .A(n1313), .B(n3282), .C(n3281), .Y(n1915) );
  AOI22X1 U4189 ( .A(\data_in<12> ), .B(n1107), .C(n3283), .D(n3292), .Y(n3284) );
  OAI21X1 U4190 ( .A(n1313), .B(n3285), .C(n3284), .Y(n1916) );
  AOI22X1 U4191 ( .A(\data_in<13> ), .B(n1107), .C(n3286), .D(n3292), .Y(n3287) );
  OAI21X1 U4192 ( .A(n1313), .B(n3288), .C(n3287), .Y(n1917) );
  AOI22X1 U4193 ( .A(\data_in<14> ), .B(n1107), .C(n3289), .D(n3292), .Y(n3290) );
  OAI21X1 U4194 ( .A(n1313), .B(n3291), .C(n3290), .Y(n1918) );
  AOI22X1 U4195 ( .A(\data_in<15> ), .B(n1107), .C(n3293), .D(n3292), .Y(n3294) );
  OAI21X1 U4196 ( .A(n1313), .B(n3295), .C(n3294), .Y(n1919) );
  OAI21X1 U4197 ( .A(n3296), .B(n1442), .C(n4496), .Y(n3319) );
  AOI22X1 U4198 ( .A(\data_in<8> ), .B(n1108), .C(n3298), .D(n3319), .Y(n3299)
         );
  OAI21X1 U4199 ( .A(n1315), .B(n3300), .C(n3299), .Y(n1920) );
  AOI22X1 U4200 ( .A(\data_in<9> ), .B(n1108), .C(n3301), .D(n3319), .Y(n3302)
         );
  OAI21X1 U4201 ( .A(n1315), .B(n3303), .C(n3302), .Y(n1921) );
  AOI22X1 U4202 ( .A(\data_in<10> ), .B(n1108), .C(n3304), .D(n3319), .Y(n3305) );
  OAI21X1 U4203 ( .A(n1315), .B(n3306), .C(n3305), .Y(n1922) );
  AOI22X1 U4204 ( .A(\data_in<11> ), .B(n1108), .C(n3307), .D(n3319), .Y(n3308) );
  OAI21X1 U4205 ( .A(n1315), .B(n3309), .C(n3308), .Y(n1923) );
  AOI22X1 U4206 ( .A(\data_in<12> ), .B(n1108), .C(n3310), .D(n3319), .Y(n3311) );
  OAI21X1 U4207 ( .A(n1315), .B(n3312), .C(n3311), .Y(n1924) );
  AOI22X1 U4208 ( .A(\data_in<13> ), .B(n1108), .C(n3313), .D(n3319), .Y(n3314) );
  OAI21X1 U4209 ( .A(n1315), .B(n3315), .C(n3314), .Y(n1925) );
  AOI22X1 U4210 ( .A(\data_in<14> ), .B(n1108), .C(n3316), .D(n3319), .Y(n3317) );
  OAI21X1 U4211 ( .A(n1315), .B(n3318), .C(n3317), .Y(n1926) );
  AOI22X1 U4212 ( .A(\data_in<15> ), .B(n1108), .C(n3320), .D(n3319), .Y(n3321) );
  OAI21X1 U4213 ( .A(n1315), .B(n3322), .C(n3321), .Y(n1927) );
  OAI21X1 U4214 ( .A(n1416), .B(n1442), .C(n1530), .Y(n3347) );
  AOI22X1 U4215 ( .A(\data_in<8> ), .B(n1109), .C(n3326), .D(n3347), .Y(n3327)
         );
  OAI21X1 U4216 ( .A(n1317), .B(n3328), .C(n3327), .Y(n1928) );
  AOI22X1 U4217 ( .A(\data_in<9> ), .B(n1109), .C(n3329), .D(n3347), .Y(n3330)
         );
  OAI21X1 U4218 ( .A(n1317), .B(n3331), .C(n3330), .Y(n1929) );
  AOI22X1 U4219 ( .A(\data_in<10> ), .B(n1109), .C(n3332), .D(n3347), .Y(n3333) );
  OAI21X1 U4220 ( .A(n1317), .B(n3334), .C(n3333), .Y(n1930) );
  AOI22X1 U4221 ( .A(\data_in<11> ), .B(n1109), .C(n3335), .D(n3347), .Y(n3336) );
  OAI21X1 U4222 ( .A(n1317), .B(n3337), .C(n3336), .Y(n1931) );
  AOI22X1 U4223 ( .A(\data_in<12> ), .B(n1109), .C(n3338), .D(n3347), .Y(n3339) );
  OAI21X1 U4224 ( .A(n1317), .B(n3340), .C(n3339), .Y(n1932) );
  AOI22X1 U4225 ( .A(\data_in<13> ), .B(n1109), .C(n3341), .D(n3347), .Y(n3342) );
  OAI21X1 U4226 ( .A(n1317), .B(n3343), .C(n3342), .Y(n1933) );
  AOI22X1 U4227 ( .A(\data_in<14> ), .B(n1109), .C(n3344), .D(n3347), .Y(n3345) );
  OAI21X1 U4228 ( .A(n1317), .B(n3346), .C(n3345), .Y(n1934) );
  AOI22X1 U4229 ( .A(\data_in<15> ), .B(n1109), .C(n3348), .D(n3347), .Y(n3349) );
  OAI21X1 U4230 ( .A(n1317), .B(n3350), .C(n3349), .Y(n1935) );
  AOI22X1 U4231 ( .A(\data_in<8> ), .B(n1110), .C(n3351), .D(n1181), .Y(n3352)
         );
  OAI21X1 U4232 ( .A(n1319), .B(n3353), .C(n3352), .Y(n1936) );
  AOI22X1 U4233 ( .A(\data_in<9> ), .B(n1110), .C(n3354), .D(n1181), .Y(n3355)
         );
  OAI21X1 U4234 ( .A(n1319), .B(n3356), .C(n3355), .Y(n1937) );
  AOI22X1 U4235 ( .A(\data_in<10> ), .B(n1110), .C(n3357), .D(n1181), .Y(n3358) );
  OAI21X1 U4236 ( .A(n1319), .B(n3359), .C(n3358), .Y(n1938) );
  AOI22X1 U4237 ( .A(\data_in<11> ), .B(n1110), .C(n3360), .D(n1181), .Y(n3361) );
  OAI21X1 U4238 ( .A(n1319), .B(n3362), .C(n3361), .Y(n1939) );
  AOI22X1 U4239 ( .A(\data_in<12> ), .B(n1110), .C(n3363), .D(n1181), .Y(n3364) );
  OAI21X1 U4240 ( .A(n1319), .B(n3365), .C(n3364), .Y(n1940) );
  AOI22X1 U4241 ( .A(\data_in<13> ), .B(n1110), .C(n3366), .D(n1181), .Y(n3367) );
  OAI21X1 U4242 ( .A(n1319), .B(n3368), .C(n3367), .Y(n1941) );
  AOI22X1 U4243 ( .A(\data_in<14> ), .B(n1110), .C(n3369), .D(n1181), .Y(n3370) );
  OAI21X1 U4244 ( .A(n1319), .B(n3371), .C(n3370), .Y(n1942) );
  AOI22X1 U4245 ( .A(\data_in<15> ), .B(n1110), .C(n3372), .D(n1181), .Y(n3373) );
  OAI21X1 U4246 ( .A(n1319), .B(n3374), .C(n3373), .Y(n1943) );
  AOI22X1 U4247 ( .A(\data_in<8> ), .B(n1111), .C(n3376), .D(n1183), .Y(n3377)
         );
  OAI21X1 U4248 ( .A(n1321), .B(n3378), .C(n3377), .Y(n1944) );
  AOI22X1 U4249 ( .A(\data_in<9> ), .B(n1111), .C(n3379), .D(n1183), .Y(n3380)
         );
  OAI21X1 U4250 ( .A(n1321), .B(n3381), .C(n3380), .Y(n1945) );
  AOI22X1 U4251 ( .A(\data_in<10> ), .B(n1111), .C(n3382), .D(n1183), .Y(n3383) );
  OAI21X1 U4252 ( .A(n1321), .B(n3384), .C(n3383), .Y(n1946) );
  AOI22X1 U4253 ( .A(\data_in<11> ), .B(n1111), .C(n3385), .D(n1183), .Y(n3386) );
  OAI21X1 U4254 ( .A(n1321), .B(n3387), .C(n3386), .Y(n1947) );
  AOI22X1 U4255 ( .A(\data_in<12> ), .B(n1111), .C(n3388), .D(n1183), .Y(n3389) );
  OAI21X1 U4256 ( .A(n1321), .B(n3390), .C(n3389), .Y(n1948) );
  AOI22X1 U4257 ( .A(\data_in<13> ), .B(n1111), .C(n3391), .D(n1183), .Y(n3392) );
  OAI21X1 U4258 ( .A(n1321), .B(n3393), .C(n3392), .Y(n1949) );
  AOI22X1 U4259 ( .A(\data_in<14> ), .B(n1111), .C(n3394), .D(n1183), .Y(n3395) );
  OAI21X1 U4260 ( .A(n1321), .B(n3396), .C(n3395), .Y(n1950) );
  AOI22X1 U4261 ( .A(\data_in<15> ), .B(n1111), .C(n3397), .D(n1183), .Y(n3398) );
  OAI21X1 U4262 ( .A(n1321), .B(n3399), .C(n3398), .Y(n1951) );
  AOI22X1 U4263 ( .A(\data_in<8> ), .B(n1112), .C(n3400), .D(n1185), .Y(n3401)
         );
  OAI21X1 U4264 ( .A(n1323), .B(n3402), .C(n3401), .Y(n1952) );
  AOI22X1 U4265 ( .A(\data_in<9> ), .B(n1112), .C(n3403), .D(n1185), .Y(n3404)
         );
  OAI21X1 U4266 ( .A(n1323), .B(n3405), .C(n3404), .Y(n1953) );
  AOI22X1 U4267 ( .A(\data_in<10> ), .B(n1112), .C(n3406), .D(n1185), .Y(n3407) );
  OAI21X1 U4268 ( .A(n1323), .B(n3408), .C(n3407), .Y(n1954) );
  AOI22X1 U4269 ( .A(\data_in<11> ), .B(n1112), .C(n3409), .D(n1185), .Y(n3410) );
  OAI21X1 U4270 ( .A(n1323), .B(n3411), .C(n3410), .Y(n1955) );
  AOI22X1 U4271 ( .A(\data_in<12> ), .B(n1112), .C(n3412), .D(n1185), .Y(n3413) );
  OAI21X1 U4272 ( .A(n1323), .B(n3414), .C(n3413), .Y(n1956) );
  AOI22X1 U4273 ( .A(\data_in<13> ), .B(n1112), .C(n3415), .D(n1185), .Y(n3416) );
  OAI21X1 U4274 ( .A(n1323), .B(n3417), .C(n3416), .Y(n1957) );
  AOI22X1 U4275 ( .A(\data_in<14> ), .B(n1112), .C(n3418), .D(n1185), .Y(n3419) );
  OAI21X1 U4276 ( .A(n1323), .B(n3420), .C(n3419), .Y(n1958) );
  AOI22X1 U4277 ( .A(\data_in<15> ), .B(n1112), .C(n3421), .D(n1185), .Y(n3422) );
  OAI21X1 U4278 ( .A(n1323), .B(n3423), .C(n3422), .Y(n1959) );
  AOI22X1 U4279 ( .A(\data_in<8> ), .B(n1113), .C(n3424), .D(n1187), .Y(n3425)
         );
  OAI21X1 U4280 ( .A(n1325), .B(n3426), .C(n3425), .Y(n1960) );
  AOI22X1 U4281 ( .A(\data_in<9> ), .B(n1113), .C(n3427), .D(n1187), .Y(n3428)
         );
  OAI21X1 U4282 ( .A(n1325), .B(n3429), .C(n3428), .Y(n1961) );
  AOI22X1 U4283 ( .A(\data_in<10> ), .B(n1113), .C(n3430), .D(n1187), .Y(n3431) );
  OAI21X1 U4284 ( .A(n1325), .B(n3432), .C(n3431), .Y(n1962) );
  AOI22X1 U4285 ( .A(\data_in<11> ), .B(n1113), .C(n3433), .D(n1187), .Y(n3434) );
  OAI21X1 U4286 ( .A(n1325), .B(n3435), .C(n3434), .Y(n1963) );
  AOI22X1 U4287 ( .A(\data_in<12> ), .B(n1113), .C(n3436), .D(n1187), .Y(n3437) );
  OAI21X1 U4288 ( .A(n1325), .B(n3438), .C(n3437), .Y(n1964) );
  AOI22X1 U4289 ( .A(\data_in<13> ), .B(n1113), .C(n3439), .D(n1187), .Y(n3440) );
  OAI21X1 U4290 ( .A(n1325), .B(n3441), .C(n3440), .Y(n1965) );
  AOI22X1 U4291 ( .A(\data_in<14> ), .B(n1113), .C(n3442), .D(n1187), .Y(n3443) );
  OAI21X1 U4292 ( .A(n1325), .B(n3444), .C(n3443), .Y(n1966) );
  AOI22X1 U4293 ( .A(\data_in<15> ), .B(n1113), .C(n3445), .D(n1187), .Y(n3446) );
  OAI21X1 U4294 ( .A(n1325), .B(n3447), .C(n3446), .Y(n1967) );
  AOI22X1 U4295 ( .A(\data_in<8> ), .B(n1114), .C(n3448), .D(n1189), .Y(n3449)
         );
  OAI21X1 U4296 ( .A(n1327), .B(n3450), .C(n3449), .Y(n1968) );
  AOI22X1 U4297 ( .A(\data_in<9> ), .B(n1114), .C(n3451), .D(n1189), .Y(n3452)
         );
  OAI21X1 U4298 ( .A(n1327), .B(n3453), .C(n3452), .Y(n1969) );
  AOI22X1 U4299 ( .A(\data_in<10> ), .B(n1114), .C(n3454), .D(n1189), .Y(n3455) );
  OAI21X1 U4300 ( .A(n1327), .B(n3456), .C(n3455), .Y(n1970) );
  AOI22X1 U4301 ( .A(\data_in<11> ), .B(n1114), .C(n3457), .D(n1189), .Y(n3458) );
  OAI21X1 U4302 ( .A(n1327), .B(n3459), .C(n3458), .Y(n1971) );
  AOI22X1 U4303 ( .A(\data_in<12> ), .B(n1114), .C(n3460), .D(n1189), .Y(n3461) );
  OAI21X1 U4304 ( .A(n1327), .B(n3462), .C(n3461), .Y(n1972) );
  AOI22X1 U4305 ( .A(\data_in<13> ), .B(n1114), .C(n3463), .D(n1189), .Y(n3464) );
  OAI21X1 U4306 ( .A(n1327), .B(n3465), .C(n3464), .Y(n1973) );
  AOI22X1 U4307 ( .A(\data_in<14> ), .B(n1114), .C(n3466), .D(n1189), .Y(n3467) );
  OAI21X1 U4308 ( .A(n1327), .B(n3468), .C(n3467), .Y(n1974) );
  AOI22X1 U4309 ( .A(\data_in<15> ), .B(n1114), .C(n3469), .D(n1189), .Y(n3470) );
  OAI21X1 U4310 ( .A(n1327), .B(n3471), .C(n3470), .Y(n1975) );
  AOI22X1 U4311 ( .A(\data_in<8> ), .B(n1115), .C(n3473), .D(n1191), .Y(n3474)
         );
  OAI21X1 U4312 ( .A(n1329), .B(n3475), .C(n3474), .Y(n1976) );
  AOI22X1 U4313 ( .A(\data_in<9> ), .B(n1115), .C(n3476), .D(n1191), .Y(n3477)
         );
  OAI21X1 U4314 ( .A(n1329), .B(n3478), .C(n3477), .Y(n1977) );
  AOI22X1 U4315 ( .A(\data_in<10> ), .B(n1115), .C(n3479), .D(n1191), .Y(n3480) );
  OAI21X1 U4316 ( .A(n1329), .B(n3481), .C(n3480), .Y(n1978) );
  AOI22X1 U4317 ( .A(\data_in<11> ), .B(n1115), .C(n3482), .D(n1191), .Y(n3483) );
  OAI21X1 U4318 ( .A(n1329), .B(n3484), .C(n3483), .Y(n1979) );
  AOI22X1 U4319 ( .A(\data_in<12> ), .B(n1115), .C(n3485), .D(n1191), .Y(n3486) );
  OAI21X1 U4320 ( .A(n1329), .B(n3487), .C(n3486), .Y(n1980) );
  AOI22X1 U4321 ( .A(\data_in<13> ), .B(n1115), .C(n3488), .D(n1191), .Y(n3489) );
  OAI21X1 U4322 ( .A(n1329), .B(n3490), .C(n3489), .Y(n1981) );
  AOI22X1 U4323 ( .A(\data_in<14> ), .B(n1115), .C(n3491), .D(n1191), .Y(n3492) );
  OAI21X1 U4324 ( .A(n1329), .B(n3493), .C(n3492), .Y(n1982) );
  AOI22X1 U4325 ( .A(\data_in<15> ), .B(n1115), .C(n3494), .D(n1191), .Y(n3495) );
  OAI21X1 U4326 ( .A(n1329), .B(n3496), .C(n3495), .Y(n1983) );
  AOI22X1 U4327 ( .A(\data_in<8> ), .B(n1116), .C(n3498), .D(n1193), .Y(n3499)
         );
  OAI21X1 U4328 ( .A(n1331), .B(n3500), .C(n3499), .Y(n1984) );
  AOI22X1 U4329 ( .A(\data_in<9> ), .B(n1116), .C(n3501), .D(n1193), .Y(n3502)
         );
  OAI21X1 U4330 ( .A(n1331), .B(n3503), .C(n3502), .Y(n1985) );
  AOI22X1 U4331 ( .A(\data_in<10> ), .B(n1116), .C(n3504), .D(n1193), .Y(n3505) );
  OAI21X1 U4332 ( .A(n1331), .B(n3506), .C(n3505), .Y(n1986) );
  AOI22X1 U4333 ( .A(\data_in<11> ), .B(n1116), .C(n3507), .D(n1193), .Y(n3508) );
  OAI21X1 U4334 ( .A(n1331), .B(n3509), .C(n3508), .Y(n1987) );
  AOI22X1 U4335 ( .A(\data_in<12> ), .B(n1116), .C(n3510), .D(n1193), .Y(n3511) );
  OAI21X1 U4336 ( .A(n1331), .B(n3512), .C(n3511), .Y(n1988) );
  AOI22X1 U4337 ( .A(\data_in<13> ), .B(n1116), .C(n3513), .D(n1193), .Y(n3514) );
  OAI21X1 U4338 ( .A(n1331), .B(n3515), .C(n3514), .Y(n1989) );
  AOI22X1 U4339 ( .A(\data_in<14> ), .B(n1116), .C(n3516), .D(n1193), .Y(n3517) );
  OAI21X1 U4340 ( .A(n1331), .B(n3518), .C(n3517), .Y(n1990) );
  AOI22X1 U4341 ( .A(\data_in<15> ), .B(n1116), .C(n3519), .D(n1193), .Y(n3520) );
  OAI21X1 U4342 ( .A(n1331), .B(n3521), .C(n3520), .Y(n1991) );
  AOI22X1 U4343 ( .A(\data_in<8> ), .B(n1117), .C(n3522), .D(n1195), .Y(n3523)
         );
  OAI21X1 U4344 ( .A(n1333), .B(n3524), .C(n3523), .Y(n1992) );
  AOI22X1 U4345 ( .A(\data_in<9> ), .B(n1117), .C(n3525), .D(n1195), .Y(n3526)
         );
  OAI21X1 U4346 ( .A(n1333), .B(n3527), .C(n3526), .Y(n1993) );
  AOI22X1 U4347 ( .A(\data_in<10> ), .B(n1117), .C(n3528), .D(n1195), .Y(n3529) );
  OAI21X1 U4348 ( .A(n1333), .B(n3530), .C(n3529), .Y(n1994) );
  AOI22X1 U4349 ( .A(\data_in<11> ), .B(n1117), .C(n3531), .D(n1195), .Y(n3532) );
  OAI21X1 U4350 ( .A(n1333), .B(n3533), .C(n3532), .Y(n1995) );
  AOI22X1 U4351 ( .A(\data_in<12> ), .B(n1117), .C(n3534), .D(n1195), .Y(n3535) );
  OAI21X1 U4352 ( .A(n1333), .B(n3536), .C(n3535), .Y(n1996) );
  AOI22X1 U4353 ( .A(\data_in<13> ), .B(n1117), .C(n3537), .D(n1195), .Y(n3538) );
  OAI21X1 U4354 ( .A(n1333), .B(n3539), .C(n3538), .Y(n1997) );
  AOI22X1 U4355 ( .A(\data_in<14> ), .B(n1117), .C(n3540), .D(n1195), .Y(n3541) );
  OAI21X1 U4356 ( .A(n1333), .B(n3542), .C(n3541), .Y(n1998) );
  AOI22X1 U4357 ( .A(\data_in<15> ), .B(n1117), .C(n3543), .D(n1195), .Y(n3544) );
  OAI21X1 U4358 ( .A(n1333), .B(n3545), .C(n3544), .Y(n1999) );
  AOI22X1 U4359 ( .A(\data_in<8> ), .B(n1118), .C(n3547), .D(n1197), .Y(n3548)
         );
  OAI21X1 U4360 ( .A(n1335), .B(n3549), .C(n3548), .Y(n2000) );
  AOI22X1 U4361 ( .A(\data_in<9> ), .B(n1118), .C(n3550), .D(n1197), .Y(n3551)
         );
  OAI21X1 U4362 ( .A(n1335), .B(n3552), .C(n3551), .Y(n2001) );
  AOI22X1 U4363 ( .A(\data_in<10> ), .B(n1118), .C(n3553), .D(n1197), .Y(n3554) );
  OAI21X1 U4364 ( .A(n1335), .B(n3555), .C(n3554), .Y(n2002) );
  AOI22X1 U4365 ( .A(\data_in<11> ), .B(n1118), .C(n3556), .D(n1197), .Y(n3557) );
  OAI21X1 U4366 ( .A(n1335), .B(n3558), .C(n3557), .Y(n2003) );
  AOI22X1 U4367 ( .A(\data_in<12> ), .B(n1118), .C(n3559), .D(n1197), .Y(n3560) );
  OAI21X1 U4368 ( .A(n1335), .B(n3561), .C(n3560), .Y(n2004) );
  AOI22X1 U4369 ( .A(\data_in<13> ), .B(n1118), .C(n3562), .D(n1197), .Y(n3563) );
  OAI21X1 U4370 ( .A(n1335), .B(n3564), .C(n3563), .Y(n2005) );
  AOI22X1 U4371 ( .A(\data_in<14> ), .B(n1118), .C(n3565), .D(n1197), .Y(n3566) );
  OAI21X1 U4372 ( .A(n1335), .B(n3567), .C(n3566), .Y(n2006) );
  AOI22X1 U4373 ( .A(\data_in<15> ), .B(n1118), .C(n3568), .D(n1197), .Y(n3569) );
  OAI21X1 U4374 ( .A(n1335), .B(n3570), .C(n3569), .Y(n2007) );
  AOI22X1 U4375 ( .A(\data_in<8> ), .B(n1119), .C(n3572), .D(n1199), .Y(n3573)
         );
  OAI21X1 U4376 ( .A(n1337), .B(n3574), .C(n3573), .Y(n2008) );
  AOI22X1 U4377 ( .A(\data_in<9> ), .B(n1119), .C(n3575), .D(n1199), .Y(n3576)
         );
  OAI21X1 U4378 ( .A(n1337), .B(n3577), .C(n3576), .Y(n2009) );
  AOI22X1 U4379 ( .A(\data_in<10> ), .B(n1119), .C(n3578), .D(n1199), .Y(n3579) );
  OAI21X1 U4380 ( .A(n1337), .B(n3580), .C(n3579), .Y(n2010) );
  AOI22X1 U4381 ( .A(\data_in<11> ), .B(n1119), .C(n3581), .D(n1199), .Y(n3582) );
  OAI21X1 U4382 ( .A(n1337), .B(n3583), .C(n3582), .Y(n2011) );
  AOI22X1 U4383 ( .A(\data_in<12> ), .B(n1119), .C(n3584), .D(n1199), .Y(n3585) );
  OAI21X1 U4384 ( .A(n1337), .B(n3586), .C(n3585), .Y(n2012) );
  AOI22X1 U4385 ( .A(\data_in<13> ), .B(n1119), .C(n3587), .D(n1199), .Y(n3588) );
  OAI21X1 U4386 ( .A(n1337), .B(n3589), .C(n3588), .Y(n2013) );
  AOI22X1 U4387 ( .A(\data_in<14> ), .B(n1119), .C(n3590), .D(n1199), .Y(n3591) );
  OAI21X1 U4388 ( .A(n1337), .B(n3592), .C(n3591), .Y(n2014) );
  AOI22X1 U4389 ( .A(\data_in<15> ), .B(n1119), .C(n3593), .D(n1199), .Y(n3594) );
  OAI21X1 U4390 ( .A(n1337), .B(n3595), .C(n3594), .Y(n2015) );
  AOI22X1 U4391 ( .A(\data_in<8> ), .B(n1120), .C(n3596), .D(n1201), .Y(n3597)
         );
  OAI21X1 U4392 ( .A(n1339), .B(n3598), .C(n3597), .Y(n2016) );
  AOI22X1 U4393 ( .A(\data_in<9> ), .B(n1120), .C(n3599), .D(n1201), .Y(n3600)
         );
  OAI21X1 U4394 ( .A(n1339), .B(n3601), .C(n3600), .Y(n2017) );
  AOI22X1 U4395 ( .A(\data_in<10> ), .B(n1120), .C(n3602), .D(n1201), .Y(n3603) );
  OAI21X1 U4396 ( .A(n1339), .B(n3604), .C(n3603), .Y(n2018) );
  AOI22X1 U4397 ( .A(\data_in<11> ), .B(n1120), .C(n3605), .D(n1201), .Y(n3606) );
  OAI21X1 U4398 ( .A(n1339), .B(n3607), .C(n3606), .Y(n2019) );
  AOI22X1 U4399 ( .A(\data_in<12> ), .B(n1120), .C(n3608), .D(n1201), .Y(n3609) );
  OAI21X1 U4400 ( .A(n1339), .B(n3610), .C(n3609), .Y(n2020) );
  AOI22X1 U4401 ( .A(\data_in<13> ), .B(n1120), .C(n3611), .D(n1201), .Y(n3612) );
  OAI21X1 U4402 ( .A(n1339), .B(n3613), .C(n3612), .Y(n2021) );
  AOI22X1 U4403 ( .A(\data_in<14> ), .B(n1120), .C(n3614), .D(n1201), .Y(n3615) );
  OAI21X1 U4404 ( .A(n1339), .B(n3616), .C(n3615), .Y(n2022) );
  AOI22X1 U4405 ( .A(\data_in<15> ), .B(n1120), .C(n3617), .D(n1201), .Y(n3618) );
  OAI21X1 U4406 ( .A(n1339), .B(n3619), .C(n3618), .Y(n2023) );
  AOI22X1 U4407 ( .A(\data_in<8> ), .B(n1121), .C(n3621), .D(n1203), .Y(n3622)
         );
  OAI21X1 U4408 ( .A(n1341), .B(n3623), .C(n3622), .Y(n2024) );
  AOI22X1 U4409 ( .A(\data_in<9> ), .B(n1121), .C(n3624), .D(n1203), .Y(n3625)
         );
  OAI21X1 U4410 ( .A(n1341), .B(n3626), .C(n3625), .Y(n2025) );
  AOI22X1 U4411 ( .A(\data_in<10> ), .B(n1121), .C(n3627), .D(n1203), .Y(n3628) );
  OAI21X1 U4412 ( .A(n1341), .B(n3629), .C(n3628), .Y(n2026) );
  AOI22X1 U4413 ( .A(\data_in<11> ), .B(n1121), .C(n3630), .D(n1203), .Y(n3631) );
  OAI21X1 U4414 ( .A(n1341), .B(n3632), .C(n3631), .Y(n2027) );
  AOI22X1 U4415 ( .A(\data_in<12> ), .B(n1121), .C(n3633), .D(n1203), .Y(n3634) );
  OAI21X1 U4416 ( .A(n1341), .B(n3635), .C(n3634), .Y(n2028) );
  AOI22X1 U4417 ( .A(\data_in<13> ), .B(n1121), .C(n3636), .D(n1203), .Y(n3637) );
  OAI21X1 U4418 ( .A(n1341), .B(n3638), .C(n3637), .Y(n2029) );
  AOI22X1 U4419 ( .A(\data_in<14> ), .B(n1121), .C(n3639), .D(n1203), .Y(n3640) );
  OAI21X1 U4420 ( .A(n1341), .B(n3641), .C(n3640), .Y(n2030) );
  AOI22X1 U4421 ( .A(\data_in<15> ), .B(n1121), .C(n3642), .D(n1203), .Y(n3643) );
  OAI21X1 U4422 ( .A(n1341), .B(n3644), .C(n3643), .Y(n2031) );
  AOI22X1 U4423 ( .A(\data_in<8> ), .B(n1122), .C(n3645), .D(n1205), .Y(n3646)
         );
  OAI21X1 U4424 ( .A(n1343), .B(n3647), .C(n3646), .Y(n2032) );
  AOI22X1 U4425 ( .A(\data_in<9> ), .B(n1122), .C(n3648), .D(n1205), .Y(n3649)
         );
  OAI21X1 U4426 ( .A(n1343), .B(n3650), .C(n3649), .Y(n2033) );
  AOI22X1 U4427 ( .A(\data_in<10> ), .B(n1122), .C(n3651), .D(n1205), .Y(n3652) );
  OAI21X1 U4428 ( .A(n1343), .B(n3653), .C(n3652), .Y(n2034) );
  AOI22X1 U4429 ( .A(\data_in<11> ), .B(n1122), .C(n3654), .D(n1205), .Y(n3655) );
  OAI21X1 U4430 ( .A(n1343), .B(n3656), .C(n3655), .Y(n2035) );
  AOI22X1 U4431 ( .A(\data_in<12> ), .B(n1122), .C(n3657), .D(n1205), .Y(n3658) );
  OAI21X1 U4432 ( .A(n1343), .B(n3659), .C(n3658), .Y(n2036) );
  AOI22X1 U4433 ( .A(\data_in<13> ), .B(n1122), .C(n3660), .D(n1205), .Y(n3661) );
  OAI21X1 U4434 ( .A(n1343), .B(n3662), .C(n3661), .Y(n2037) );
  AOI22X1 U4435 ( .A(\data_in<14> ), .B(n1122), .C(n3663), .D(n1205), .Y(n3664) );
  OAI21X1 U4436 ( .A(n1343), .B(n3665), .C(n3664), .Y(n2038) );
  AOI22X1 U4437 ( .A(\data_in<15> ), .B(n1122), .C(n3666), .D(n1205), .Y(n3667) );
  OAI21X1 U4438 ( .A(n1343), .B(n3668), .C(n3667), .Y(n2039) );
  AOI22X1 U4439 ( .A(\data_in<8> ), .B(n1123), .C(n3670), .D(n1207), .Y(n3671)
         );
  OAI21X1 U4440 ( .A(n1345), .B(n3672), .C(n3671), .Y(n2040) );
  AOI22X1 U4441 ( .A(\data_in<9> ), .B(n1123), .C(n3673), .D(n1207), .Y(n3674)
         );
  OAI21X1 U4442 ( .A(n1345), .B(n3675), .C(n3674), .Y(n2041) );
  AOI22X1 U4443 ( .A(\data_in<10> ), .B(n1123), .C(n3676), .D(n1207), .Y(n3677) );
  OAI21X1 U4444 ( .A(n1345), .B(n3678), .C(n3677), .Y(n2042) );
  AOI22X1 U4445 ( .A(\data_in<11> ), .B(n1123), .C(n3679), .D(n1207), .Y(n3680) );
  OAI21X1 U4446 ( .A(n1345), .B(n3681), .C(n3680), .Y(n2043) );
  AOI22X1 U4447 ( .A(\data_in<12> ), .B(n1123), .C(n3682), .D(n1207), .Y(n3683) );
  OAI21X1 U4448 ( .A(n1345), .B(n3684), .C(n3683), .Y(n2044) );
  AOI22X1 U4449 ( .A(\data_in<13> ), .B(n1123), .C(n3685), .D(n1207), .Y(n3686) );
  OAI21X1 U4450 ( .A(n1345), .B(n3687), .C(n3686), .Y(n2045) );
  AOI22X1 U4451 ( .A(\data_in<14> ), .B(n1123), .C(n3688), .D(n1207), .Y(n3689) );
  OAI21X1 U4452 ( .A(n1345), .B(n3690), .C(n3689), .Y(n2046) );
  AOI22X1 U4453 ( .A(\data_in<15> ), .B(n1123), .C(n3691), .D(n1207), .Y(n3692) );
  OAI21X1 U4454 ( .A(n1345), .B(n3693), .C(n3692), .Y(n2047) );
  AOI22X1 U4455 ( .A(\data_in<8> ), .B(n1124), .C(n3694), .D(n1209), .Y(n3695)
         );
  OAI21X1 U4456 ( .A(n1347), .B(n3696), .C(n3695), .Y(n2048) );
  AOI22X1 U4457 ( .A(\data_in<9> ), .B(n1124), .C(n3697), .D(n1209), .Y(n3698)
         );
  OAI21X1 U4458 ( .A(n1347), .B(n3699), .C(n3698), .Y(n2049) );
  AOI22X1 U4459 ( .A(\data_in<10> ), .B(n1124), .C(n3700), .D(n1209), .Y(n3701) );
  OAI21X1 U4460 ( .A(n1347), .B(n3702), .C(n3701), .Y(n2050) );
  AOI22X1 U4461 ( .A(\data_in<11> ), .B(n1124), .C(n3703), .D(n1209), .Y(n3704) );
  OAI21X1 U4462 ( .A(n1347), .B(n3705), .C(n3704), .Y(n2051) );
  AOI22X1 U4463 ( .A(\data_in<12> ), .B(n1124), .C(n3706), .D(n1209), .Y(n3707) );
  OAI21X1 U4464 ( .A(n1347), .B(n3708), .C(n3707), .Y(n2052) );
  AOI22X1 U4465 ( .A(\data_in<13> ), .B(n1124), .C(n3709), .D(n1209), .Y(n3710) );
  OAI21X1 U4466 ( .A(n1347), .B(n3711), .C(n3710), .Y(n2053) );
  AOI22X1 U4467 ( .A(\data_in<14> ), .B(n1124), .C(n3712), .D(n1209), .Y(n3713) );
  OAI21X1 U4468 ( .A(n1347), .B(n3714), .C(n3713), .Y(n2054) );
  AOI22X1 U4469 ( .A(\data_in<15> ), .B(n1124), .C(n3715), .D(n1209), .Y(n3716) );
  OAI21X1 U4470 ( .A(n1347), .B(n3717), .C(n3716), .Y(n2055) );
  AOI22X1 U4471 ( .A(\data_in<8> ), .B(n1125), .C(n3719), .D(n1211), .Y(n3720)
         );
  OAI21X1 U4472 ( .A(n1349), .B(n3721), .C(n3720), .Y(n2056) );
  AOI22X1 U4473 ( .A(\data_in<9> ), .B(n1125), .C(n3722), .D(n1211), .Y(n3723)
         );
  OAI21X1 U4474 ( .A(n1349), .B(n3724), .C(n3723), .Y(n2057) );
  AOI22X1 U4475 ( .A(\data_in<10> ), .B(n1125), .C(n3725), .D(n1211), .Y(n3726) );
  OAI21X1 U4476 ( .A(n1349), .B(n3727), .C(n3726), .Y(n2058) );
  AOI22X1 U4477 ( .A(\data_in<11> ), .B(n1125), .C(n3728), .D(n1211), .Y(n3729) );
  OAI21X1 U4478 ( .A(n1349), .B(n3730), .C(n3729), .Y(n2059) );
  AOI22X1 U4479 ( .A(\data_in<12> ), .B(n1125), .C(n3731), .D(n1211), .Y(n3732) );
  OAI21X1 U4480 ( .A(n1349), .B(n3733), .C(n3732), .Y(n2060) );
  AOI22X1 U4481 ( .A(\data_in<13> ), .B(n1125), .C(n3734), .D(n1211), .Y(n3735) );
  OAI21X1 U4482 ( .A(n1349), .B(n3736), .C(n3735), .Y(n2061) );
  AOI22X1 U4483 ( .A(\data_in<14> ), .B(n1125), .C(n3737), .D(n1211), .Y(n3738) );
  OAI21X1 U4484 ( .A(n1349), .B(n3739), .C(n3738), .Y(n2062) );
  AOI22X1 U4485 ( .A(\data_in<15> ), .B(n1125), .C(n3740), .D(n1211), .Y(n3741) );
  OAI21X1 U4486 ( .A(n1349), .B(n3742), .C(n3741), .Y(n2063) );
  AOI22X1 U4487 ( .A(\data_in<8> ), .B(n1126), .C(n3743), .D(n1213), .Y(n3744)
         );
  OAI21X1 U4488 ( .A(n1351), .B(n3745), .C(n3744), .Y(n2064) );
  AOI22X1 U4489 ( .A(\data_in<9> ), .B(n1126), .C(n3746), .D(n1213), .Y(n3747)
         );
  OAI21X1 U4490 ( .A(n1351), .B(n3748), .C(n3747), .Y(n2065) );
  AOI22X1 U4491 ( .A(\data_in<10> ), .B(n1126), .C(n3749), .D(n1213), .Y(n3750) );
  OAI21X1 U4492 ( .A(n1351), .B(n3751), .C(n3750), .Y(n2066) );
  AOI22X1 U4493 ( .A(\data_in<11> ), .B(n1126), .C(n3752), .D(n1213), .Y(n3753) );
  OAI21X1 U4494 ( .A(n1351), .B(n3754), .C(n3753), .Y(n2067) );
  AOI22X1 U4495 ( .A(\data_in<12> ), .B(n1126), .C(n3755), .D(n1213), .Y(n3756) );
  OAI21X1 U4496 ( .A(n1351), .B(n3757), .C(n3756), .Y(n2068) );
  AOI22X1 U4497 ( .A(\data_in<13> ), .B(n1126), .C(n3758), .D(n1213), .Y(n3759) );
  OAI21X1 U4498 ( .A(n1351), .B(n3760), .C(n3759), .Y(n2069) );
  AOI22X1 U4499 ( .A(\data_in<14> ), .B(n1126), .C(n3761), .D(n1213), .Y(n3762) );
  OAI21X1 U4500 ( .A(n1351), .B(n3763), .C(n3762), .Y(n2070) );
  AOI22X1 U4501 ( .A(\data_in<15> ), .B(n1126), .C(n3764), .D(n1213), .Y(n3765) );
  OAI21X1 U4502 ( .A(n1351), .B(n3766), .C(n3765), .Y(n2071) );
  OAI21X1 U4503 ( .A(n3793), .B(n788), .C(n1530), .Y(n3789) );
  AOI22X1 U4504 ( .A(\data_in<8> ), .B(n1127), .C(n3768), .D(n3789), .Y(n3769)
         );
  OAI21X1 U4505 ( .A(n1353), .B(n3770), .C(n3769), .Y(n2072) );
  AOI22X1 U4506 ( .A(\data_in<9> ), .B(n1127), .C(n3771), .D(n3789), .Y(n3772)
         );
  OAI21X1 U4507 ( .A(n1353), .B(n3773), .C(n3772), .Y(n2073) );
  AOI22X1 U4508 ( .A(\data_in<10> ), .B(n1127), .C(n3774), .D(n3789), .Y(n3775) );
  OAI21X1 U4509 ( .A(n1353), .B(n3776), .C(n3775), .Y(n2074) );
  AOI22X1 U4510 ( .A(\data_in<11> ), .B(n1127), .C(n3777), .D(n3789), .Y(n3778) );
  OAI21X1 U4511 ( .A(n1353), .B(n3779), .C(n3778), .Y(n2075) );
  AOI22X1 U4512 ( .A(\data_in<12> ), .B(n1127), .C(n3780), .D(n3789), .Y(n3781) );
  OAI21X1 U4513 ( .A(n1353), .B(n3782), .C(n3781), .Y(n2076) );
  AOI22X1 U4514 ( .A(\data_in<13> ), .B(n1127), .C(n3783), .D(n3789), .Y(n3784) );
  OAI21X1 U4515 ( .A(n1353), .B(n3785), .C(n3784), .Y(n2077) );
  AOI22X1 U4516 ( .A(\data_in<14> ), .B(n1127), .C(n3786), .D(n3789), .Y(n3787) );
  OAI21X1 U4517 ( .A(n1353), .B(n3788), .C(n3787), .Y(n2078) );
  AOI22X1 U4518 ( .A(\data_in<15> ), .B(n1127), .C(n3790), .D(n3789), .Y(n3791) );
  OAI21X1 U4519 ( .A(n1353), .B(n3792), .C(n3791), .Y(n2079) );
  OAI21X1 U4520 ( .A(n3793), .B(n1418), .C(n1530), .Y(n3817) );
  AOI22X1 U4521 ( .A(\data_in<8> ), .B(n1128), .C(n3796), .D(n3817), .Y(n3797)
         );
  OAI21X1 U4522 ( .A(n1355), .B(n3798), .C(n3797), .Y(n2080) );
  AOI22X1 U4523 ( .A(\data_in<9> ), .B(n1128), .C(n3799), .D(n3817), .Y(n3800)
         );
  OAI21X1 U4524 ( .A(n1355), .B(n3801), .C(n3800), .Y(n2081) );
  AOI22X1 U4525 ( .A(\data_in<10> ), .B(n1128), .C(n3802), .D(n3817), .Y(n3803) );
  OAI21X1 U4526 ( .A(n1355), .B(n3804), .C(n3803), .Y(n2082) );
  AOI22X1 U4527 ( .A(\data_in<11> ), .B(n1128), .C(n3805), .D(n3817), .Y(n3806) );
  OAI21X1 U4528 ( .A(n1355), .B(n3807), .C(n3806), .Y(n2083) );
  AOI22X1 U4529 ( .A(\data_in<12> ), .B(n1128), .C(n3808), .D(n3817), .Y(n3809) );
  OAI21X1 U4530 ( .A(n1355), .B(n3810), .C(n3809), .Y(n2084) );
  AOI22X1 U4531 ( .A(\data_in<13> ), .B(n1128), .C(n3811), .D(n3817), .Y(n3812) );
  OAI21X1 U4532 ( .A(n1355), .B(n3813), .C(n3812), .Y(n2085) );
  AOI22X1 U4533 ( .A(\data_in<14> ), .B(n1128), .C(n3814), .D(n3817), .Y(n3815) );
  OAI21X1 U4534 ( .A(n1355), .B(n3816), .C(n3815), .Y(n2086) );
  AOI22X1 U4535 ( .A(\data_in<15> ), .B(n1128), .C(n3818), .D(n3817), .Y(n3819) );
  OAI21X1 U4536 ( .A(n1355), .B(n3820), .C(n3819), .Y(n2087) );
  OAI21X1 U4537 ( .A(n804), .B(n1418), .C(n4496), .Y(n3843) );
  AOI22X1 U4538 ( .A(\data_in<8> ), .B(n1129), .C(n3822), .D(n3843), .Y(n3823)
         );
  OAI21X1 U4539 ( .A(n1357), .B(n3824), .C(n3823), .Y(n2088) );
  AOI22X1 U4540 ( .A(\data_in<9> ), .B(n1129), .C(n3825), .D(n3843), .Y(n3826)
         );
  OAI21X1 U4541 ( .A(n1357), .B(n3827), .C(n3826), .Y(n2089) );
  AOI22X1 U4542 ( .A(\data_in<10> ), .B(n1129), .C(n3828), .D(n3843), .Y(n3829) );
  OAI21X1 U4543 ( .A(n1357), .B(n3830), .C(n3829), .Y(n2090) );
  AOI22X1 U4544 ( .A(\data_in<11> ), .B(n1129), .C(n3831), .D(n3843), .Y(n3832) );
  OAI21X1 U4545 ( .A(n1357), .B(n3833), .C(n3832), .Y(n2091) );
  AOI22X1 U4546 ( .A(\data_in<12> ), .B(n1129), .C(n3834), .D(n3843), .Y(n3835) );
  OAI21X1 U4547 ( .A(n1357), .B(n3836), .C(n3835), .Y(n2092) );
  AOI22X1 U4548 ( .A(\data_in<13> ), .B(n1129), .C(n3837), .D(n3843), .Y(n3838) );
  OAI21X1 U4549 ( .A(n1357), .B(n3839), .C(n3838), .Y(n2093) );
  AOI22X1 U4550 ( .A(\data_in<14> ), .B(n1129), .C(n3840), .D(n3843), .Y(n3841) );
  OAI21X1 U4551 ( .A(n1357), .B(n3842), .C(n3841), .Y(n2094) );
  AOI22X1 U4552 ( .A(\data_in<15> ), .B(n1129), .C(n3844), .D(n3843), .Y(n3845) );
  OAI21X1 U4553 ( .A(n1357), .B(n3846), .C(n3845), .Y(n2095) );
  OAI21X1 U4554 ( .A(n804), .B(n1507), .C(n1530), .Y(n3869) );
  AOI22X1 U4555 ( .A(\data_in<8> ), .B(n1130), .C(n3848), .D(n3869), .Y(n3849)
         );
  OAI21X1 U4556 ( .A(n1359), .B(n3850), .C(n3849), .Y(n2096) );
  AOI22X1 U4557 ( .A(\data_in<9> ), .B(n1130), .C(n3851), .D(n3869), .Y(n3852)
         );
  OAI21X1 U4558 ( .A(n1359), .B(n3853), .C(n3852), .Y(n2097) );
  AOI22X1 U4559 ( .A(\data_in<10> ), .B(n1130), .C(n3854), .D(n3869), .Y(n3855) );
  OAI21X1 U4560 ( .A(n1359), .B(n3856), .C(n3855), .Y(n2098) );
  AOI22X1 U4561 ( .A(\data_in<11> ), .B(n1130), .C(n3857), .D(n3869), .Y(n3858) );
  OAI21X1 U4562 ( .A(n1359), .B(n3859), .C(n3858), .Y(n2099) );
  AOI22X1 U4563 ( .A(\data_in<12> ), .B(n1130), .C(n3860), .D(n3869), .Y(n3861) );
  OAI21X1 U4564 ( .A(n1359), .B(n3862), .C(n3861), .Y(n2100) );
  AOI22X1 U4565 ( .A(\data_in<13> ), .B(n1130), .C(n3863), .D(n3869), .Y(n3864) );
  OAI21X1 U4566 ( .A(n1359), .B(n3865), .C(n3864), .Y(n2101) );
  AOI22X1 U4567 ( .A(\data_in<14> ), .B(n1130), .C(n3866), .D(n3869), .Y(n3867) );
  OAI21X1 U4568 ( .A(n1359), .B(n3868), .C(n3867), .Y(n2102) );
  AOI22X1 U4569 ( .A(\data_in<15> ), .B(n1130), .C(n3870), .D(n3869), .Y(n3871) );
  OAI21X1 U4570 ( .A(n1359), .B(n3872), .C(n3871), .Y(n2103) );
  OAI21X1 U4571 ( .A(n836), .B(n1507), .C(n1530), .Y(n3895) );
  AOI22X1 U4572 ( .A(\data_in<8> ), .B(n1131), .C(n3874), .D(n3895), .Y(n3875)
         );
  OAI21X1 U4573 ( .A(n1361), .B(n3876), .C(n3875), .Y(n2104) );
  AOI22X1 U4574 ( .A(\data_in<9> ), .B(n1131), .C(n3877), .D(n3895), .Y(n3878)
         );
  OAI21X1 U4575 ( .A(n1361), .B(n3879), .C(n3878), .Y(n2105) );
  AOI22X1 U4576 ( .A(\data_in<10> ), .B(n1131), .C(n3880), .D(n3895), .Y(n3881) );
  OAI21X1 U4577 ( .A(n1361), .B(n3882), .C(n3881), .Y(n2106) );
  AOI22X1 U4578 ( .A(\data_in<11> ), .B(n1131), .C(n3883), .D(n3895), .Y(n3884) );
  OAI21X1 U4579 ( .A(n1361), .B(n3885), .C(n3884), .Y(n2107) );
  AOI22X1 U4580 ( .A(\data_in<12> ), .B(n1131), .C(n3886), .D(n3895), .Y(n3887) );
  OAI21X1 U4581 ( .A(n1361), .B(n3888), .C(n3887), .Y(n2108) );
  AOI22X1 U4582 ( .A(\data_in<13> ), .B(n1131), .C(n3889), .D(n3895), .Y(n3890) );
  OAI21X1 U4583 ( .A(n1361), .B(n3891), .C(n3890), .Y(n2109) );
  AOI22X1 U4584 ( .A(\data_in<14> ), .B(n1131), .C(n3892), .D(n3895), .Y(n3893) );
  OAI21X1 U4585 ( .A(n1361), .B(n3894), .C(n3893), .Y(n2110) );
  AOI22X1 U4586 ( .A(\data_in<15> ), .B(n1131), .C(n3896), .D(n3895), .Y(n3897) );
  OAI21X1 U4587 ( .A(n1361), .B(n3898), .C(n3897), .Y(n2111) );
  OAI21X1 U4588 ( .A(n836), .B(n825), .C(n4496), .Y(n3922) );
  AOI22X1 U4589 ( .A(\data_in<8> ), .B(n1132), .C(n3901), .D(n3922), .Y(n3902)
         );
  OAI21X1 U4590 ( .A(n1363), .B(n3903), .C(n3902), .Y(n2112) );
  AOI22X1 U4591 ( .A(\data_in<9> ), .B(n1132), .C(n3904), .D(n3922), .Y(n3905)
         );
  OAI21X1 U4592 ( .A(n1363), .B(n3906), .C(n3905), .Y(n2113) );
  AOI22X1 U4593 ( .A(\data_in<10> ), .B(n1132), .C(n3907), .D(n3922), .Y(n3908) );
  OAI21X1 U4594 ( .A(n1363), .B(n3909), .C(n3908), .Y(n2114) );
  AOI22X1 U4595 ( .A(\data_in<11> ), .B(n1132), .C(n3910), .D(n3922), .Y(n3911) );
  OAI21X1 U4596 ( .A(n1363), .B(n3912), .C(n3911), .Y(n2115) );
  AOI22X1 U4597 ( .A(\data_in<12> ), .B(n1132), .C(n3913), .D(n3922), .Y(n3914) );
  OAI21X1 U4598 ( .A(n1363), .B(n3915), .C(n3914), .Y(n2116) );
  AOI22X1 U4599 ( .A(\data_in<13> ), .B(n1132), .C(n3916), .D(n3922), .Y(n3917) );
  OAI21X1 U4600 ( .A(n1363), .B(n3918), .C(n3917), .Y(n2117) );
  AOI22X1 U4601 ( .A(\data_in<14> ), .B(n1132), .C(n3919), .D(n3922), .Y(n3920) );
  OAI21X1 U4602 ( .A(n1363), .B(n3921), .C(n3920), .Y(n2118) );
  AOI22X1 U4603 ( .A(\data_in<15> ), .B(n1132), .C(n3923), .D(n3922), .Y(n3924) );
  OAI21X1 U4604 ( .A(n1363), .B(n3925), .C(n3924), .Y(n2119) );
  OAI21X1 U4605 ( .A(n3926), .B(n825), .C(n1530), .Y(n3949) );
  AOI22X1 U4606 ( .A(\data_in<8> ), .B(n1133), .C(n3928), .D(n3949), .Y(n3929)
         );
  OAI21X1 U4607 ( .A(n1365), .B(n3930), .C(n3929), .Y(n2120) );
  AOI22X1 U4608 ( .A(\data_in<9> ), .B(n1133), .C(n3931), .D(n3949), .Y(n3932)
         );
  OAI21X1 U4609 ( .A(n1365), .B(n3933), .C(n3932), .Y(n2121) );
  AOI22X1 U4610 ( .A(\data_in<10> ), .B(n1133), .C(n3934), .D(n3949), .Y(n3935) );
  OAI21X1 U4611 ( .A(n1365), .B(n3936), .C(n3935), .Y(n2122) );
  AOI22X1 U4612 ( .A(\data_in<11> ), .B(n1133), .C(n3937), .D(n3949), .Y(n3938) );
  OAI21X1 U4613 ( .A(n1365), .B(n3939), .C(n3938), .Y(n2123) );
  AOI22X1 U4614 ( .A(\data_in<12> ), .B(n1133), .C(n3940), .D(n3949), .Y(n3941) );
  OAI21X1 U4615 ( .A(n1365), .B(n3942), .C(n3941), .Y(n2124) );
  AOI22X1 U4616 ( .A(\data_in<13> ), .B(n1133), .C(n3943), .D(n3949), .Y(n3944) );
  OAI21X1 U4617 ( .A(n1365), .B(n3945), .C(n3944), .Y(n2125) );
  AOI22X1 U4618 ( .A(\data_in<14> ), .B(n1133), .C(n3946), .D(n3949), .Y(n3947) );
  OAI21X1 U4619 ( .A(n1365), .B(n3948), .C(n3947), .Y(n2126) );
  AOI22X1 U4620 ( .A(\data_in<15> ), .B(n1133), .C(n3950), .D(n3949), .Y(n3951) );
  OAI21X1 U4621 ( .A(n1365), .B(n3952), .C(n3951), .Y(n2127) );
  AOI22X1 U4622 ( .A(\data_in<8> ), .B(n1134), .C(n3953), .D(n1215), .Y(n3954)
         );
  OAI21X1 U4623 ( .A(n1367), .B(n3955), .C(n3954), .Y(n2128) );
  AOI22X1 U4624 ( .A(\data_in<9> ), .B(n1134), .C(n3956), .D(n1215), .Y(n3957)
         );
  OAI21X1 U4625 ( .A(n1367), .B(n3958), .C(n3957), .Y(n2129) );
  AOI22X1 U4626 ( .A(\data_in<10> ), .B(n1134), .C(n3959), .D(n1215), .Y(n3960) );
  OAI21X1 U4627 ( .A(n1367), .B(n3961), .C(n3960), .Y(n2130) );
  AOI22X1 U4628 ( .A(\data_in<11> ), .B(n1134), .C(n3962), .D(n1215), .Y(n3963) );
  OAI21X1 U4629 ( .A(n1367), .B(n3964), .C(n3963), .Y(n2131) );
  AOI22X1 U4630 ( .A(\data_in<12> ), .B(n1134), .C(n3965), .D(n1215), .Y(n3966) );
  OAI21X1 U4631 ( .A(n1367), .B(n3967), .C(n3966), .Y(n2132) );
  AOI22X1 U4632 ( .A(\data_in<13> ), .B(n1134), .C(n3968), .D(n1215), .Y(n3969) );
  OAI21X1 U4633 ( .A(n1367), .B(n3970), .C(n3969), .Y(n2133) );
  AOI22X1 U4634 ( .A(\data_in<14> ), .B(n1134), .C(n3971), .D(n1215), .Y(n3972) );
  OAI21X1 U4635 ( .A(n1367), .B(n3973), .C(n3972), .Y(n2134) );
  AOI22X1 U4636 ( .A(\data_in<15> ), .B(n1134), .C(n3974), .D(n1215), .Y(n3975) );
  OAI21X1 U4637 ( .A(n1367), .B(n3976), .C(n3975), .Y(n2135) );
  AOI22X1 U4638 ( .A(\data_in<8> ), .B(n1135), .C(n3977), .D(n1217), .Y(n3978)
         );
  OAI21X1 U4639 ( .A(n1369), .B(n3979), .C(n3978), .Y(n2136) );
  AOI22X1 U4640 ( .A(\data_in<9> ), .B(n1135), .C(n3980), .D(n1217), .Y(n3981)
         );
  OAI21X1 U4641 ( .A(n1369), .B(n3982), .C(n3981), .Y(n2137) );
  AOI22X1 U4642 ( .A(\data_in<10> ), .B(n1135), .C(n3983), .D(n1217), .Y(n3984) );
  OAI21X1 U4643 ( .A(n1369), .B(n3985), .C(n3984), .Y(n2138) );
  AOI22X1 U4644 ( .A(\data_in<11> ), .B(n1135), .C(n3986), .D(n1217), .Y(n3987) );
  OAI21X1 U4645 ( .A(n1369), .B(n3988), .C(n3987), .Y(n2139) );
  AOI22X1 U4646 ( .A(\data_in<12> ), .B(n1135), .C(n3989), .D(n1217), .Y(n3990) );
  OAI21X1 U4647 ( .A(n1369), .B(n3991), .C(n3990), .Y(n2140) );
  AOI22X1 U4648 ( .A(\data_in<13> ), .B(n1135), .C(n3992), .D(n1217), .Y(n3993) );
  OAI21X1 U4649 ( .A(n1369), .B(n3994), .C(n3993), .Y(n2141) );
  AOI22X1 U4650 ( .A(\data_in<14> ), .B(n1135), .C(n3995), .D(n1217), .Y(n3996) );
  OAI21X1 U4651 ( .A(n1369), .B(n3997), .C(n3996), .Y(n2142) );
  AOI22X1 U4652 ( .A(\data_in<15> ), .B(n1135), .C(n3998), .D(n1217), .Y(n3999) );
  OAI21X1 U4653 ( .A(n1369), .B(n4000), .C(n3999), .Y(n2143) );
  AOI22X1 U4654 ( .A(\data_in<8> ), .B(n1136), .C(n4001), .D(n1219), .Y(n4002)
         );
  OAI21X1 U4655 ( .A(n1371), .B(n4003), .C(n4002), .Y(n2144) );
  AOI22X1 U4656 ( .A(\data_in<9> ), .B(n1136), .C(n4004), .D(n1219), .Y(n4005)
         );
  OAI21X1 U4657 ( .A(n1371), .B(n4006), .C(n4005), .Y(n2145) );
  AOI22X1 U4658 ( .A(\data_in<10> ), .B(n1136), .C(n4007), .D(n1219), .Y(n4008) );
  OAI21X1 U4659 ( .A(n1371), .B(n4009), .C(n4008), .Y(n2146) );
  AOI22X1 U4660 ( .A(\data_in<11> ), .B(n1136), .C(n4010), .D(n1219), .Y(n4011) );
  OAI21X1 U4661 ( .A(n1371), .B(n4012), .C(n4011), .Y(n2147) );
  AOI22X1 U4662 ( .A(\data_in<12> ), .B(n1136), .C(n4013), .D(n1219), .Y(n4014) );
  OAI21X1 U4663 ( .A(n1371), .B(n4015), .C(n4014), .Y(n2148) );
  AOI22X1 U4664 ( .A(\data_in<13> ), .B(n1136), .C(n4016), .D(n1219), .Y(n4017) );
  OAI21X1 U4665 ( .A(n1371), .B(n4018), .C(n4017), .Y(n2149) );
  AOI22X1 U4666 ( .A(\data_in<14> ), .B(n1136), .C(n4019), .D(n1219), .Y(n4020) );
  OAI21X1 U4667 ( .A(n1371), .B(n4021), .C(n4020), .Y(n2150) );
  AOI22X1 U4668 ( .A(\data_in<15> ), .B(n1136), .C(n4022), .D(n1219), .Y(n4023) );
  OAI21X1 U4669 ( .A(n1371), .B(n4024), .C(n4023), .Y(n2151) );
  AOI22X1 U4670 ( .A(\data_in<8> ), .B(n1137), .C(n4026), .D(n1221), .Y(n4027)
         );
  OAI21X1 U4671 ( .A(n1373), .B(n4028), .C(n4027), .Y(n2152) );
  AOI22X1 U4672 ( .A(\data_in<9> ), .B(n1137), .C(n4029), .D(n1221), .Y(n4030)
         );
  OAI21X1 U4673 ( .A(n1373), .B(n4031), .C(n4030), .Y(n2153) );
  AOI22X1 U4674 ( .A(\data_in<10> ), .B(n1137), .C(n4032), .D(n1221), .Y(n4033) );
  OAI21X1 U4675 ( .A(n1373), .B(n4034), .C(n4033), .Y(n2154) );
  AOI22X1 U4676 ( .A(\data_in<11> ), .B(n1137), .C(n4035), .D(n1221), .Y(n4036) );
  OAI21X1 U4677 ( .A(n1373), .B(n4037), .C(n4036), .Y(n2155) );
  AOI22X1 U4678 ( .A(\data_in<12> ), .B(n1137), .C(n4038), .D(n1221), .Y(n4039) );
  OAI21X1 U4679 ( .A(n1373), .B(n4040), .C(n4039), .Y(n2156) );
  AOI22X1 U4680 ( .A(\data_in<13> ), .B(n1137), .C(n4041), .D(n1221), .Y(n4042) );
  OAI21X1 U4681 ( .A(n1373), .B(n4043), .C(n4042), .Y(n2157) );
  AOI22X1 U4682 ( .A(\data_in<14> ), .B(n1137), .C(n4044), .D(n1221), .Y(n4045) );
  OAI21X1 U4683 ( .A(n1373), .B(n4046), .C(n4045), .Y(n2158) );
  AOI22X1 U4684 ( .A(\data_in<15> ), .B(n1137), .C(n4047), .D(n1221), .Y(n4048) );
  OAI21X1 U4685 ( .A(n1373), .B(n4049), .C(n4048), .Y(n2159) );
  AOI22X1 U4686 ( .A(\data_in<8> ), .B(n1138), .C(n4051), .D(n1223), .Y(n4052)
         );
  OAI21X1 U4687 ( .A(n1375), .B(n4053), .C(n4052), .Y(n2160) );
  AOI22X1 U4688 ( .A(\data_in<9> ), .B(n1138), .C(n4054), .D(n1223), .Y(n4055)
         );
  OAI21X1 U4689 ( .A(n1375), .B(n4056), .C(n4055), .Y(n2161) );
  AOI22X1 U4690 ( .A(\data_in<10> ), .B(n1138), .C(n4057), .D(n1223), .Y(n4058) );
  OAI21X1 U4691 ( .A(n1375), .B(n4059), .C(n4058), .Y(n2162) );
  AOI22X1 U4692 ( .A(\data_in<11> ), .B(n1138), .C(n4060), .D(n1223), .Y(n4061) );
  OAI21X1 U4693 ( .A(n1375), .B(n4062), .C(n4061), .Y(n2163) );
  AOI22X1 U4694 ( .A(\data_in<12> ), .B(n1138), .C(n4063), .D(n1223), .Y(n4064) );
  OAI21X1 U4695 ( .A(n1375), .B(n4065), .C(n4064), .Y(n2164) );
  AOI22X1 U4696 ( .A(\data_in<13> ), .B(n1138), .C(n4066), .D(n1223), .Y(n4067) );
  OAI21X1 U4697 ( .A(n1375), .B(n4068), .C(n4067), .Y(n2165) );
  AOI22X1 U4698 ( .A(\data_in<14> ), .B(n1138), .C(n4069), .D(n1223), .Y(n4070) );
  OAI21X1 U4699 ( .A(n1375), .B(n4071), .C(n4070), .Y(n2166) );
  AOI22X1 U4700 ( .A(\data_in<15> ), .B(n1138), .C(n4072), .D(n1223), .Y(n4073) );
  OAI21X1 U4701 ( .A(n1375), .B(n4074), .C(n4073), .Y(n2167) );
  AOI22X1 U4702 ( .A(\data_in<8> ), .B(n1139), .C(n4076), .D(n1225), .Y(n4077)
         );
  OAI21X1 U4703 ( .A(n1377), .B(n4078), .C(n4077), .Y(n2168) );
  AOI22X1 U4704 ( .A(\data_in<9> ), .B(n1139), .C(n4079), .D(n1225), .Y(n4080)
         );
  OAI21X1 U4705 ( .A(n1377), .B(n4081), .C(n4080), .Y(n2169) );
  AOI22X1 U4706 ( .A(\data_in<10> ), .B(n1139), .C(n4082), .D(n1225), .Y(n4083) );
  OAI21X1 U4707 ( .A(n1377), .B(n4084), .C(n4083), .Y(n2170) );
  AOI22X1 U4708 ( .A(\data_in<11> ), .B(n1139), .C(n4085), .D(n1225), .Y(n4086) );
  OAI21X1 U4709 ( .A(n1377), .B(n4087), .C(n4086), .Y(n2171) );
  AOI22X1 U4710 ( .A(\data_in<12> ), .B(n1139), .C(n4088), .D(n1225), .Y(n4089) );
  OAI21X1 U4711 ( .A(n1377), .B(n4090), .C(n4089), .Y(n2172) );
  AOI22X1 U4712 ( .A(\data_in<13> ), .B(n1139), .C(n4091), .D(n1225), .Y(n4092) );
  OAI21X1 U4713 ( .A(n1377), .B(n4093), .C(n4092), .Y(n2173) );
  AOI22X1 U4714 ( .A(\data_in<14> ), .B(n1139), .C(n4094), .D(n1225), .Y(n4095) );
  OAI21X1 U4715 ( .A(n1377), .B(n4096), .C(n4095), .Y(n2174) );
  AOI22X1 U4716 ( .A(\data_in<15> ), .B(n1139), .C(n4097), .D(n1225), .Y(n4098) );
  OAI21X1 U4717 ( .A(n1377), .B(n4099), .C(n4098), .Y(n2175) );
  AOI22X1 U4718 ( .A(\data_in<8> ), .B(n1140), .C(n4100), .D(n1227), .Y(n4101)
         );
  OAI21X1 U4719 ( .A(n1379), .B(n4102), .C(n4101), .Y(n2176) );
  AOI22X1 U4720 ( .A(\data_in<9> ), .B(n1140), .C(n4103), .D(n1227), .Y(n4104)
         );
  OAI21X1 U4721 ( .A(n1379), .B(n4105), .C(n4104), .Y(n2177) );
  AOI22X1 U4722 ( .A(\data_in<10> ), .B(n1140), .C(n4106), .D(n1227), .Y(n4107) );
  OAI21X1 U4723 ( .A(n1379), .B(n4108), .C(n4107), .Y(n2178) );
  AOI22X1 U4724 ( .A(\data_in<11> ), .B(n1140), .C(n4109), .D(n1227), .Y(n4110) );
  OAI21X1 U4725 ( .A(n1379), .B(n4111), .C(n4110), .Y(n2179) );
  AOI22X1 U4726 ( .A(\data_in<12> ), .B(n1140), .C(n4112), .D(n1227), .Y(n4113) );
  OAI21X1 U4727 ( .A(n1379), .B(n4114), .C(n4113), .Y(n2180) );
  AOI22X1 U4728 ( .A(\data_in<13> ), .B(n1140), .C(n4115), .D(n1227), .Y(n4116) );
  OAI21X1 U4729 ( .A(n1379), .B(n4117), .C(n4116), .Y(n2181) );
  AOI22X1 U4730 ( .A(\data_in<14> ), .B(n1140), .C(n4118), .D(n1227), .Y(n4119) );
  OAI21X1 U4731 ( .A(n1379), .B(n4120), .C(n4119), .Y(n2182) );
  AOI22X1 U4732 ( .A(\data_in<15> ), .B(n1140), .C(n4121), .D(n1227), .Y(n4122) );
  OAI21X1 U4733 ( .A(n1379), .B(n4123), .C(n4122), .Y(n2183) );
  AOI22X1 U4734 ( .A(\data_in<8> ), .B(n1141), .C(n4124), .D(n1229), .Y(n4125)
         );
  OAI21X1 U4735 ( .A(n1381), .B(n4126), .C(n4125), .Y(n2184) );
  AOI22X1 U4736 ( .A(\data_in<9> ), .B(n1141), .C(n4127), .D(n1229), .Y(n4128)
         );
  OAI21X1 U4737 ( .A(n1381), .B(n4129), .C(n4128), .Y(n2185) );
  AOI22X1 U4738 ( .A(\data_in<10> ), .B(n1141), .C(n4130), .D(n1229), .Y(n4131) );
  OAI21X1 U4739 ( .A(n1381), .B(n4132), .C(n4131), .Y(n2186) );
  AOI22X1 U4740 ( .A(\data_in<11> ), .B(n1141), .C(n4133), .D(n1229), .Y(n4134) );
  OAI21X1 U4741 ( .A(n1381), .B(n4135), .C(n4134), .Y(n2187) );
  AOI22X1 U4742 ( .A(\data_in<12> ), .B(n1141), .C(n4136), .D(n1229), .Y(n4137) );
  OAI21X1 U4743 ( .A(n1381), .B(n4138), .C(n4137), .Y(n2188) );
  AOI22X1 U4744 ( .A(\data_in<13> ), .B(n1141), .C(n4139), .D(n1229), .Y(n4140) );
  OAI21X1 U4745 ( .A(n1381), .B(n4141), .C(n4140), .Y(n2189) );
  AOI22X1 U4746 ( .A(\data_in<14> ), .B(n1141), .C(n4142), .D(n1229), .Y(n4143) );
  OAI21X1 U4747 ( .A(n1381), .B(n4144), .C(n4143), .Y(n2190) );
  AOI22X1 U4748 ( .A(\data_in<15> ), .B(n1141), .C(n4145), .D(n1229), .Y(n4146) );
  OAI21X1 U4749 ( .A(n1381), .B(n4147), .C(n4146), .Y(n2191) );
  AOI22X1 U4750 ( .A(\data_in<8> ), .B(n1142), .C(n4150), .D(n1231), .Y(n4151)
         );
  OAI21X1 U4751 ( .A(n1383), .B(n4152), .C(n4151), .Y(n2192) );
  AOI22X1 U4752 ( .A(\data_in<9> ), .B(n1142), .C(n4153), .D(n1231), .Y(n4154)
         );
  OAI21X1 U4753 ( .A(n1383), .B(n4155), .C(n4154), .Y(n2193) );
  AOI22X1 U4754 ( .A(\data_in<10> ), .B(n1142), .C(n4156), .D(n1231), .Y(n4157) );
  OAI21X1 U4755 ( .A(n1383), .B(n4158), .C(n4157), .Y(n2194) );
  AOI22X1 U4756 ( .A(\data_in<11> ), .B(n1142), .C(n4159), .D(n1231), .Y(n4160) );
  OAI21X1 U4757 ( .A(n1383), .B(n4161), .C(n4160), .Y(n2195) );
  AOI22X1 U4758 ( .A(\data_in<12> ), .B(n1142), .C(n4162), .D(n1231), .Y(n4163) );
  OAI21X1 U4759 ( .A(n1383), .B(n4164), .C(n4163), .Y(n2196) );
  AOI22X1 U4760 ( .A(\data_in<13> ), .B(n1142), .C(n4165), .D(n1231), .Y(n4166) );
  OAI21X1 U4761 ( .A(n1383), .B(n4167), .C(n4166), .Y(n2197) );
  AOI22X1 U4762 ( .A(\data_in<14> ), .B(n1142), .C(n4168), .D(n1231), .Y(n4169) );
  OAI21X1 U4763 ( .A(n1383), .B(n4170), .C(n4169), .Y(n2198) );
  AOI22X1 U4764 ( .A(\data_in<15> ), .B(n1142), .C(n4171), .D(n1231), .Y(n4172) );
  OAI21X1 U4765 ( .A(n1383), .B(n4173), .C(n4172), .Y(n2199) );
  AOI22X1 U4766 ( .A(\data_in<8> ), .B(n1143), .C(n4174), .D(n1233), .Y(n4175)
         );
  OAI21X1 U4767 ( .A(n1385), .B(n4176), .C(n4175), .Y(n2200) );
  AOI22X1 U4768 ( .A(\data_in<9> ), .B(n1143), .C(n4177), .D(n1233), .Y(n4178)
         );
  OAI21X1 U4769 ( .A(n1385), .B(n4179), .C(n4178), .Y(n2201) );
  AOI22X1 U4770 ( .A(\data_in<10> ), .B(n1143), .C(n4180), .D(n1233), .Y(n4181) );
  OAI21X1 U4771 ( .A(n1385), .B(n4182), .C(n4181), .Y(n2202) );
  AOI22X1 U4772 ( .A(\data_in<11> ), .B(n1143), .C(n4183), .D(n1233), .Y(n4184) );
  OAI21X1 U4773 ( .A(n1385), .B(n4185), .C(n4184), .Y(n2203) );
  AOI22X1 U4774 ( .A(\data_in<12> ), .B(n1143), .C(n4186), .D(n1233), .Y(n4187) );
  OAI21X1 U4775 ( .A(n1385), .B(n4188), .C(n4187), .Y(n2204) );
  AOI22X1 U4776 ( .A(\data_in<13> ), .B(n1143), .C(n4189), .D(n1233), .Y(n4190) );
  OAI21X1 U4777 ( .A(n1385), .B(n4191), .C(n4190), .Y(n2205) );
  AOI22X1 U4778 ( .A(\data_in<14> ), .B(n1143), .C(n4192), .D(n1233), .Y(n4193) );
  OAI21X1 U4779 ( .A(n1385), .B(n4194), .C(n4193), .Y(n2206) );
  AOI22X1 U4780 ( .A(\data_in<15> ), .B(n1143), .C(n4195), .D(n1233), .Y(n4196) );
  OAI21X1 U4781 ( .A(n1385), .B(n4197), .C(n4196), .Y(n2207) );
  AOI22X1 U4782 ( .A(\data_in<8> ), .B(n1144), .C(n4200), .D(n1235), .Y(n4201)
         );
  OAI21X1 U4783 ( .A(n1387), .B(n4202), .C(n4201), .Y(n2208) );
  AOI22X1 U4784 ( .A(\data_in<9> ), .B(n1144), .C(n4203), .D(n1235), .Y(n4204)
         );
  OAI21X1 U4785 ( .A(n1387), .B(n4205), .C(n4204), .Y(n2209) );
  AOI22X1 U4786 ( .A(\data_in<10> ), .B(n1144), .C(n4206), .D(n1235), .Y(n4207) );
  OAI21X1 U4787 ( .A(n1387), .B(n4208), .C(n4207), .Y(n2210) );
  AOI22X1 U4788 ( .A(\data_in<11> ), .B(n1144), .C(n4209), .D(n1235), .Y(n4210) );
  OAI21X1 U4789 ( .A(n1387), .B(n4211), .C(n4210), .Y(n2211) );
  AOI22X1 U4790 ( .A(\data_in<12> ), .B(n1144), .C(n4212), .D(n1235), .Y(n4213) );
  OAI21X1 U4791 ( .A(n1387), .B(n4214), .C(n4213), .Y(n2212) );
  AOI22X1 U4792 ( .A(\data_in<13> ), .B(n1144), .C(n4215), .D(n1235), .Y(n4216) );
  OAI21X1 U4793 ( .A(n1387), .B(n4217), .C(n4216), .Y(n2213) );
  AOI22X1 U4794 ( .A(\data_in<14> ), .B(n1144), .C(n4218), .D(n1235), .Y(n4219) );
  OAI21X1 U4795 ( .A(n1387), .B(n4220), .C(n4219), .Y(n2214) );
  AOI22X1 U4796 ( .A(\data_in<15> ), .B(n1144), .C(n4221), .D(n1235), .Y(n4222) );
  OAI21X1 U4797 ( .A(n1387), .B(n4223), .C(n4222), .Y(n2215) );
  AOI22X1 U4798 ( .A(\data_in<8> ), .B(n1145), .C(n4224), .D(n1237), .Y(n4225)
         );
  OAI21X1 U4799 ( .A(n1389), .B(n4226), .C(n4225), .Y(n2216) );
  AOI22X1 U4800 ( .A(\data_in<9> ), .B(n1145), .C(n4227), .D(n1237), .Y(n4228)
         );
  OAI21X1 U4801 ( .A(n1389), .B(n4229), .C(n4228), .Y(n2217) );
  AOI22X1 U4802 ( .A(\data_in<10> ), .B(n1145), .C(n4230), .D(n1237), .Y(n4231) );
  OAI21X1 U4803 ( .A(n1389), .B(n4232), .C(n4231), .Y(n2218) );
  AOI22X1 U4804 ( .A(\data_in<11> ), .B(n1145), .C(n4233), .D(n1237), .Y(n4234) );
  OAI21X1 U4805 ( .A(n1389), .B(n4235), .C(n4234), .Y(n2219) );
  AOI22X1 U4806 ( .A(\data_in<12> ), .B(n1145), .C(n4236), .D(n1237), .Y(n4237) );
  OAI21X1 U4807 ( .A(n1389), .B(n4238), .C(n4237), .Y(n2220) );
  AOI22X1 U4808 ( .A(\data_in<13> ), .B(n1145), .C(n4239), .D(n1237), .Y(n4240) );
  OAI21X1 U4809 ( .A(n1389), .B(n4241), .C(n4240), .Y(n2221) );
  AOI22X1 U4810 ( .A(\data_in<14> ), .B(n1145), .C(n4242), .D(n1237), .Y(n4243) );
  OAI21X1 U4811 ( .A(n1389), .B(n4244), .C(n4243), .Y(n2222) );
  AOI22X1 U4812 ( .A(\data_in<15> ), .B(n1145), .C(n4245), .D(n1237), .Y(n4246) );
  OAI21X1 U4813 ( .A(n1389), .B(n4247), .C(n4246), .Y(n2223) );
  AOI22X1 U4814 ( .A(\data_in<8> ), .B(n1146), .C(n4248), .D(n1239), .Y(n4249)
         );
  OAI21X1 U4815 ( .A(n1391), .B(n4250), .C(n4249), .Y(n2224) );
  AOI22X1 U4816 ( .A(\data_in<9> ), .B(n1146), .C(n4251), .D(n1239), .Y(n4252)
         );
  OAI21X1 U4817 ( .A(n1391), .B(n4253), .C(n4252), .Y(n2225) );
  AOI22X1 U4818 ( .A(\data_in<10> ), .B(n1146), .C(n4254), .D(n1239), .Y(n4255) );
  OAI21X1 U4819 ( .A(n1391), .B(n4256), .C(n4255), .Y(n2226) );
  AOI22X1 U4820 ( .A(\data_in<11> ), .B(n1146), .C(n4257), .D(n1239), .Y(n4258) );
  OAI21X1 U4821 ( .A(n1391), .B(n4259), .C(n4258), .Y(n2227) );
  AOI22X1 U4822 ( .A(\data_in<12> ), .B(n1146), .C(n4260), .D(n1239), .Y(n4261) );
  OAI21X1 U4823 ( .A(n1391), .B(n4262), .C(n4261), .Y(n2228) );
  AOI22X1 U4824 ( .A(\data_in<13> ), .B(n1146), .C(n4263), .D(n1239), .Y(n4264) );
  OAI21X1 U4825 ( .A(n1391), .B(n4265), .C(n4264), .Y(n2229) );
  AOI22X1 U4826 ( .A(\data_in<14> ), .B(n1146), .C(n4266), .D(n1239), .Y(n4267) );
  OAI21X1 U4827 ( .A(n1391), .B(n4268), .C(n4267), .Y(n2230) );
  AOI22X1 U4828 ( .A(\data_in<15> ), .B(n1146), .C(n4269), .D(n1239), .Y(n4270) );
  OAI21X1 U4829 ( .A(n1391), .B(n4271), .C(n4270), .Y(n2231) );
  AOI22X1 U4830 ( .A(\data_in<8> ), .B(n1147), .C(n4273), .D(n1241), .Y(n4274)
         );
  OAI21X1 U4831 ( .A(n1393), .B(n4275), .C(n4274), .Y(n2232) );
  AOI22X1 U4832 ( .A(\data_in<9> ), .B(n1147), .C(n4276), .D(n1241), .Y(n4277)
         );
  OAI21X1 U4833 ( .A(n1393), .B(n4278), .C(n4277), .Y(n2233) );
  AOI22X1 U4834 ( .A(\data_in<10> ), .B(n1147), .C(n4279), .D(n1241), .Y(n4280) );
  OAI21X1 U4835 ( .A(n1393), .B(n4281), .C(n4280), .Y(n2234) );
  AOI22X1 U4836 ( .A(\data_in<11> ), .B(n1147), .C(n4282), .D(n1241), .Y(n4283) );
  OAI21X1 U4837 ( .A(n1393), .B(n4284), .C(n4283), .Y(n2235) );
  AOI22X1 U4838 ( .A(\data_in<12> ), .B(n1147), .C(n4285), .D(n1241), .Y(n4286) );
  OAI21X1 U4839 ( .A(n1393), .B(n4287), .C(n4286), .Y(n2236) );
  AOI22X1 U4840 ( .A(\data_in<13> ), .B(n1147), .C(n4288), .D(n1241), .Y(n4289) );
  OAI21X1 U4841 ( .A(n1393), .B(n4290), .C(n4289), .Y(n2237) );
  AOI22X1 U4842 ( .A(\data_in<14> ), .B(n1147), .C(n4291), .D(n1241), .Y(n4292) );
  OAI21X1 U4843 ( .A(n1393), .B(n4293), .C(n4292), .Y(n2238) );
  AOI22X1 U4844 ( .A(\data_in<15> ), .B(n1147), .C(n4294), .D(n1241), .Y(n4295) );
  OAI21X1 U4845 ( .A(n1393), .B(n4296), .C(n4295), .Y(n2239) );
  AOI22X1 U4846 ( .A(\data_in<8> ), .B(n1148), .C(n4298), .D(n1243), .Y(n4299)
         );
  OAI21X1 U4847 ( .A(n1395), .B(n4300), .C(n4299), .Y(n2240) );
  AOI22X1 U4848 ( .A(\data_in<9> ), .B(n1148), .C(n4301), .D(n1243), .Y(n4302)
         );
  OAI21X1 U4849 ( .A(n1395), .B(n4303), .C(n4302), .Y(n2241) );
  AOI22X1 U4850 ( .A(\data_in<10> ), .B(n1148), .C(n4304), .D(n1243), .Y(n4305) );
  OAI21X1 U4851 ( .A(n1395), .B(n4306), .C(n4305), .Y(n2242) );
  AOI22X1 U4852 ( .A(\data_in<11> ), .B(n1148), .C(n4307), .D(n1243), .Y(n4308) );
  OAI21X1 U4853 ( .A(n1395), .B(n4309), .C(n4308), .Y(n2243) );
  AOI22X1 U4854 ( .A(\data_in<12> ), .B(n1148), .C(n4310), .D(n1243), .Y(n4311) );
  OAI21X1 U4855 ( .A(n1395), .B(n4312), .C(n4311), .Y(n2244) );
  AOI22X1 U4856 ( .A(\data_in<13> ), .B(n1148), .C(n4313), .D(n1243), .Y(n4314) );
  OAI21X1 U4857 ( .A(n1395), .B(n4315), .C(n4314), .Y(n2245) );
  AOI22X1 U4858 ( .A(\data_in<14> ), .B(n1148), .C(n4316), .D(n1243), .Y(n4317) );
  OAI21X1 U4859 ( .A(n1395), .B(n4318), .C(n4317), .Y(n2246) );
  AOI22X1 U4860 ( .A(\data_in<15> ), .B(n1148), .C(n4319), .D(n1243), .Y(n4320) );
  OAI21X1 U4861 ( .A(n1395), .B(n4321), .C(n4320), .Y(n2247) );
  AOI22X1 U4862 ( .A(\data_in<8> ), .B(n1149), .C(n4322), .D(n1245), .Y(n4323)
         );
  OAI21X1 U4863 ( .A(n1397), .B(n4324), .C(n4323), .Y(n2248) );
  AOI22X1 U4864 ( .A(\data_in<9> ), .B(n1149), .C(n4325), .D(n1245), .Y(n4326)
         );
  OAI21X1 U4865 ( .A(n1397), .B(n4327), .C(n4326), .Y(n2249) );
  AOI22X1 U4866 ( .A(\data_in<10> ), .B(n1149), .C(n4328), .D(n1245), .Y(n4329) );
  OAI21X1 U4867 ( .A(n1397), .B(n4330), .C(n4329), .Y(n2250) );
  AOI22X1 U4868 ( .A(\data_in<11> ), .B(n1149), .C(n4331), .D(n1245), .Y(n4332) );
  OAI21X1 U4869 ( .A(n1397), .B(n4333), .C(n4332), .Y(n2251) );
  AOI22X1 U4870 ( .A(\data_in<12> ), .B(n1149), .C(n4334), .D(n1245), .Y(n4335) );
  OAI21X1 U4871 ( .A(n1397), .B(n4336), .C(n4335), .Y(n2252) );
  AOI22X1 U4872 ( .A(\data_in<13> ), .B(n1149), .C(n4337), .D(n1245), .Y(n4338) );
  OAI21X1 U4873 ( .A(n1397), .B(n4339), .C(n4338), .Y(n2253) );
  AOI22X1 U4874 ( .A(\data_in<14> ), .B(n1149), .C(n4340), .D(n1245), .Y(n4341) );
  OAI21X1 U4875 ( .A(n1397), .B(n4342), .C(n4341), .Y(n2254) );
  AOI22X1 U4876 ( .A(\data_in<15> ), .B(n1149), .C(n4343), .D(n1245), .Y(n4344) );
  OAI21X1 U4877 ( .A(n1397), .B(n4345), .C(n4344), .Y(n2255) );
  AOI22X1 U4878 ( .A(\data_in<8> ), .B(n1150), .C(n4347), .D(n1247), .Y(n4348)
         );
  OAI21X1 U4879 ( .A(n1399), .B(n4349), .C(n4348), .Y(n2256) );
  AOI22X1 U4880 ( .A(\data_in<9> ), .B(n1150), .C(n4350), .D(n1247), .Y(n4351)
         );
  OAI21X1 U4881 ( .A(n1399), .B(n4352), .C(n4351), .Y(n2257) );
  AOI22X1 U4882 ( .A(\data_in<10> ), .B(n1150), .C(n4353), .D(n1247), .Y(n4354) );
  OAI21X1 U4883 ( .A(n1399), .B(n4355), .C(n4354), .Y(n2258) );
  AOI22X1 U4884 ( .A(\data_in<11> ), .B(n1150), .C(n4356), .D(n1247), .Y(n4357) );
  OAI21X1 U4885 ( .A(n1399), .B(n4358), .C(n4357), .Y(n2259) );
  AOI22X1 U4886 ( .A(\data_in<12> ), .B(n1150), .C(n4359), .D(n1247), .Y(n4360) );
  OAI21X1 U4887 ( .A(n1399), .B(n4361), .C(n4360), .Y(n2260) );
  AOI22X1 U4888 ( .A(\data_in<13> ), .B(n1150), .C(n4362), .D(n1247), .Y(n4363) );
  OAI21X1 U4889 ( .A(n1399), .B(n4364), .C(n4363), .Y(n2261) );
  AOI22X1 U4890 ( .A(\data_in<14> ), .B(n1150), .C(n4365), .D(n1247), .Y(n4366) );
  OAI21X1 U4891 ( .A(n1399), .B(n4367), .C(n4366), .Y(n2262) );
  AOI22X1 U4892 ( .A(\data_in<15> ), .B(n1150), .C(n4368), .D(n1247), .Y(n4369) );
  OAI21X1 U4893 ( .A(n1399), .B(n4370), .C(n4369), .Y(n2263) );
  AOI22X1 U4894 ( .A(\data_in<8> ), .B(n1151), .C(n4372), .D(n1249), .Y(n4373)
         );
  OAI21X1 U4895 ( .A(n1401), .B(n4374), .C(n4373), .Y(n2264) );
  AOI22X1 U4896 ( .A(\data_in<9> ), .B(n1151), .C(n4375), .D(n1249), .Y(n4376)
         );
  OAI21X1 U4897 ( .A(n1401), .B(n4377), .C(n4376), .Y(n2265) );
  AOI22X1 U4898 ( .A(\data_in<10> ), .B(n1151), .C(n4378), .D(n1249), .Y(n4379) );
  OAI21X1 U4899 ( .A(n1401), .B(n4380), .C(n4379), .Y(n2266) );
  AOI22X1 U4900 ( .A(\data_in<11> ), .B(n1151), .C(n4381), .D(n1249), .Y(n4382) );
  OAI21X1 U4901 ( .A(n1401), .B(n4383), .C(n4382), .Y(n2267) );
  AOI22X1 U4902 ( .A(\data_in<12> ), .B(n1151), .C(n4384), .D(n1249), .Y(n4385) );
  OAI21X1 U4903 ( .A(n1401), .B(n4386), .C(n4385), .Y(n2268) );
  AOI22X1 U4904 ( .A(\data_in<13> ), .B(n1151), .C(n4387), .D(n1249), .Y(n4388) );
  OAI21X1 U4905 ( .A(n1401), .B(n4389), .C(n4388), .Y(n2269) );
  AOI22X1 U4906 ( .A(\data_in<14> ), .B(n1151), .C(n4390), .D(n1249), .Y(n4391) );
  OAI21X1 U4907 ( .A(n1401), .B(n4392), .C(n4391), .Y(n2270) );
  AOI22X1 U4908 ( .A(\data_in<15> ), .B(n1151), .C(n4393), .D(n1249), .Y(n4394) );
  OAI21X1 U4909 ( .A(n1401), .B(n4395), .C(n4394), .Y(n2271) );
  AOI22X1 U4910 ( .A(\data_in<8> ), .B(n1152), .C(n4397), .D(n1251), .Y(n4398)
         );
  OAI21X1 U4911 ( .A(n1403), .B(n4399), .C(n4398), .Y(n2272) );
  AOI22X1 U4912 ( .A(\data_in<9> ), .B(n1152), .C(n4400), .D(n1251), .Y(n4401)
         );
  OAI21X1 U4913 ( .A(n1403), .B(n4402), .C(n4401), .Y(n2273) );
  AOI22X1 U4914 ( .A(\data_in<10> ), .B(n1152), .C(n4403), .D(n1251), .Y(n4404) );
  OAI21X1 U4915 ( .A(n1403), .B(n4405), .C(n4404), .Y(n2274) );
  AOI22X1 U4916 ( .A(\data_in<11> ), .B(n1152), .C(n4406), .D(n1251), .Y(n4407) );
  OAI21X1 U4917 ( .A(n1403), .B(n4408), .C(n4407), .Y(n2275) );
  AOI22X1 U4918 ( .A(\data_in<12> ), .B(n1152), .C(n4409), .D(n1251), .Y(n4410) );
  OAI21X1 U4919 ( .A(n1403), .B(n4411), .C(n4410), .Y(n2276) );
  AOI22X1 U4920 ( .A(\data_in<13> ), .B(n1152), .C(n4412), .D(n1251), .Y(n4413) );
  OAI21X1 U4921 ( .A(n1403), .B(n4414), .C(n4413), .Y(n2277) );
  AOI22X1 U4922 ( .A(\data_in<14> ), .B(n1152), .C(n4415), .D(n1251), .Y(n4416) );
  OAI21X1 U4923 ( .A(n1403), .B(n4417), .C(n4416), .Y(n2278) );
  AOI22X1 U4924 ( .A(\data_in<15> ), .B(n1152), .C(n4418), .D(n1251), .Y(n4419) );
  OAI21X1 U4925 ( .A(n1403), .B(n4420), .C(n4419), .Y(n2279) );
  AOI22X1 U4926 ( .A(\data_in<8> ), .B(n1153), .C(n4421), .D(n1253), .Y(n4422)
         );
  OAI21X1 U4927 ( .A(n1405), .B(n4423), .C(n4422), .Y(n2280) );
  AOI22X1 U4928 ( .A(\data_in<9> ), .B(n1153), .C(n4424), .D(n1253), .Y(n4425)
         );
  OAI21X1 U4929 ( .A(n1405), .B(n4426), .C(n4425), .Y(n2281) );
  AOI22X1 U4930 ( .A(\data_in<10> ), .B(n1153), .C(n4427), .D(n1253), .Y(n4428) );
  OAI21X1 U4931 ( .A(n1405), .B(n4429), .C(n4428), .Y(n2282) );
  AOI22X1 U4932 ( .A(\data_in<11> ), .B(n1153), .C(n4430), .D(n1253), .Y(n4431) );
  OAI21X1 U4933 ( .A(n1405), .B(n4432), .C(n4431), .Y(n2283) );
  AOI22X1 U4934 ( .A(\data_in<12> ), .B(n1153), .C(n4433), .D(n1253), .Y(n4434) );
  OAI21X1 U4935 ( .A(n1405), .B(n4435), .C(n4434), .Y(n2284) );
  AOI22X1 U4936 ( .A(\data_in<13> ), .B(n1153), .C(n4436), .D(n1253), .Y(n4437) );
  OAI21X1 U4937 ( .A(n1405), .B(n4438), .C(n4437), .Y(n2285) );
  AOI22X1 U4938 ( .A(\data_in<14> ), .B(n1153), .C(n4439), .D(n1253), .Y(n4440) );
  OAI21X1 U4939 ( .A(n1405), .B(n4441), .C(n4440), .Y(n2286) );
  AOI22X1 U4940 ( .A(\data_in<15> ), .B(n1153), .C(n4442), .D(n1253), .Y(n4443) );
  OAI21X1 U4941 ( .A(n1405), .B(n4444), .C(n4443), .Y(n2287) );
  AOI22X1 U4942 ( .A(\data_in<8> ), .B(n1154), .C(n4446), .D(n1255), .Y(n4447)
         );
  OAI21X1 U4943 ( .A(n1407), .B(n4448), .C(n4447), .Y(n2288) );
  AOI22X1 U4944 ( .A(\data_in<9> ), .B(n1154), .C(n4449), .D(n1255), .Y(n4450)
         );
  OAI21X1 U4945 ( .A(n1407), .B(n4451), .C(n4450), .Y(n2289) );
  AOI22X1 U4946 ( .A(\data_in<10> ), .B(n1154), .C(n4452), .D(n1255), .Y(n4453) );
  OAI21X1 U4947 ( .A(n1407), .B(n4454), .C(n4453), .Y(n2290) );
  AOI22X1 U4948 ( .A(\data_in<11> ), .B(n1154), .C(n4455), .D(n1255), .Y(n4456) );
  OAI21X1 U4949 ( .A(n1407), .B(n4457), .C(n4456), .Y(n2291) );
  AOI22X1 U4950 ( .A(\data_in<12> ), .B(n1154), .C(n4458), .D(n1255), .Y(n4459) );
  OAI21X1 U4951 ( .A(n1407), .B(n4460), .C(n4459), .Y(n2292) );
  AOI22X1 U4952 ( .A(\data_in<13> ), .B(n1154), .C(n4461), .D(n1255), .Y(n4462) );
  OAI21X1 U4953 ( .A(n1407), .B(n4463), .C(n4462), .Y(n2293) );
  AOI22X1 U4954 ( .A(\data_in<14> ), .B(n1154), .C(n4464), .D(n1255), .Y(n4465) );
  OAI21X1 U4955 ( .A(n1407), .B(n4466), .C(n4465), .Y(n2294) );
  AOI22X1 U4956 ( .A(\data_in<15> ), .B(n1154), .C(n4467), .D(n1255), .Y(n4468) );
  OAI21X1 U4957 ( .A(n1407), .B(n4469), .C(n4468), .Y(n2295) );
  AOI22X1 U4958 ( .A(\data_in<8> ), .B(n1155), .C(n4472), .D(n1257), .Y(n4473)
         );
  OAI21X1 U4959 ( .A(n1409), .B(n4474), .C(n4473), .Y(n2296) );
  AOI22X1 U4960 ( .A(\data_in<9> ), .B(n1155), .C(n4475), .D(n1257), .Y(n4476)
         );
  OAI21X1 U4961 ( .A(n1409), .B(n4477), .C(n4476), .Y(n2297) );
  AOI22X1 U4962 ( .A(\data_in<10> ), .B(n1155), .C(n4478), .D(n1257), .Y(n4479) );
  OAI21X1 U4963 ( .A(n1409), .B(n4480), .C(n4479), .Y(n2298) );
  AOI22X1 U4964 ( .A(\data_in<11> ), .B(n1155), .C(n4481), .D(n1257), .Y(n4482) );
  OAI21X1 U4965 ( .A(n1409), .B(n4483), .C(n4482), .Y(n2299) );
  AOI22X1 U4966 ( .A(\data_in<12> ), .B(n1155), .C(n4484), .D(n1257), .Y(n4485) );
  OAI21X1 U4967 ( .A(n1409), .B(n4486), .C(n4485), .Y(n2300) );
  AOI22X1 U4968 ( .A(\data_in<13> ), .B(n1155), .C(n4487), .D(n1257), .Y(n4488) );
  OAI21X1 U4969 ( .A(n1409), .B(n4489), .C(n4488), .Y(n2301) );
  AOI22X1 U4970 ( .A(\data_in<14> ), .B(n1155), .C(n4490), .D(n1257), .Y(n4491) );
  OAI21X1 U4971 ( .A(n1409), .B(n4492), .C(n4491), .Y(n2302) );
  AOI22X1 U4972 ( .A(\data_in<15> ), .B(n1155), .C(n4493), .D(n1257), .Y(n4494) );
  OAI21X1 U4973 ( .A(n1409), .B(n4495), .C(n4494), .Y(n2303) );
  AOI22X1 U4974 ( .A(\data_in<8> ), .B(n1156), .C(n4497), .D(n1259), .Y(n4498)
         );
  OAI21X1 U4975 ( .A(n1411), .B(n4499), .C(n4498), .Y(n2304) );
  AOI22X1 U4976 ( .A(\data_in<9> ), .B(n1156), .C(n4500), .D(n1259), .Y(n4501)
         );
  OAI21X1 U4977 ( .A(n1411), .B(n4502), .C(n4501), .Y(n2305) );
  AOI22X1 U4978 ( .A(\data_in<10> ), .B(n1156), .C(n4503), .D(n1259), .Y(n4504) );
  OAI21X1 U4979 ( .A(n1411), .B(n4505), .C(n4504), .Y(n2306) );
  AOI22X1 U4980 ( .A(\data_in<11> ), .B(n1156), .C(n4506), .D(n1259), .Y(n4507) );
  OAI21X1 U4981 ( .A(n1411), .B(n4508), .C(n4507), .Y(n2307) );
  AOI22X1 U4982 ( .A(\data_in<12> ), .B(n1156), .C(n4509), .D(n1259), .Y(n4510) );
  OAI21X1 U4983 ( .A(n1411), .B(n4511), .C(n4510), .Y(n2308) );
  AOI22X1 U4984 ( .A(\data_in<13> ), .B(n1156), .C(n4512), .D(n1259), .Y(n4513) );
  OAI21X1 U4985 ( .A(n1411), .B(n4514), .C(n4513), .Y(n2309) );
  AOI22X1 U4986 ( .A(\data_in<14> ), .B(n1156), .C(n4515), .D(n1259), .Y(n4516) );
  OAI21X1 U4987 ( .A(n1411), .B(n4517), .C(n4516), .Y(n2310) );
  AOI22X1 U4988 ( .A(\data_in<15> ), .B(n1156), .C(n4518), .D(n1259), .Y(n4519) );
  OAI21X1 U4989 ( .A(n1411), .B(n4520), .C(n4519), .Y(n2311) );
  OAI21X1 U4990 ( .A(n4521), .B(n1282), .C(n1262), .Y(n4543) );
  NOR2X1 U4991 ( .A(n4543), .B(n4573), .Y(n4522) );
  AOI21X1 U4992 ( .A(\data_in<8> ), .B(n1157), .C(n4522), .Y(n4523) );
  OAI21X1 U4993 ( .A(n1413), .B(n4524), .C(n956), .Y(n2312) );
  NOR2X1 U4994 ( .A(n4543), .B(n4572), .Y(n4525) );
  AOI21X1 U4995 ( .A(\data_in<9> ), .B(n1157), .C(n4525), .Y(n4526) );
  OAI21X1 U4996 ( .A(n1413), .B(n4527), .C(n957), .Y(n2313) );
  NOR2X1 U4997 ( .A(n4543), .B(n4571), .Y(n4528) );
  AOI21X1 U4998 ( .A(\data_in<10> ), .B(n1157), .C(n4528), .Y(n4529) );
  OAI21X1 U4999 ( .A(n1413), .B(n4530), .C(n958), .Y(n2314) );
  NOR2X1 U5000 ( .A(n4543), .B(n4570), .Y(n4531) );
  AOI21X1 U5001 ( .A(\data_in<11> ), .B(n1157), .C(n4531), .Y(n4532) );
  OAI21X1 U5002 ( .A(n1413), .B(n4533), .C(n959), .Y(n2315) );
  NOR2X1 U5003 ( .A(n4543), .B(n4569), .Y(n4534) );
  AOI21X1 U5004 ( .A(\data_in<12> ), .B(n1157), .C(n4534), .Y(n4535) );
  OAI21X1 U5005 ( .A(n1413), .B(n4536), .C(n960), .Y(n2316) );
  NOR2X1 U5006 ( .A(n4543), .B(n4568), .Y(n4537) );
  AOI21X1 U5007 ( .A(\data_in<13> ), .B(n1157), .C(n4537), .Y(n4538) );
  OAI21X1 U5008 ( .A(n1413), .B(n4539), .C(n961), .Y(n2317) );
  NOR2X1 U5009 ( .A(n4543), .B(n4567), .Y(n4540) );
  AOI21X1 U5010 ( .A(\data_in<14> ), .B(n1157), .C(n4540), .Y(n4541) );
  OAI21X1 U5011 ( .A(n1413), .B(n4542), .C(n962), .Y(n2318) );
  NOR2X1 U5012 ( .A(n4543), .B(n4566), .Y(n4544) );
  AOI21X1 U5013 ( .A(\data_in<15> ), .B(n1157), .C(n4544), .Y(n4545) );
  OAI21X1 U5014 ( .A(n1413), .B(n4546), .C(n963), .Y(n2319) );
  MUX2X1 U5015 ( .B(n4565), .A(n4547), .S(n1261), .Y(n2320) );
  MUX2X1 U5016 ( .B(n4564), .A(n4548), .S(n1261), .Y(n2321) );
  MUX2X1 U5017 ( .B(n4563), .A(n4549), .S(n1261), .Y(n2322) );
  MUX2X1 U5018 ( .B(n4562), .A(n4550), .S(n1261), .Y(n2323) );
  MUX2X1 U5019 ( .B(n4561), .A(n4551), .S(n1261), .Y(n2324) );
  MUX2X1 U5020 ( .B(n4560), .A(n4552), .S(n1261), .Y(n2325) );
  MUX2X1 U5021 ( .B(n4559), .A(n4553), .S(n1261), .Y(n2326) );
  MUX2X1 U5022 ( .B(n4558), .A(n4554), .S(n1261), .Y(n2327) );
endmodule


module adder_2 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Overflow, Cout, .Sum({\Sum<15> , \Sum<14> , \Sum<13> , 
        \Sum<12> , \Sum<11> , \Sum<10> , \Sum<9> , \Sum<8> , \Sum<7> , 
        \Sum<6> , \Sum<5> , \Sum<4> , \Sum<3> , \Sum<2> , \Sum<1> , \Sum<0> })
 );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Overflow, Cout, \Sum<15> , \Sum<14> , \Sum<13> , \Sum<12> , \Sum<11> ,
         \Sum<10> , \Sum<9> , \Sum<8> , \Sum<7> , \Sum<6> , \Sum<5> , \Sum<4> ,
         \Sum<3> , \Sum<2> , \Sum<1> , \Sum<0> ;
  wire   c12, p12, g12, c8, p8, g8, c4, p4, g4, p0, g0, n1;

  FAX1 U1 ( .A(\B<15> ), .B(\A<15> ), .C(n1), .YC(), .YS(Overflow) );
  XOR2X1 U2 ( .A(\Sum<15> ), .B(Cout), .Y(n1) );
  cla_4_11 add1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(c12), .p(p12), .g(g12), .S({
        \Sum<15> , \Sum<14> , \Sum<13> , \Sum<12> }), .Cout() );
  cla_4_10 add2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(c8), .p(p8), .g(g8), .S({\Sum<11> , \Sum<10> , 
        \Sum<9> , \Sum<8> }), .Cout() );
  cla_4_9 add3 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(c4), .p(p4), .g(g4), .S({\Sum<7> , \Sum<6> , 
        \Sum<5> , \Sum<4> }), .Cout() );
  cla_4_8 add4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .p(p0), .g(g0), .S({\Sum<3> , \Sum<2> , 
        \Sum<1> , \Sum<0> }), .Cout() );
  groupcla_14 cla ( .p({p12, p8, p4, p0}), .g({g12, g8, g4, g0}), .Cin(Cin), 
        .c({Cout, c12, c8, c4}), .pg(), .gg() );
endmodule


module control ( .instr({\instr<4> , \instr<3> , \instr<2> , \instr<1> , 
        \instr<0> }), .func({\func<1> , \func<0> }), .regDst({\regDst<1> , 
        \regDst<0> }), regWrite, .whichImm({\whichImm<1> , \whichImm<0> }), 
        toExt, jump, jumpReg, branch, .branchOp({\branchOp<1> , \branchOp<0> }
        ), memRead, memWrite, memToReg, .ALUOp({\ALUOp<3> , \ALUOp<2> , 
        \ALUOp<1> , \ALUOp<0> }), ALUSrc, invSrc1, invSrc2, sub, halt, 
        passthrough, reverse, err );
  input \instr<4> , \instr<3> , \instr<2> , \instr<1> , \instr<0> , \func<1> ,
         \func<0> ;
  output \regDst<1> , \regDst<0> , regWrite, \whichImm<1> , \whichImm<0> ,
         toExt, jump, jumpReg, branch, \branchOp<1> , \branchOp<0> , memRead,
         memWrite, memToReg, \ALUOp<3> , \ALUOp<2> , \ALUOp<1> , \ALUOp<0> ,
         ALUSrc, invSrc1, invSrc2, sub, halt, passthrough, reverse, err;
  wire   n195, N7, N10, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n16, n18, n19, n20, n22, n24, n26, n27, n28, n29, n31, n32, n33,
         n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n110, n112, n113, n114, n115, n116, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n143, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n194;
  assign err = 1'b0;
  assign \regDst<1>  = N7;
  assign \regDst<0>  = N10;

  INVX1 U2 ( .A(n91), .Y(n1) );
  INVX1 U3 ( .A(n152), .Y(n2) );
  INVX4 U4 ( .A(n157), .Y(\ALUOp<2> ) );
  OR2X2 U5 ( .A(n4), .B(n46), .Y(\ALUOp<0> ) );
  INVX1 U6 ( .A(n169), .Y(n4) );
  INVX1 U7 ( .A(n115), .Y(n165) );
  INVX1 U8 ( .A(n24), .Y(\whichImm<1> ) );
  INVX1 U9 ( .A(memToReg), .Y(n143) );
  INVX1 U10 ( .A(n143), .Y(memRead) );
  AND2X2 U11 ( .A(n75), .B(n155), .Y(n5) );
  INVX1 U12 ( .A(n71), .Y(n6) );
  INVX4 U13 ( .A(\instr<4> ), .Y(n190) );
  MUX2X1 U14 ( .B(n62), .A(n38), .S(n125), .Y(n188) );
  INVX2 U15 ( .A(\instr<0> ), .Y(n141) );
  INVX1 U16 ( .A(n190), .Y(n7) );
  INVX1 U17 ( .A(\instr<2> ), .Y(n8) );
  AND2X2 U18 ( .A(n127), .B(n153), .Y(n9) );
  INVX1 U19 ( .A(n9), .Y(n65) );
  INVX2 U20 ( .A(\instr<1> ), .Y(n127) );
  INVX1 U21 ( .A(n11), .Y(n10) );
  INVX1 U22 ( .A(\func<0> ), .Y(n11) );
  INVX1 U23 ( .A(n11), .Y(n12) );
  INVX1 U24 ( .A(n1), .Y(n13) );
  AND2X2 U25 ( .A(n99), .B(n28), .Y(n14) );
  INVX1 U26 ( .A(n14), .Y(regWrite) );
  OR2X2 U27 ( .A(n74), .B(n119), .Y(n16) );
  INVX1 U28 ( .A(n16), .Y(reverse) );
  OR2X2 U29 ( .A(n93), .B(n51), .Y(n18) );
  INVX1 U30 ( .A(n18), .Y(n19) );
  AND2X2 U31 ( .A(n181), .B(n180), .Y(n20) );
  INVX1 U32 ( .A(n20), .Y(\ALUOp<3> ) );
  AND2X2 U33 ( .A(n50), .B(n45), .Y(n22) );
  INVX1 U34 ( .A(n22), .Y(\whichImm<0> ) );
  AND2X2 U35 ( .A(n43), .B(n188), .Y(n24) );
  OR2X2 U36 ( .A(n87), .B(n101), .Y(n26) );
  INVX1 U37 ( .A(n26), .Y(n27) );
  AND2X2 U38 ( .A(n114), .B(n95), .Y(n28) );
  OR2X2 U39 ( .A(n81), .B(n119), .Y(n29) );
  INVX1 U40 ( .A(n29), .Y(passthrough) );
  AND2X2 U41 ( .A(n126), .B(n160), .Y(n31) );
  AND2X2 U42 ( .A(n136), .B(n161), .Y(n32) );
  OR2X2 U43 ( .A(n88), .B(n120), .Y(n33) );
  INVX1 U44 ( .A(n33), .Y(n34) );
  AND2X2 U45 ( .A(n73), .B(n148), .Y(memToReg) );
  OR2X2 U46 ( .A(n93), .B(n154), .Y(n36) );
  OR2X2 U47 ( .A(n163), .B(n8), .Y(n37) );
  INVX1 U48 ( .A(n37), .Y(n38) );
  BUFX2 U49 ( .A(n170), .Y(n39) );
  BUFX2 U50 ( .A(n176), .Y(n40) );
  AND2X2 U51 ( .A(n161), .B(n91), .Y(n41) );
  INVX1 U52 ( .A(n41), .Y(n42) );
  BUFX2 U53 ( .A(n189), .Y(n43) );
  AND2X2 U54 ( .A(n48), .B(n158), .Y(n44) );
  INVX1 U55 ( .A(n44), .Y(n45) );
  AND2X2 U56 ( .A(n92), .B(n167), .Y(n46) );
  AND2X2 U57 ( .A(n141), .B(n150), .Y(n47) );
  INVX1 U58 ( .A(n47), .Y(n48) );
  AND2X2 U59 ( .A(n132), .B(n89), .Y(n49) );
  INVX1 U60 ( .A(n49), .Y(n50) );
  BUFX2 U61 ( .A(n171), .Y(n51) );
  AND2X2 U62 ( .A(n149), .B(n92), .Y(n52) );
  INVX1 U63 ( .A(n52), .Y(n53) );
  AND2X2 U64 ( .A(n190), .B(n156), .Y(n54) );
  INVX1 U65 ( .A(n54), .Y(n55) );
  BUFX2 U66 ( .A(n173), .Y(n56) );
  AND2X2 U67 ( .A(n10), .B(n91), .Y(n57) );
  INVX1 U68 ( .A(n57), .Y(n58) );
  OR2X2 U69 ( .A(n121), .B(n186), .Y(n59) );
  INVX1 U70 ( .A(n59), .Y(n60) );
  OR2X2 U71 ( .A(n186), .B(n147), .Y(n61) );
  INVX1 U72 ( .A(n61), .Y(n62) );
  AND2X2 U73 ( .A(n163), .B(n2), .Y(n63) );
  INVX1 U74 ( .A(n63), .Y(n64) );
  AND2X2 U75 ( .A(n165), .B(n164), .Y(n66) );
  INVX1 U76 ( .A(n66), .Y(n67) );
  AND2X2 U77 ( .A(n183), .B(n31), .Y(n68) );
  INVX1 U78 ( .A(n68), .Y(n69) );
  AND2X2 U79 ( .A(n182), .B(n31), .Y(n70) );
  INVX1 U80 ( .A(n70), .Y(n71) );
  INVX1 U81 ( .A(n70), .Y(n72) );
  AND2X2 U82 ( .A(n139), .B(n9), .Y(n73) );
  INVX1 U83 ( .A(n73), .Y(n74) );
  AND2X2 U84 ( .A(\func<1> ), .B(\func<0> ), .Y(n75) );
  INVX1 U85 ( .A(n75), .Y(n76) );
  AND2X2 U86 ( .A(n39), .B(n69), .Y(n77) );
  INVX1 U87 ( .A(n77), .Y(n78) );
  INVX1 U88 ( .A(n77), .Y(n79) );
  AND2X2 U89 ( .A(n182), .B(n9), .Y(n80) );
  INVX1 U90 ( .A(n80), .Y(n81) );
  INVX1 U91 ( .A(n80), .Y(n82) );
  AND2X2 U92 ( .A(n153), .B(n148), .Y(n83) );
  BUFX2 U93 ( .A(n178), .Y(n84) );
  INVX1 U94 ( .A(n84), .Y(n85) );
  INVX1 U95 ( .A(n84), .Y(jumpReg) );
  INVX1 U96 ( .A(n32), .Y(n87) );
  INVX1 U97 ( .A(n32), .Y(n88) );
  INVX2 U98 ( .A(n156), .Y(n151) );
  AND2X2 U99 ( .A(n134), .B(n190), .Y(n89) );
  INVX1 U100 ( .A(n190), .Y(n90) );
  INVX1 U101 ( .A(n152), .Y(n91) );
  INVX2 U102 ( .A(n141), .Y(n136) );
  AND2X2 U103 ( .A(n136), .B(n159), .Y(n92) );
  BUFX2 U104 ( .A(n161), .Y(n93) );
  AND2X2 U105 ( .A(n130), .B(n82), .Y(n94) );
  INVX1 U106 ( .A(n94), .Y(n95) );
  OR2X2 U107 ( .A(n118), .B(n136), .Y(n96) );
  INVX1 U108 ( .A(n96), .Y(n97) );
  AND2X2 U109 ( .A(n93), .B(n151), .Y(n98) );
  INVX1 U110 ( .A(n98), .Y(n99) );
  AND2X2 U111 ( .A(n126), .B(n163), .Y(n100) );
  INVX1 U112 ( .A(n100), .Y(n101) );
  AND2X2 U113 ( .A(n149), .B(n155), .Y(n102) );
  INVX1 U114 ( .A(n102), .Y(n103) );
  OR2X2 U115 ( .A(n183), .B(n136), .Y(n104) );
  INVX1 U116 ( .A(n104), .Y(n105) );
  INVX1 U117 ( .A(n174), .Y(n106) );
  INVX1 U118 ( .A(n106), .Y(n107) );
  OR2X2 U119 ( .A(n123), .B(n183), .Y(n108) );
  INVX1 U120 ( .A(n108), .Y(\branchOp<1> ) );
  INVX1 U121 ( .A(n195), .Y(n110) );
  INVX1 U122 ( .A(n110), .Y(memWrite) );
  INVX1 U123 ( .A(n83), .Y(n112) );
  AND2X2 U124 ( .A(n132), .B(n134), .Y(n113) );
  INVX1 U125 ( .A(n113), .Y(n114) );
  INVX1 U126 ( .A(n113), .Y(n115) );
  OR2X2 U127 ( .A(n123), .B(n182), .Y(n116) );
  INVX1 U128 ( .A(n116), .Y(\branchOp<0> ) );
  INVX1 U129 ( .A(n122), .Y(n118) );
  INVX1 U130 ( .A(n160), .Y(n119) );
  INVX1 U131 ( .A(n122), .Y(n120) );
  NOR3X1 U132 ( .A(n182), .B(n67), .C(n166), .Y(invSrc1) );
  INVX2 U133 ( .A(n125), .Y(n182) );
  INVX1 U134 ( .A(n124), .Y(n121) );
  AND2X2 U135 ( .A(n124), .B(n7), .Y(n122) );
  INVX1 U136 ( .A(n184), .Y(n194) );
  INVX1 U137 ( .A(branch), .Y(n123) );
  INVX1 U138 ( .A(n133), .Y(n124) );
  INVX4 U139 ( .A(n175), .Y(\ALUOp<1> ) );
  INVX1 U140 ( .A(n141), .Y(n125) );
  INVX1 U141 ( .A(n187), .Y(n126) );
  INVX1 U142 ( .A(n127), .Y(n128) );
  BUFX2 U143 ( .A(n194), .Y(branch) );
  BUFX2 U144 ( .A(n163), .Y(n130) );
  INVX1 U145 ( .A(n71), .Y(n179) );
  INVX1 U146 ( .A(n153), .Y(n131) );
  INVX1 U147 ( .A(n131), .Y(n132) );
  INVX1 U148 ( .A(\instr<2> ), .Y(n153) );
  INVX1 U149 ( .A(\instr<3> ), .Y(n133) );
  INVX1 U150 ( .A(n145), .Y(n134) );
  INVX1 U151 ( .A(n190), .Y(n135) );
  INVX1 U152 ( .A(n89), .Y(n137) );
  INVX1 U153 ( .A(n125), .Y(n138) );
  INVX1 U154 ( .A(n138), .Y(n139) );
  AND2X2 U155 ( .A(n89), .B(n132), .Y(n140) );
  INVX1 U156 ( .A(n186), .Y(n159) );
  BUFX2 U157 ( .A(invSrc1), .Y(sub) );
  INVX1 U158 ( .A(\instr<3> ), .Y(n145) );
  INVX1 U159 ( .A(n133), .Y(n146) );
  INVX1 U160 ( .A(n158), .Y(n147) );
  INVX1 U161 ( .A(n147), .Y(n148) );
  BUFX2 U162 ( .A(n146), .Y(n149) );
  AND2X2 U163 ( .A(n187), .B(\instr<1> ), .Y(n150) );
  INVX1 U164 ( .A(n150), .Y(n186) );
  INVX1 U165 ( .A(\func<1> ), .Y(n152) );
  AND2X2 U166 ( .A(n9), .B(n141), .Y(n185) );
  INVX1 U167 ( .A(\instr<2> ), .Y(n187) );
  INVX1 U168 ( .A(n128), .Y(n183) );
  BUFX2 U169 ( .A(n139), .Y(n154) );
  INVX1 U170 ( .A(n186), .Y(n155) );
  BUFX2 U171 ( .A(\instr<3> ), .Y(n162) );
  INVX1 U172 ( .A(n13), .Y(n172) );
  BUFX2 U173 ( .A(n128), .Y(n161) );
  OR2X2 U174 ( .A(n162), .B(n8), .Y(n156) );
  AND2X2 U175 ( .A(n40), .B(n177), .Y(n157) );
  AND2X2 U176 ( .A(\instr<4> ), .B(n145), .Y(n158) );
  INVX1 U177 ( .A(n158), .Y(n191) );
  AND2X2 U178 ( .A(n124), .B(n135), .Y(n160) );
  BUFX4 U179 ( .A(\instr<4> ), .Y(n163) );
  NOR3X1 U180 ( .A(n130), .B(n82), .C(n149), .Y(halt) );
  OAI21X1 U181 ( .A(n183), .B(n12), .C(n42), .Y(n166) );
  XNOR2X1 U182 ( .A(n161), .B(n163), .Y(n164) );
  AOI21X1 U183 ( .A(n90), .B(n58), .C(n53), .Y(invSrc2) );
  NAND3X1 U184 ( .A(n146), .B(n163), .C(n65), .Y(ALUSrc) );
  OAI21X1 U185 ( .A(n120), .B(n76), .C(n137), .Y(n167) );
  OAI21X1 U186 ( .A(n10), .B(n64), .C(n191), .Y(n168) );
  AOI21X1 U187 ( .A(n168), .B(n105), .C(n6), .Y(n169) );
  NAND3X1 U188 ( .A(n122), .B(n92), .C(n13), .Y(n170) );
  NAND3X1 U189 ( .A(n139), .B(n163), .C(n151), .Y(n171) );
  NAND3X1 U190 ( .A(n12), .B(n182), .C(n172), .Y(n173) );
  AOI21X1 U191 ( .A(n130), .B(n56), .C(n103), .Y(n174) );
  NOR3X1 U192 ( .A(n78), .B(n19), .C(n107), .Y(n175) );
  AND2X2 U193 ( .A(n69), .B(n72), .Y(n177) );
  AOI21X1 U194 ( .A(n97), .B(n5), .C(n27), .Y(n176) );
  NAND3X1 U195 ( .A(n136), .B(n151), .C(n190), .Y(n178) );
  NOR3X1 U196 ( .A(n85), .B(n140), .C(n79), .Y(n181) );
  NOR3X1 U197 ( .A(n83), .B(n34), .C(n179), .Y(n180) );
  AOI21X1 U198 ( .A(n87), .B(n36), .C(n112), .Y(n195) );
  NAND3X1 U199 ( .A(n126), .B(n162), .C(n190), .Y(n184) );
  NOR3X1 U200 ( .A(n154), .B(n156), .C(n130), .Y(jump) );
  MUX2X1 U201 ( .B(n60), .A(n151), .S(n163), .Y(toExt) );
  AOI21X1 U202 ( .A(n185), .B(n122), .C(n194), .Y(n189) );
  OAI21X1 U203 ( .A(n155), .B(n146), .C(n130), .Y(N10) );
  NAND3X1 U204 ( .A(n55), .B(n191), .C(n82), .Y(N7) );
endmodule


module rf ( .read1data({\read1data<15> , \read1data<14> , \read1data<13> , 
        \read1data<12> , \read1data<11> , \read1data<10> , \read1data<9> , 
        \read1data<8> , \read1data<7> , \read1data<6> , \read1data<5> , 
        \read1data<4> , \read1data<3> , \read1data<2> , \read1data<1> , 
        \read1data<0> }), .read2data({\read2data<15> , \read2data<14> , 
        \read2data<13> , \read2data<12> , \read2data<11> , \read2data<10> , 
        \read2data<9> , \read2data<8> , \read2data<7> , \read2data<6> , 
        \read2data<5> , \read2data<4> , \read2data<3> , \read2data<2> , 
        \read2data<1> , \read2data<0> }), err, clk, rst, .read1regsel({
        \read1regsel<2> , \read1regsel<1> , \read1regsel<0> }), .read2regsel({
        \read2regsel<2> , \read2regsel<1> , \read2regsel<0> }), .writeregsel({
        \writeregsel<2> , \writeregsel<1> , \writeregsel<0> }), .writedata({
        \writedata<15> , \writedata<14> , \writedata<13> , \writedata<12> , 
        \writedata<11> , \writedata<10> , \writedata<9> , \writedata<8> , 
        \writedata<7> , \writedata<6> , \writedata<5> , \writedata<4> , 
        \writedata<3> , \writedata<2> , \writedata<1> , \writedata<0> }), 
        write );
  input clk, rst, \read1regsel<2> , \read1regsel<1> , \read1regsel<0> ,
         \read2regsel<2> , \read2regsel<1> , \read2regsel<0> ,
         \writeregsel<2> , \writeregsel<1> , \writeregsel<0> , \writedata<15> ,
         \writedata<14> , \writedata<13> , \writedata<12> , \writedata<11> ,
         \writedata<10> , \writedata<9> , \writedata<8> , \writedata<7> ,
         \writedata<6> , \writedata<5> , \writedata<4> , \writedata<3> ,
         \writedata<2> , \writedata<1> , \writedata<0> , write;
  output \read1data<15> , \read1data<14> , \read1data<13> , \read1data<12> ,
         \read1data<11> , \read1data<10> , \read1data<9> , \read1data<8> ,
         \read1data<7> , \read1data<6> , \read1data<5> , \read1data<4> ,
         \read1data<3> , \read1data<2> , \read1data<1> , \read1data<0> ,
         \read2data<15> , \read2data<14> , \read2data<13> , \read2data<12> ,
         \read2data<11> , \read2data<10> , \read2data<9> , \read2data<8> ,
         \read2data<7> , \read2data<6> , \read2data<5> , \read2data<4> ,
         \read2data<3> , \read2data<2> , \read2data<1> , \read2data<0> , err;
  wire   \r7in<15> , \r7in<14> , \r7in<13> , \r7in<12> , \r7in<10> , \r7in<8> ,
         \r7in<5> , \r7in<4> , \r6in<15> , \r6in<14> , \r6in<13> , \r6in<12> ,
         \r6in<10> , \r6in<8> , \r6in<7> , \r6in<6> , \r6in<5> , \r6in<4> ,
         \r6in<2> , \r5in<15> , \r5in<14> , \r5in<13> , \r5in<12> , \r5in<10> ,
         \r5in<8> , \r5in<7> , \r5in<5> , \r5in<4> , \r5in<2> , \r4in<15> ,
         \r4in<14> , \r4in<13> , \r4in<12> , \r4in<10> , \r4in<8> , \r4in<7> ,
         \r4in<6> , \r4in<5> , \r4in<4> , \r4in<2> , \r3in<15> , \r3in<14> ,
         \r3in<13> , \r3in<12> , \r3in<8> , \r3in<7> , \r3in<5> , \r3in<4> ,
         \r2in<15> , \r2in<14> , \r2in<13> , \r2in<12> , \r2in<10> , \r2in<8> ,
         \r2in<7> , \r2in<6> , \r2in<5> , \r2in<4> , \r2in<2> , \r2in<1> ,
         \r2in<0> , \r1in<15> , \r1in<14> , \r1in<13> , \r1in<12> , \r1in<10> ,
         \r1in<8> , \r1in<7> , \r1in<6> , \r1in<5> , \r1in<4> , \r1in<1> ,
         \r1in<0> , \r0in<15> , \r0in<14> , \r0in<13> , \r0in<12> , \r0in<10> ,
         \r0in<8> , \r0in<7> , \r0in<6> , \r0in<5> , \r0in<4> , \r0in<0> , n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225;
  assign err = 1'b0;
  assign \read2data<0>  = 1'b0;
  assign \read2data<1>  = 1'b0;
  assign \read2data<2>  = 1'b0;
  assign \read2data<3>  = 1'b0;
  assign \read2data<4>  = 1'b0;
  assign \read2data<5>  = 1'b0;
  assign \read2data<6>  = 1'b0;
  assign \read2data<7>  = 1'b0;
  assign \read2data<8>  = 1'b0;
  assign \read2data<9>  = 1'b0;
  assign \read2data<10>  = 1'b0;
  assign \read2data<11>  = 1'b0;
  assign \read2data<12>  = 1'b0;
  assign \read2data<13>  = 1'b0;
  assign \read2data<14>  = 1'b0;
  assign \read2data<15>  = 1'b0;
  assign \read1data<0>  = 1'b0;
  assign \read1data<1>  = 1'b0;
  assign \read1data<2>  = 1'b0;
  assign \read1data<3>  = 1'b0;
  assign \read1data<4>  = 1'b0;
  assign \read1data<5>  = 1'b0;
  assign \read1data<6>  = 1'b0;
  assign \read1data<7>  = 1'b0;
  assign \read1data<8>  = 1'b0;
  assign \read1data<9>  = 1'b0;
  assign \read1data<10>  = 1'b0;
  assign \read1data<11>  = 1'b0;
  assign \read1data<12>  = 1'b0;
  assign \read1data<13>  = 1'b0;
  assign \read1data<14>  = 1'b0;
  assign \read1data<15>  = 1'b0;

  register_7 r7 ( .in({\r7in<15> , \r7in<14> , \r7in<13> , \r7in<12> , n128, 
        \r7in<10> , n130, \r7in<8> , n60, n58, \r7in<5> , \r7in<4> , n64, n70, 
        n66, n68}), .clk(clk), .rst(n213), .out({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  register_6 r6 ( .in({\r6in<15> , \r6in<14> , \r6in<13> , \r6in<12> , n124, 
        \r6in<10> , n126, \r6in<8> , \r6in<7> , \r6in<6> , \r6in<5> , 
        \r6in<4> , n86, \r6in<2> , n88, n92}), .clk(clk), .rst(n212), .out({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  register_5 r5 ( .in({\r5in<15> , \r5in<14> , \r5in<13> , \r5in<12> , n120, 
        \r5in<10> , n122, \r5in<8> , \r5in<7> , n38, \r5in<5> , \r5in<4> , n44, 
        \r5in<2> , n37, n78}), .clk(clk), .rst(n212), .out({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}) );
  register_4 r4 ( .in({\r4in<15> , \r4in<14> , \r4in<13> , \r4in<12> , n116, 
        \r4in<10> , n118, \r4in<8> , \r4in<7> , \r4in<6> , \r4in<5> , 
        \r4in<4> , n80, \r4in<2> , n82, n84}), .clk(clk), .rst(n212), .out({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  register_3 r3 ( .in({\r3in<15> , \r3in<14> , \r3in<13> , \r3in<12> , n112, 
        n143, n114, \r3in<8> , \r3in<7> , n62, \r3in<5> , \r3in<4> , n54, n76, 
        n72, n74}), .clk(clk), .rst(n212), .out({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  register_2 r2 ( .in({\r2in<15> , \r2in<14> , \r2in<13> , \r2in<12> , n108, 
        \r2in<10> , n110, \r2in<8> , \r2in<7> , \r2in<6> , \r2in<5> , 
        \r2in<4> , n98, \r2in<2> , \r2in<1> , \r2in<0> }), .clk(clk), .rst(
        n213), .out({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  register_1 r1 ( .in({\r1in<15> , \r1in<14> , \r1in<13> , \r1in<12> , n104, 
        \r1in<10> , n106, \r1in<8> , \r1in<7> , \r1in<6> , \r1in<5> , 
        \r1in<4> , n90, n96, \r1in<1> , \r1in<0> }), .clk(clk), .rst(n213), 
        .out({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  register_0 r0 ( .in({\r0in<15> , \r0in<14> , \r0in<13> , \r0in<12> , n100, 
        \r0in<10> , n102, \r0in<8> , \r0in<7> , \r0in<6> , \r0in<5> , 
        \r0in<4> , n56, n42, n94, \r0in<0> }), .clk(clk), .rst(n213), .out({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}) );
  INVX1 U34 ( .A(\writedata<9> ), .Y(n33) );
  INVX1 U35 ( .A(\writedata<10> ), .Y(n34) );
  INVX1 U36 ( .A(n34), .Y(n35) );
  INVX1 U37 ( .A(n209), .Y(n36) );
  AND2X1 U38 ( .A(n52), .B(n45), .Y(n37) );
  INVX4 U39 ( .A(n137), .Y(n45) );
  INVX2 U40 ( .A(n176), .Y(n225) );
  BUFX2 U41 ( .A(rst), .Y(n212) );
  BUFX2 U42 ( .A(rst), .Y(n213) );
  INVX1 U43 ( .A(write), .Y(n214) );
  INVX2 U44 ( .A(n170), .Y(n224) );
  INVX2 U45 ( .A(n166), .Y(n222) );
  INVX2 U46 ( .A(n155), .Y(n219) );
  INVX2 U47 ( .A(n158), .Y(n218) );
  INVX2 U48 ( .A(n163), .Y(n217) );
  INVX1 U49 ( .A(n145), .Y(n223) );
  INVX1 U50 ( .A(n215), .Y(n220) );
  AND2X1 U51 ( .A(n148), .B(n45), .Y(n38) );
  INVX1 U52 ( .A(n40), .Y(n39) );
  INVX1 U53 ( .A(\writedata<7> ), .Y(n40) );
  INVX1 U54 ( .A(n180), .Y(n41) );
  AND2X2 U55 ( .A(\writedata<2> ), .B(n162), .Y(n42) );
  INVX1 U56 ( .A(\writedata<6> ), .Y(n43) );
  AND2X2 U57 ( .A(n51), .B(n45), .Y(n44) );
  INVX1 U58 ( .A(n204), .Y(n46) );
  BUFX2 U59 ( .A(\writedata<2> ), .Y(n47) );
  INVX1 U60 ( .A(\writedata<4> ), .Y(n48) );
  INVX1 U61 ( .A(n48), .Y(n49) );
  INVX1 U62 ( .A(\writedata<3> ), .Y(n50) );
  INVX1 U63 ( .A(n50), .Y(n51) );
  INVX1 U64 ( .A(n187), .Y(n52) );
  INVX1 U65 ( .A(n194), .Y(n53) );
  AND2X2 U66 ( .A(n175), .B(n51), .Y(n54) );
  INVX4 U67 ( .A(n175), .Y(n174) );
  OR2X2 U68 ( .A(n181), .B(n164), .Y(n55) );
  INVX1 U69 ( .A(n55), .Y(n56) );
  OR2X2 U70 ( .A(n204), .B(n178), .Y(n57) );
  INVX1 U71 ( .A(n57), .Y(n58) );
  OR2X2 U72 ( .A(n40), .B(n177), .Y(n59) );
  INVX1 U73 ( .A(n59), .Y(n60) );
  OR2X2 U74 ( .A(n43), .B(n174), .Y(n61) );
  INVX1 U75 ( .A(n61), .Y(n62) );
  OR2X2 U76 ( .A(n182), .B(n178), .Y(n63) );
  INVX1 U77 ( .A(n63), .Y(n64) );
  OR2X2 U78 ( .A(n183), .B(n177), .Y(n65) );
  INVX1 U79 ( .A(n65), .Y(n66) );
  OR2X2 U80 ( .A(n184), .B(n178), .Y(n67) );
  INVX1 U81 ( .A(n67), .Y(n68) );
  OR2X2 U82 ( .A(n185), .B(n177), .Y(n69) );
  INVX1 U83 ( .A(n69), .Y(n70) );
  OR2X2 U84 ( .A(n183), .B(n174), .Y(n71) );
  INVX1 U85 ( .A(n71), .Y(n72) );
  OR2X2 U86 ( .A(n184), .B(n174), .Y(n73) );
  INVX1 U87 ( .A(n73), .Y(n74) );
  OR2X2 U88 ( .A(n186), .B(n174), .Y(n75) );
  INVX1 U89 ( .A(n75), .Y(n76) );
  OR2X2 U90 ( .A(n188), .B(n137), .Y(n77) );
  INVX1 U91 ( .A(n77), .Y(n78) );
  OR2X2 U92 ( .A(n189), .B(n167), .Y(n79) );
  INVX1 U93 ( .A(n79), .Y(n80) );
  OR2X2 U94 ( .A(n190), .B(n167), .Y(n81) );
  INVX1 U95 ( .A(n81), .Y(n82) );
  OR2X2 U96 ( .A(n188), .B(n167), .Y(n83) );
  INVX1 U97 ( .A(n83), .Y(n84) );
  OR2X2 U98 ( .A(n191), .B(n171), .Y(n85) );
  INVX1 U99 ( .A(n85), .Y(n86) );
  OR2X2 U100 ( .A(n192), .B(n171), .Y(n87) );
  INVX1 U101 ( .A(n87), .Y(n88) );
  OR2X2 U102 ( .A(n193), .B(n159), .Y(n89) );
  INVX1 U103 ( .A(n89), .Y(n90) );
  OR2X2 U104 ( .A(n194), .B(n171), .Y(n91) );
  INVX1 U105 ( .A(n91), .Y(n92) );
  OR2X2 U106 ( .A(n192), .B(n164), .Y(n93) );
  INVX1 U107 ( .A(n93), .Y(n94) );
  OR2X2 U108 ( .A(n195), .B(n159), .Y(n95) );
  INVX1 U109 ( .A(n95), .Y(n96) );
  OR2X2 U110 ( .A(n196), .B(n156), .Y(n97) );
  INVX1 U111 ( .A(n97), .Y(n98) );
  OR2X2 U112 ( .A(n164), .B(n198), .Y(n99) );
  INVX1 U113 ( .A(n99), .Y(n100) );
  OR2X2 U114 ( .A(n199), .B(n164), .Y(n101) );
  INVX1 U115 ( .A(n101), .Y(n102) );
  OR2X2 U116 ( .A(n159), .B(n198), .Y(n103) );
  INVX1 U117 ( .A(n103), .Y(n104) );
  OR2X2 U118 ( .A(n201), .B(n159), .Y(n105) );
  INVX1 U119 ( .A(n105), .Y(n106) );
  OR2X2 U120 ( .A(n156), .B(n202), .Y(n107) );
  INVX1 U121 ( .A(n107), .Y(n108) );
  OR2X2 U122 ( .A(n201), .B(n156), .Y(n109) );
  INVX1 U123 ( .A(n109), .Y(n110) );
  OR2X2 U124 ( .A(n174), .B(n200), .Y(n111) );
  INVX1 U125 ( .A(n111), .Y(n112) );
  OR2X2 U126 ( .A(n197), .B(n174), .Y(n113) );
  INVX1 U127 ( .A(n113), .Y(n114) );
  OR2X2 U128 ( .A(n167), .B(n203), .Y(n115) );
  INVX1 U129 ( .A(n115), .Y(n116) );
  OR2X2 U130 ( .A(n33), .B(n167), .Y(n117) );
  INVX1 U131 ( .A(n117), .Y(n118) );
  OR2X2 U132 ( .A(n137), .B(n202), .Y(n119) );
  INVX1 U133 ( .A(n119), .Y(n120) );
  OR2X2 U134 ( .A(n199), .B(n137), .Y(n121) );
  INVX1 U135 ( .A(n121), .Y(n122) );
  OR2X2 U136 ( .A(n171), .B(n203), .Y(n123) );
  INVX1 U137 ( .A(n123), .Y(n124) );
  OR2X2 U138 ( .A(n197), .B(n171), .Y(n125) );
  INVX1 U139 ( .A(n125), .Y(n126) );
  OR2X2 U140 ( .A(n178), .B(n200), .Y(n127) );
  INVX1 U141 ( .A(n127), .Y(n128) );
  OR2X2 U142 ( .A(n33), .B(n177), .Y(n129) );
  INVX1 U143 ( .A(n129), .Y(n130) );
  OR2X2 U144 ( .A(n157), .B(n133), .Y(n131) );
  INVX1 U145 ( .A(n131), .Y(n132) );
  OR2X2 U146 ( .A(n145), .B(n215), .Y(n133) );
  OR2X2 U147 ( .A(n161), .B(n136), .Y(n134) );
  INVX1 U148 ( .A(n134), .Y(n135) );
  OR2X2 U149 ( .A(n160), .B(n215), .Y(n136) );
  OR2X2 U150 ( .A(n161), .B(n138), .Y(n137) );
  OR2X2 U151 ( .A(n168), .B(n169), .Y(n138) );
  OR2X2 U152 ( .A(n173), .B(n141), .Y(n139) );
  INVX1 U153 ( .A(n139), .Y(n140) );
  OR2X2 U154 ( .A(n145), .B(n172), .Y(n141) );
  OR2X2 U155 ( .A(n180), .B(n174), .Y(n142) );
  INVX1 U156 ( .A(n142), .Y(n143) );
  BUFX2 U157 ( .A(\writeregsel<2> ), .Y(n144) );
  BUFX2 U158 ( .A(\writeregsel<0> ), .Y(n145) );
  BUFX2 U159 ( .A(\writeregsel<1> ), .Y(n146) );
  AND2X2 U160 ( .A(write), .B(n144), .Y(n147) );
  INVX1 U161 ( .A(n204), .Y(n148) );
  INVX1 U162 ( .A(\writedata<4> ), .Y(n149) );
  INVX1 U163 ( .A(n149), .Y(n150) );
  INVX1 U164 ( .A(n205), .Y(n151) );
  AND2X1 U165 ( .A(\writedata<15> ), .B(n175), .Y(\r3in<15> ) );
  INVX1 U166 ( .A(\writedata<12> ), .Y(n152) );
  INVX1 U167 ( .A(n152), .Y(n153) );
  AND2X2 U168 ( .A(n146), .B(n145), .Y(n154) );
  AND2X1 U169 ( .A(n154), .B(n147), .Y(n179) );
  INVX1 U170 ( .A(n132), .Y(n155) );
  INVX1 U171 ( .A(n132), .Y(n156) );
  INVX1 U172 ( .A(n146), .Y(n157) );
  INVX1 U173 ( .A(n135), .Y(n158) );
  INVX1 U174 ( .A(n135), .Y(n159) );
  INVX1 U175 ( .A(n173), .Y(n160) );
  INVX1 U176 ( .A(n145), .Y(n161) );
  INVX1 U177 ( .A(n216), .Y(n162) );
  INVX1 U178 ( .A(n162), .Y(n163) );
  INVX1 U179 ( .A(n162), .Y(n164) );
  INVX1 U180 ( .A(n221), .Y(n165) );
  INVX1 U181 ( .A(n165), .Y(n166) );
  INVX1 U182 ( .A(n165), .Y(n167) );
  INVX1 U183 ( .A(n157), .Y(n168) );
  INVX1 U184 ( .A(n147), .Y(n169) );
  INVX1 U185 ( .A(n140), .Y(n170) );
  INVX1 U186 ( .A(n140), .Y(n171) );
  INVX1 U187 ( .A(n147), .Y(n172) );
  INVX1 U188 ( .A(n146), .Y(n173) );
  AND2X2 U189 ( .A(n220), .B(n154), .Y(n175) );
  INVX1 U190 ( .A(n179), .Y(n176) );
  INVX1 U191 ( .A(n179), .Y(n177) );
  INVX1 U192 ( .A(n179), .Y(n178) );
  INVX1 U193 ( .A(\writedata<10> ), .Y(n180) );
  INVX1 U194 ( .A(\writedata<3> ), .Y(n181) );
  INVX1 U195 ( .A(\writedata<3> ), .Y(n182) );
  INVX1 U196 ( .A(\writedata<1> ), .Y(n183) );
  INVX1 U197 ( .A(\writedata<0> ), .Y(n184) );
  INVX1 U198 ( .A(\writedata<2> ), .Y(n185) );
  INVX1 U199 ( .A(\writedata<2> ), .Y(n186) );
  INVX1 U200 ( .A(\writedata<1> ), .Y(n187) );
  INVX1 U201 ( .A(\writedata<0> ), .Y(n188) );
  INVX1 U202 ( .A(\writedata<3> ), .Y(n189) );
  INVX1 U203 ( .A(\writedata<1> ), .Y(n190) );
  INVX1 U204 ( .A(\writedata<3> ), .Y(n191) );
  INVX1 U205 ( .A(\writedata<1> ), .Y(n192) );
  INVX1 U206 ( .A(\writedata<3> ), .Y(n193) );
  INVX1 U207 ( .A(\writedata<0> ), .Y(n194) );
  INVX1 U208 ( .A(\writedata<2> ), .Y(n195) );
  INVX1 U209 ( .A(\writedata<3> ), .Y(n196) );
  INVX1 U210 ( .A(\writedata<9> ), .Y(n197) );
  INVX1 U211 ( .A(\writedata<11> ), .Y(n198) );
  INVX1 U212 ( .A(\writedata<9> ), .Y(n199) );
  INVX1 U213 ( .A(\writedata<11> ), .Y(n200) );
  INVX1 U214 ( .A(\writedata<9> ), .Y(n201) );
  INVX1 U215 ( .A(\writedata<11> ), .Y(n202) );
  INVX1 U216 ( .A(\writedata<11> ), .Y(n203) );
  AND2X2 U217 ( .A(\writedata<8> ), .B(n225), .Y(\r7in<8> ) );
  INVX1 U218 ( .A(\writedata<6> ), .Y(n204) );
  INVX1 U219 ( .A(\writedata<4> ), .Y(n205) );
  INVX1 U220 ( .A(n207), .Y(n206) );
  AND2X2 U221 ( .A(\writedata<12> ), .B(n225), .Y(\r7in<12> ) );
  INVX1 U222 ( .A(\writedata<12> ), .Y(n207) );
  INVX1 U223 ( .A(n207), .Y(n208) );
  INVX1 U224 ( .A(\writedata<7> ), .Y(n209) );
  INVX1 U225 ( .A(n209), .Y(n210) );
  INVX1 U226 ( .A(n204), .Y(n211) );
  OR2X2 U227 ( .A(n144), .B(n214), .Y(n215) );
  NAND3X1 U228 ( .A(n223), .B(n220), .C(n157), .Y(n216) );
  AND2X2 U229 ( .A(\writedata<15> ), .B(n217), .Y(\r0in<15> ) );
  AND2X2 U230 ( .A(\writedata<14> ), .B(n217), .Y(\r0in<14> ) );
  AND2X2 U231 ( .A(\writedata<13> ), .B(n217), .Y(\r0in<13> ) );
  AND2X2 U232 ( .A(n153), .B(n217), .Y(\r0in<12> ) );
  AND2X2 U233 ( .A(n35), .B(n217), .Y(\r0in<10> ) );
  AND2X2 U234 ( .A(\writedata<8> ), .B(n217), .Y(\r0in<8> ) );
  AND2X2 U235 ( .A(n39), .B(n217), .Y(\r0in<7> ) );
  AND2X2 U236 ( .A(n148), .B(n217), .Y(\r0in<6> ) );
  AND2X2 U237 ( .A(\writedata<5> ), .B(n217), .Y(\r0in<5> ) );
  AND2X2 U238 ( .A(n49), .B(n217), .Y(\r0in<4> ) );
  AND2X2 U239 ( .A(n53), .B(n217), .Y(\r0in<0> ) );
  AND2X2 U240 ( .A(\writedata<15> ), .B(n218), .Y(\r1in<15> ) );
  AND2X2 U241 ( .A(\writedata<14> ), .B(n218), .Y(\r1in<14> ) );
  AND2X2 U242 ( .A(\writedata<13> ), .B(n218), .Y(\r1in<13> ) );
  AND2X2 U243 ( .A(n153), .B(n218), .Y(\r1in<12> ) );
  AND2X2 U244 ( .A(\writedata<10> ), .B(n218), .Y(\r1in<10> ) );
  AND2X2 U245 ( .A(\writedata<8> ), .B(n218), .Y(\r1in<8> ) );
  AND2X2 U246 ( .A(n36), .B(n218), .Y(\r1in<7> ) );
  AND2X2 U247 ( .A(n46), .B(n218), .Y(\r1in<6> ) );
  AND2X2 U248 ( .A(\writedata<5> ), .B(n218), .Y(\r1in<5> ) );
  AND2X2 U249 ( .A(n150), .B(n218), .Y(\r1in<4> ) );
  AND2X2 U250 ( .A(n52), .B(n218), .Y(\r1in<1> ) );
  AND2X2 U251 ( .A(n53), .B(n218), .Y(\r1in<0> ) );
  AND2X2 U252 ( .A(\writedata<15> ), .B(n219), .Y(\r2in<15> ) );
  AND2X2 U253 ( .A(\writedata<14> ), .B(n219), .Y(\r2in<14> ) );
  AND2X2 U254 ( .A(\writedata<13> ), .B(n219), .Y(\r2in<13> ) );
  AND2X2 U255 ( .A(n206), .B(n219), .Y(\r2in<12> ) );
  AND2X2 U256 ( .A(n35), .B(n219), .Y(\r2in<10> ) );
  AND2X2 U257 ( .A(\writedata<8> ), .B(n219), .Y(\r2in<8> ) );
  AND2X2 U258 ( .A(n39), .B(n219), .Y(\r2in<7> ) );
  AND2X2 U259 ( .A(n211), .B(n219), .Y(\r2in<6> ) );
  AND2X2 U260 ( .A(\writedata<5> ), .B(n219), .Y(\r2in<5> ) );
  AND2X2 U261 ( .A(n150), .B(n219), .Y(\r2in<4> ) );
  AND2X2 U262 ( .A(n47), .B(n219), .Y(\r2in<2> ) );
  AND2X2 U263 ( .A(n52), .B(n219), .Y(\r2in<1> ) );
  AND2X2 U264 ( .A(n53), .B(n219), .Y(\r2in<0> ) );
  AND2X2 U265 ( .A(\writedata<14> ), .B(n175), .Y(\r3in<14> ) );
  AND2X2 U266 ( .A(\writedata<13> ), .B(n175), .Y(\r3in<13> ) );
  AND2X2 U267 ( .A(n206), .B(n175), .Y(\r3in<12> ) );
  AND2X2 U268 ( .A(\writedata<8> ), .B(n175), .Y(\r3in<8> ) );
  AND2X2 U269 ( .A(n210), .B(n175), .Y(\r3in<7> ) );
  AND2X2 U270 ( .A(\writedata<5> ), .B(n175), .Y(\r3in<5> ) );
  AND2X2 U271 ( .A(n150), .B(n175), .Y(\r3in<4> ) );
  NAND3X1 U272 ( .A(n223), .B(n147), .C(n173), .Y(n221) );
  AND2X2 U273 ( .A(\writedata<15> ), .B(n222), .Y(\r4in<15> ) );
  AND2X2 U274 ( .A(\writedata<14> ), .B(n222), .Y(\r4in<14> ) );
  AND2X2 U275 ( .A(\writedata<13> ), .B(n222), .Y(\r4in<13> ) );
  AND2X2 U276 ( .A(n208), .B(n222), .Y(\r4in<12> ) );
  AND2X2 U277 ( .A(\writedata<10> ), .B(n222), .Y(\r4in<10> ) );
  AND2X2 U278 ( .A(\writedata<8> ), .B(n222), .Y(\r4in<8> ) );
  AND2X2 U279 ( .A(n210), .B(n222), .Y(\r4in<7> ) );
  AND2X2 U280 ( .A(n211), .B(n222), .Y(\r4in<6> ) );
  AND2X2 U281 ( .A(\writedata<5> ), .B(n222), .Y(\r4in<5> ) );
  AND2X2 U282 ( .A(n151), .B(n222), .Y(\r4in<4> ) );
  AND2X2 U283 ( .A(n47), .B(n222), .Y(\r4in<2> ) );
  AND2X2 U284 ( .A(\writedata<15> ), .B(n45), .Y(\r5in<15> ) );
  AND2X2 U285 ( .A(\writedata<14> ), .B(n45), .Y(\r5in<14> ) );
  AND2X2 U286 ( .A(\writedata<13> ), .B(n45), .Y(\r5in<13> ) );
  AND2X2 U287 ( .A(n208), .B(n45), .Y(\r5in<12> ) );
  AND2X2 U288 ( .A(n35), .B(n45), .Y(\r5in<10> ) );
  AND2X2 U289 ( .A(\writedata<8> ), .B(n45), .Y(\r5in<8> ) );
  AND2X2 U290 ( .A(n36), .B(n45), .Y(\r5in<7> ) );
  AND2X2 U291 ( .A(\writedata<5> ), .B(n45), .Y(\r5in<5> ) );
  AND2X2 U292 ( .A(n151), .B(n45), .Y(\r5in<4> ) );
  AND2X2 U293 ( .A(n47), .B(n45), .Y(\r5in<2> ) );
  AND2X2 U294 ( .A(\writedata<15> ), .B(n224), .Y(\r6in<15> ) );
  AND2X2 U295 ( .A(\writedata<14> ), .B(n224), .Y(\r6in<14> ) );
  AND2X2 U296 ( .A(\writedata<13> ), .B(n224), .Y(\r6in<13> ) );
  AND2X2 U297 ( .A(n208), .B(n224), .Y(\r6in<12> ) );
  AND2X2 U298 ( .A(n41), .B(n224), .Y(\r6in<10> ) );
  AND2X2 U299 ( .A(\writedata<8> ), .B(n224), .Y(\r6in<8> ) );
  AND2X2 U300 ( .A(n39), .B(n224), .Y(\r6in<7> ) );
  AND2X2 U301 ( .A(n46), .B(n224), .Y(\r6in<6> ) );
  AND2X2 U302 ( .A(\writedata<5> ), .B(n224), .Y(\r6in<5> ) );
  AND2X2 U303 ( .A(n49), .B(n224), .Y(\r6in<4> ) );
  AND2X2 U304 ( .A(n47), .B(n224), .Y(\r6in<2> ) );
  AND2X2 U305 ( .A(\writedata<15> ), .B(n225), .Y(\r7in<15> ) );
  AND2X2 U306 ( .A(\writedata<14> ), .B(n225), .Y(\r7in<14> ) );
  AND2X2 U307 ( .A(\writedata<13> ), .B(n225), .Y(\r7in<13> ) );
  AND2X2 U308 ( .A(n41), .B(n225), .Y(\r7in<10> ) );
  AND2X2 U309 ( .A(\writedata<5> ), .B(n225), .Y(\r7in<5> ) );
  AND2X2 U310 ( .A(n151), .B(n225), .Y(\r7in<4> ) );
endmodule


module alu ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , 
        \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> 
        }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , 
        \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> 
        }), Cin, .Op({\Op<3> , \Op<2> , \Op<1> , \Op<0> }), passthrough, 
        reverse, invA, invB, sign, .Out({\Out<15> , \Out<14> , \Out<13> , 
        \Out<12> , \Out<11> , \Out<10> , \Out<9> , \Out<8> , \Out<7> , 
        \Out<6> , \Out<5> , \Out<4> , \Out<3> , \Out<2> , \Out<1> , \Out<0> }), 
        Ofl, zero );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin,
         \Op<3> , \Op<2> , \Op<1> , \Op<0> , passthrough, reverse, invA, invB,
         sign;
  output \Out<15> , \Out<14> , \Out<13> , \Out<12> , \Out<11> , \Out<10> ,
         \Out<9> , \Out<8> , \Out<7> , \Out<6> , \Out<5> , \Out<4> , \Out<3> ,
         \Out<2> , \Out<1> , \Out<0> , Ofl, zero;
  wire   \A_inv<0> , overflow, Cout, \shift_out<15> , \shift_out<14> ,
         \shift_out<13> , \shift_out<12> , \shift_out<11> , \shift_out<10> ,
         \shift_out<9> , \shift_out<8> , \shift_out<7> , \shift_out<6> ,
         \shift_out<5> , \shift_out<4> , \shift_out<3> , \shift_out<2> ,
         \shift_out<1> , \shift_out<0> , \sum<15> , \sum<14> , \sum<13> ,
         \sum<12> , \sum<11> , \sum<10> , \sum<9> , \sum<8> , \sum<7> ,
         \sum<6> , \sum<5> , \sum<4> , \sum<3> , \sum<2> , \sum<1> , \sum<0> ,
         n231, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44,
         n45, n46, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n191, n192, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n378, n379, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621;

  AOI22X1 U214 ( .A(n396), .B(n621), .C(sign), .D(overflow), .Y(n231) );
  shifter shift ( .In({n13, n620, n619, n618, n617, n400, n616, n215, n349, 
        n604, n381, n602, n209, n355, n399, \A_inv<0> }), .Cnt({n609, n608, 
        n598, n607}), .Op({\Op<2> , \Op<1> , \Op<0> }), .Out({\shift_out<15> , 
        \shift_out<14> , \shift_out<13> , \shift_out<12> , \shift_out<11> , 
        \shift_out<10> , \shift_out<9> , \shift_out<8> , \shift_out<7> , 
        \shift_out<6> , \shift_out<5> , \shift_out<4> , \shift_out<3> , 
        \shift_out<2> , \shift_out<1> , \shift_out<0> }) );
  adder_0 add ( .A({n606, n620, n619, n618, n617, n400, n369, n215, n605, n604, 
        n603, n244, n601, n355, n399, n366}), .B({n387, n615, n16, n6, n36, 
        n38, n614, n242, n613, n612, n611, n610, n609, n608, n34, n393}), 
        .Cin(Cin), .Overflow(overflow), .Cout(Cout), .Sum({\sum<15> , 
        \sum<14> , \sum<13> , \sum<12> , \sum<11> , \sum<10> , \sum<9> , 
        \sum<8> , \sum<7> , \sum<6> , \sum<5> , \sum<4> , \sum<3> , \sum<2> , 
        \sum<1> , \sum<0> }) );
  INVX4 U2 ( .A(n413), .Y(n355) );
  INVX1 U3 ( .A(n405), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  BUFX2 U5 ( .A(n415), .Y(n3) );
  INVX1 U6 ( .A(\Out<6> ), .Y(n4) );
  INVX1 U7 ( .A(n4), .Y(n5) );
  INVX4 U8 ( .A(n453), .Y(n604) );
  INVX4 U9 ( .A(n414), .Y(n399) );
  INVX2 U10 ( .A(n210), .Y(n601) );
  INVX2 U11 ( .A(n367), .Y(n358) );
  INVX2 U12 ( .A(invB), .Y(n367) );
  INVX4 U13 ( .A(n403), .Y(n379) );
  XOR2X1 U14 ( .A(\B<12> ), .B(n358), .Y(n6) );
  INVX2 U15 ( .A(\B<4> ), .Y(n526) );
  INVX4 U16 ( .A(n168), .Y(\Out<1> ) );
  INVX4 U17 ( .A(n419), .Y(n611) );
  BUFX2 U18 ( .A(\Op<0> ), .Y(n7) );
  AND2X2 U19 ( .A(n94), .B(n270), .Y(n138) );
  INVX1 U20 ( .A(\A<14> ), .Y(n553) );
  INVX1 U21 ( .A(\A<12> ), .Y(n547) );
  INVX1 U22 ( .A(\A<0> ), .Y(n522) );
  AND2X1 U23 ( .A(n250), .B(n248), .Y(n306) );
  INVX1 U24 ( .A(\A<4> ), .Y(n520) );
  INVX1 U25 ( .A(\A<15> ), .Y(n516) );
  AND2X1 U26 ( .A(n299), .B(n321), .Y(n44) );
  INVX1 U27 ( .A(\A<10> ), .Y(n541) );
  INVX1 U28 ( .A(\A<11> ), .Y(n543) );
  INVX1 U29 ( .A(\A<1> ), .Y(n523) );
  INVX1 U30 ( .A(n474), .Y(n475) );
  INVX1 U31 ( .A(\A<2> ), .Y(n521) );
  INVX1 U32 ( .A(\A<15> ), .Y(n14) );
  AND2X1 U33 ( .A(n571), .B(n570), .Y(n187) );
  INVX1 U34 ( .A(\A<3> ), .Y(n525) );
  INVX1 U35 ( .A(\A<6> ), .Y(n531) );
  INVX1 U36 ( .A(\A<7> ), .Y(n533) );
  INVX1 U37 ( .A(n556), .Y(n20) );
  INVX1 U38 ( .A(n411), .Y(n603) );
  INVX1 U39 ( .A(n574), .Y(n445) );
  AND2X1 U40 ( .A(\sum<1> ), .B(n592), .Y(n55) );
  AND2X1 U41 ( .A(n390), .B(n246), .Y(n389) );
  INVX1 U42 ( .A(\A<5> ), .Y(n519) );
  INVX1 U43 ( .A(n578), .Y(n454) );
  INVX1 U44 ( .A(sign), .Y(n621) );
  INVX1 U45 ( .A(n555), .Y(n581) );
  AND2X1 U46 ( .A(n314), .B(n293), .Y(n220) );
  INVX2 U47 ( .A(n22), .Y(\Out<12> ) );
  INVX1 U48 ( .A(n452), .Y(n10) );
  BUFX2 U49 ( .A(\B<13> ), .Y(n8) );
  AND2X2 U50 ( .A(n21), .B(n10), .Y(n9) );
  INVX8 U51 ( .A(n9), .Y(\Out<5> ) );
  NOR3X1 U52 ( .A(\Out<5> ), .B(\Out<1> ), .C(n5), .Y(n11) );
  AND2X1 U53 ( .A(\sum<7> ), .B(n592), .Y(n207) );
  NOR3X1 U54 ( .A(n200), .B(n374), .C(n45), .Y(n12) );
  XNOR2X1 U55 ( .A(n405), .B(n14), .Y(n13) );
  BUFX4 U56 ( .A(\B<5> ), .Y(n15) );
  XNOR2X1 U57 ( .A(n372), .B(n379), .Y(n509) );
  XOR2X1 U58 ( .A(\B<13> ), .B(n233), .Y(n16) );
  BUFX2 U59 ( .A(n6), .Y(n17) );
  BUFX2 U60 ( .A(\B<12> ), .Y(n18) );
  NOR3X1 U61 ( .A(n294), .B(n177), .C(n20), .Y(n19) );
  INVX2 U62 ( .A(n19), .Y(n582) );
  NOR3X1 U63 ( .A(n287), .B(n310), .C(n181), .Y(n21) );
  NOR3X1 U64 ( .A(n289), .B(n178), .C(n23), .Y(n22) );
  INVX1 U65 ( .A(n462), .Y(n23) );
  NOR3X1 U66 ( .A(n25), .B(n311), .C(n319), .Y(n24) );
  INVX2 U67 ( .A(n24), .Y(\Out<6> ) );
  INVX1 U68 ( .A(n458), .Y(n25) );
  NOR3X1 U69 ( .A(n27), .B(n332), .C(n335), .Y(n26) );
  INVX1 U70 ( .A(n26), .Y(\Out<8> ) );
  INVX1 U71 ( .A(n471), .Y(n27) );
  BUFX2 U72 ( .A(\Out<8> ), .Y(n28) );
  BUFX2 U73 ( .A(\B<10> ), .Y(n29) );
  BUFX2 U74 ( .A(n2), .Y(n30) );
  BUFX2 U75 ( .A(\B<1> ), .Y(n385) );
  BUFX2 U76 ( .A(invA), .Y(n404) );
  BUFX2 U77 ( .A(invA), .Y(n405) );
  INVX1 U78 ( .A(n57), .Y(\Out<2> ) );
  NOR3X1 U79 ( .A(n291), .B(n312), .C(n182), .Y(n31) );
  INVX1 U80 ( .A(n31), .Y(n483) );
  INVX8 U81 ( .A(n217), .Y(\Out<4> ) );
  INVX2 U82 ( .A(n216), .Y(n217) );
  BUFX2 U83 ( .A(invB), .Y(n403) );
  AND2X2 U84 ( .A(n124), .B(n116), .Y(n33) );
  INVX1 U85 ( .A(n33), .Y(n34) );
  AND2X2 U86 ( .A(n128), .B(n118), .Y(n35) );
  INVX1 U87 ( .A(n35), .Y(n36) );
  AND2X2 U88 ( .A(n130), .B(n120), .Y(n37) );
  INVX1 U89 ( .A(n37), .Y(n38) );
  INVX1 U90 ( .A(n143), .Y(\Out<7> ) );
  AND2X2 U91 ( .A(n213), .B(n297), .Y(n40) );
  AND2X2 U92 ( .A(n40), .B(n214), .Y(n41) );
  INVX1 U93 ( .A(n41), .Y(n42) );
  OR2X2 U94 ( .A(n64), .B(n62), .Y(n43) );
  INVX1 U95 ( .A(n147), .Y(n45) );
  AND2X2 U96 ( .A(\A<3> ), .B(n2), .Y(n46) );
  INVX1 U97 ( .A(n46), .Y(n47) );
  OR2X2 U98 ( .A(n394), .B(n395), .Y(\Out<14> ) );
  OR2X2 U99 ( .A(n132), .B(n569), .Y(n49) );
  AND2X2 U100 ( .A(n276), .B(n114), .Y(n50) );
  AND2X2 U101 ( .A(n435), .B(n222), .Y(n51) );
  AND2X2 U102 ( .A(n232), .B(n429), .Y(n52) );
  AND2X2 U103 ( .A(n435), .B(n581), .Y(n53) );
  AND2X2 U104 ( .A(n329), .B(n345), .Y(n54) );
  INVX1 U105 ( .A(n55), .Y(n56) );
  AND2X2 U106 ( .A(n266), .B(n122), .Y(n57) );
  INVX1 U107 ( .A(n57), .Y(n58) );
  OR2X2 U108 ( .A(n340), .B(n497), .Y(n59) );
  INVX1 U109 ( .A(n59), .Y(n60) );
  OR2X2 U110 ( .A(n521), .B(\B<2> ), .Y(n61) );
  INVX1 U111 ( .A(n61), .Y(n62) );
  OR2X2 U112 ( .A(n523), .B(n352), .Y(n63) );
  INVX1 U113 ( .A(n63), .Y(n64) );
  OR2X2 U114 ( .A(n541), .B(n29), .Y(n65) );
  INVX1 U115 ( .A(n65), .Y(n66) );
  AND2X2 U116 ( .A(n18), .B(n547), .Y(n67) );
  INVX1 U117 ( .A(n67), .Y(n68) );
  AND2X2 U118 ( .A(n126), .B(n580), .Y(n69) );
  INVX1 U119 ( .A(n69), .Y(n70) );
  BUFX2 U120 ( .A(n456), .Y(n71) );
  BUFX2 U121 ( .A(n505), .Y(n72) );
  AND2X2 U122 ( .A(\A<8> ), .B(n2), .Y(n73) );
  INVX1 U123 ( .A(n73), .Y(n74) );
  AND2X2 U124 ( .A(\shift_out<9> ), .B(n401), .Y(n75) );
  INVX1 U125 ( .A(n75), .Y(n76) );
  BUFX2 U126 ( .A(n515), .Y(n77) );
  BUFX2 U127 ( .A(n444), .Y(n78) );
  BUFX2 U128 ( .A(n485), .Y(n79) );
  BUFX2 U129 ( .A(n493), .Y(n80) );
  BUFX2 U130 ( .A(n585), .Y(n81) );
  BUFX2 U131 ( .A(n594), .Y(n82) );
  AND2X2 U132 ( .A(n236), .B(n237), .Y(n83) );
  INVX1 U133 ( .A(n83), .Y(n84) );
  AND2X2 U134 ( .A(n528), .B(n225), .Y(n85) );
  INVX1 U135 ( .A(n85), .Y(n86) );
  AND2X2 U136 ( .A(n386), .B(n237), .Y(n87) );
  INVX1 U137 ( .A(n87), .Y(n88) );
  AND2X2 U138 ( .A(n592), .B(\sum<15> ), .Y(n89) );
  INVX1 U139 ( .A(n89), .Y(n90) );
  AND2X2 U140 ( .A(n241), .B(n341), .Y(n91) );
  INVX1 U141 ( .A(n91), .Y(n92) );
  AND2X2 U142 ( .A(n401), .B(\shift_out<13> ), .Y(n93) );
  INVX1 U143 ( .A(n93), .Y(n94) );
  AND2X2 U144 ( .A(\shift_out<3> ), .B(n401), .Y(n95) );
  INVX1 U145 ( .A(n95), .Y(n96) );
  AND2X2 U146 ( .A(\sum<10> ), .B(n592), .Y(n97) );
  INVX1 U147 ( .A(n97), .Y(n98) );
  OR2X2 U148 ( .A(n567), .B(n149), .Y(n99) );
  INVX1 U149 ( .A(n99), .Y(n100) );
  BUFX2 U150 ( .A(n433), .Y(n101) );
  BUFX2 U151 ( .A(n441), .Y(n102) );
  BUFX2 U152 ( .A(n464), .Y(n103) );
  BUFX2 U153 ( .A(n476), .Y(n104) );
  BUFX2 U154 ( .A(n486), .Y(n105) );
  BUFX2 U155 ( .A(n494), .Y(n106) );
  BUFX2 U156 ( .A(n503), .Y(n107) );
  BUFX2 U157 ( .A(n511), .Y(n108) );
  BUFX2 U158 ( .A(n587), .Y(n109) );
  AND2X2 U159 ( .A(\sum<12> ), .B(n592), .Y(n110) );
  INVX1 U160 ( .A(n110), .Y(n111) );
  AND2X2 U161 ( .A(n532), .B(\A<8> ), .Y(n112) );
  INVX1 U162 ( .A(n112), .Y(n113) );
  BUFX2 U163 ( .A(n514), .Y(n114) );
  AND2X2 U164 ( .A(n238), .B(n239), .Y(n115) );
  INVX1 U165 ( .A(n115), .Y(n116) );
  AND2X2 U166 ( .A(n370), .B(n403), .Y(n117) );
  INVX1 U167 ( .A(n117), .Y(n118) );
  AND2X2 U168 ( .A(n378), .B(n234), .Y(n119) );
  INVX1 U169 ( .A(n119), .Y(n120) );
  AND2X2 U170 ( .A(\shift_out<2> ), .B(n401), .Y(n121) );
  INVX1 U171 ( .A(n121), .Y(n122) );
  AND2X2 U172 ( .A(n385), .B(n367), .Y(n123) );
  INVX1 U173 ( .A(n123), .Y(n124) );
  OR2X2 U174 ( .A(n49), .B(n205), .Y(n125) );
  INVX1 U175 ( .A(n125), .Y(n126) );
  AND2X2 U176 ( .A(\B<11> ), .B(n379), .Y(n127) );
  INVX1 U177 ( .A(n127), .Y(n128) );
  AND2X2 U178 ( .A(\B<10> ), .B(n379), .Y(n129) );
  INVX1 U179 ( .A(n129), .Y(n130) );
  AND2X2 U180 ( .A(n559), .B(n558), .Y(n131) );
  INVX1 U181 ( .A(n131), .Y(n132) );
  BUFX2 U182 ( .A(n524), .Y(n133) );
  AND2X2 U183 ( .A(n220), .B(n96), .Y(n134) );
  INVX1 U184 ( .A(n134), .Y(n135) );
  AND2X2 U185 ( .A(n584), .B(n81), .Y(n136) );
  INVX1 U186 ( .A(n136), .Y(n137) );
  INVX1 U187 ( .A(n138), .Y(n139) );
  AND2X2 U188 ( .A(n582), .B(n70), .Y(n140) );
  INVX1 U189 ( .A(n140), .Y(n141) );
  BUFX2 U190 ( .A(n391), .Y(\Out<9> ) );
  AND2X2 U191 ( .A(n327), .B(n208), .Y(n143) );
  INVX1 U192 ( .A(n143), .Y(n144) );
  OR2X2 U193 ( .A(Cout), .B(n141), .Y(n145) );
  INVX1 U194 ( .A(n145), .Y(n146) );
  AND2X2 U195 ( .A(n197), .B(n221), .Y(n147) );
  INVX1 U196 ( .A(n147), .Y(n148) );
  BUFX2 U197 ( .A(n566), .Y(n149) );
  AND2X2 U198 ( .A(n268), .B(n78), .Y(n150) );
  INVX1 U199 ( .A(n150), .Y(n151) );
  OR2X2 U200 ( .A(n571), .B(n402), .Y(n152) );
  INVX1 U201 ( .A(n152), .Y(n153) );
  OR2X2 U202 ( .A(n570), .B(n402), .Y(n154) );
  INVX1 U203 ( .A(n154), .Y(n155) );
  AND2X2 U204 ( .A(n272), .B(n79), .Y(n156) );
  INVX1 U205 ( .A(n156), .Y(n157) );
  OR2X2 U206 ( .A(n573), .B(n402), .Y(n158) );
  INVX1 U207 ( .A(n158), .Y(n159) );
  AND2X2 U208 ( .A(n274), .B(n80), .Y(n160) );
  INVX1 U209 ( .A(n160), .Y(n161) );
  OR2X2 U210 ( .A(n519), .B(n15), .Y(n162) );
  INVX1 U211 ( .A(n162), .Y(n163) );
  BUFX2 U212 ( .A(n398), .Y(n164) );
  BUFX2 U213 ( .A(n446), .Y(n165) );
  OR2X2 U215 ( .A(n42), .B(\Out<12> ), .Y(n166) );
  INVX1 U216 ( .A(n166), .Y(n167) );
  BUFX2 U217 ( .A(n448), .Y(n168) );
  OR2X2 U218 ( .A(n340), .B(n362), .Y(n169) );
  INVX1 U219 ( .A(n169), .Y(n170) );
  OR2X2 U220 ( .A(n340), .B(n437), .Y(n171) );
  INVX1 U221 ( .A(n171), .Y(n172) );
  AND2X2 U222 ( .A(n227), .B(n86), .Y(n173) );
  INVX1 U223 ( .A(n173), .Y(n174) );
  BUFX2 U224 ( .A(n540), .Y(n175) );
  BUFX2 U225 ( .A(n552), .Y(n176) );
  AND2X2 U226 ( .A(n554), .B(n44), .Y(n177) );
  OR2X2 U227 ( .A(n280), .B(n461), .Y(n178) );
  OR2X2 U228 ( .A(n133), .B(n43), .Y(n179) );
  INVX1 U229 ( .A(n179), .Y(n180) );
  AND2X2 U230 ( .A(n401), .B(\shift_out<5> ), .Y(n181) );
  AND2X2 U231 ( .A(\shift_out<4> ), .B(n401), .Y(n182) );
  BUFX2 U232 ( .A(n597), .Y(n183) );
  BUFX2 U233 ( .A(n579), .Y(n184) );
  AND2X2 U234 ( .A(n217), .B(n408), .Y(n185) );
  INVX1 U235 ( .A(n185), .Y(n186) );
  INVX1 U236 ( .A(n187), .Y(n188) );
  AND2X2 U237 ( .A(n265), .B(n90), .Y(n189) );
  INVX1 U238 ( .A(n189), .Y(\Out<15> ) );
  INVX1 U239 ( .A(n189), .Y(n191) );
  AND2X2 U240 ( .A(n72), .B(n98), .Y(n192) );
  INVX1 U241 ( .A(n192), .Y(\Out<10> ) );
  INVX1 U242 ( .A(n192), .Y(n194) );
  AND2X2 U243 ( .A(\sum<11> ), .B(n592), .Y(n195) );
  BUFX2 U244 ( .A(n596), .Y(n196) );
  BUFX2 U245 ( .A(n593), .Y(n197) );
  OR2X2 U246 ( .A(n137), .B(n146), .Y(n198) );
  INVX1 U247 ( .A(n198), .Y(n199) );
  INVX1 U248 ( .A(n198), .Y(n200) );
  BUFX2 U249 ( .A(n583), .Y(n201) );
  AND2X2 U250 ( .A(n50), .B(n77), .Y(n202) );
  INVX1 U251 ( .A(n202), .Y(n203) );
  AND2X2 U252 ( .A(n568), .B(n100), .Y(n204) );
  INVX1 U253 ( .A(n204), .Y(n205) );
  INVX1 U254 ( .A(n204), .Y(n206) );
  BUFX2 U255 ( .A(n588), .Y(n402) );
  INVX1 U256 ( .A(n207), .Y(n208) );
  AND2X2 U257 ( .A(n47), .B(n88), .Y(n209) );
  INVX1 U258 ( .A(n209), .Y(n210) );
  OR2X2 U259 ( .A(n139), .B(n465), .Y(n211) );
  INVX1 U260 ( .A(n211), .Y(n212) );
  INVX1 U261 ( .A(n211), .Y(n213) );
  BUFX2 U262 ( .A(n466), .Y(n214) );
  AND2X2 U263 ( .A(n74), .B(n84), .Y(n215) );
  OR2X2 U264 ( .A(n483), .B(n484), .Y(n216) );
  BUFX2 U265 ( .A(n479), .Y(n218) );
  BUFX2 U266 ( .A(reverse), .Y(n406) );
  AND2X2 U267 ( .A(n278), .B(n82), .Y(n221) );
  AND2X2 U268 ( .A(\Op<1> ), .B(n7), .Y(n222) );
  BUFX2 U269 ( .A(n527), .Y(n223) );
  INVX1 U270 ( .A(n529), .Y(n224) );
  INVX1 U271 ( .A(n224), .Y(n225) );
  INVX1 U272 ( .A(n530), .Y(n226) );
  INVX1 U273 ( .A(n226), .Y(n227) );
  INVX1 U274 ( .A(n12), .Y(n228) );
  INVX1 U275 ( .A(\Op<3> ), .Y(n229) );
  INVX1 U276 ( .A(n229), .Y(n230) );
  INVX1 U277 ( .A(n425), .Y(n232) );
  INVX1 U278 ( .A(passthrough), .Y(n425) );
  INVX1 U279 ( .A(\Op<1> ), .Y(n428) );
  INVX1 U280 ( .A(n379), .Y(n233) );
  INVX1 U281 ( .A(n367), .Y(n234) );
  BUFX2 U282 ( .A(\B<0> ), .Y(n235) );
  INVX1 U283 ( .A(\A<8> ), .Y(n236) );
  INVX1 U284 ( .A(n405), .Y(n237) );
  INVX1 U285 ( .A(n385), .Y(n238) );
  INVX1 U286 ( .A(n367), .Y(n239) );
  INVX2 U287 ( .A(n418), .Y(n613) );
  INVX1 U288 ( .A(n518), .Y(n240) );
  INVX1 U289 ( .A(n518), .Y(n241) );
  INVX2 U290 ( .A(n417), .Y(n242) );
  BUFX2 U291 ( .A(n242), .Y(n243) );
  INVX2 U292 ( .A(n412), .Y(n244) );
  INVX1 U293 ( .A(n412), .Y(n602) );
  XOR2X1 U294 ( .A(\B<8> ), .B(n379), .Y(n417) );
  AND2X2 U295 ( .A(\B<9> ), .B(n52), .Y(n245) );
  INVX1 U296 ( .A(n245), .Y(n246) );
  AND2X2 U297 ( .A(\B<2> ), .B(n521), .Y(n247) );
  INVX1 U298 ( .A(n247), .Y(n248) );
  AND2X2 U299 ( .A(\B<3> ), .B(n525), .Y(n249) );
  INVX1 U300 ( .A(n249), .Y(n250) );
  BUFX2 U301 ( .A(n550), .Y(n251) );
  BUFX2 U302 ( .A(n431), .Y(n252) );
  BUFX2 U303 ( .A(n439), .Y(n253) );
  BUFX2 U304 ( .A(n449), .Y(n254) );
  BUFX2 U305 ( .A(n480), .Y(n255) );
  BUFX2 U306 ( .A(n489), .Y(n256) );
  BUFX2 U307 ( .A(n500), .Y(n257) );
  BUFX2 U308 ( .A(n538), .Y(n258) );
  AND2X2 U309 ( .A(n407), .B(\A<7> ), .Y(n259) );
  INVX1 U310 ( .A(n259), .Y(n260) );
  AND2X2 U311 ( .A(\B<8> ), .B(n536), .Y(n261) );
  INVX1 U312 ( .A(n261), .Y(n262) );
  AND2X2 U313 ( .A(n542), .B(\A<12> ), .Y(n263) );
  INVX1 U314 ( .A(n263), .Y(n264) );
  BUFX2 U315 ( .A(n436), .Y(n265) );
  BUFX2 U316 ( .A(n488), .Y(n266) );
  AND2X2 U317 ( .A(n406), .B(\A<14> ), .Y(n267) );
  INVX1 U318 ( .A(n267), .Y(n268) );
  AND2X2 U319 ( .A(n8), .B(n52), .Y(n269) );
  INVX1 U320 ( .A(n269), .Y(n270) );
  AND2X2 U321 ( .A(n407), .B(\A<13> ), .Y(n271) );
  INVX1 U322 ( .A(n271), .Y(n272) );
  AND2X2 U323 ( .A(n407), .B(\A<8> ), .Y(n273) );
  INVX1 U324 ( .A(n273), .Y(n274) );
  AND2X2 U325 ( .A(n407), .B(\A<4> ), .Y(n275) );
  INVX1 U326 ( .A(n275), .Y(n276) );
  AND2X2 U327 ( .A(n407), .B(\A<15> ), .Y(n277) );
  INVX1 U328 ( .A(n277), .Y(n278) );
  OR2X2 U329 ( .A(n429), .B(n384), .Y(n279) );
  INVX1 U330 ( .A(n279), .Y(n280) );
  BUFX2 U331 ( .A(n231), .Y(n281) );
  BUFX2 U332 ( .A(n447), .Y(n282) );
  AND2X2 U333 ( .A(n71), .B(n92), .Y(n283) );
  INVX1 U334 ( .A(n283), .Y(n284) );
  OR2X2 U335 ( .A(n525), .B(\B<3> ), .Y(n285) );
  INVX1 U336 ( .A(n285), .Y(n286) );
  INVX1 U337 ( .A(n288), .Y(n287) );
  BUFX2 U338 ( .A(n451), .Y(n288) );
  INVX1 U339 ( .A(n290), .Y(n289) );
  BUFX2 U340 ( .A(n463), .Y(n290) );
  INVX1 U341 ( .A(n292), .Y(n291) );
  BUFX2 U342 ( .A(n482), .Y(n292) );
  BUFX2 U343 ( .A(n491), .Y(n293) );
  INVX1 U344 ( .A(n295), .Y(n294) );
  BUFX2 U345 ( .A(n557), .Y(n295) );
  AND2X2 U346 ( .A(n407), .B(\A<2> ), .Y(n296) );
  INVX1 U347 ( .A(n296), .Y(n297) );
  AND2X2 U348 ( .A(n517), .B(\A<15> ), .Y(n298) );
  INVX1 U349 ( .A(n298), .Y(n299) );
  INVX4 U350 ( .A(n437), .Y(n620) );
  BUFX2 U351 ( .A(n535), .Y(n300) );
  BUFX2 U352 ( .A(n545), .Y(n301) );
  OR2X2 U353 ( .A(n340), .B(n459), .Y(n302) );
  INVX1 U354 ( .A(n302), .Y(n303) );
  OR2X2 U355 ( .A(n340), .B(n354), .Y(n304) );
  INVX1 U356 ( .A(n304), .Y(n305) );
  INVX1 U357 ( .A(n306), .Y(n307) );
  AND2X2 U358 ( .A(n342), .B(n385), .Y(n308) );
  INVX1 U359 ( .A(n308), .Y(n309) );
  AND2X2 U360 ( .A(n15), .B(n343), .Y(n310) );
  AND2X2 U361 ( .A(n406), .B(\A<9> ), .Y(n311) );
  AND2X2 U362 ( .A(\B<4> ), .B(n342), .Y(n312) );
  AND2X2 U363 ( .A(\B<3> ), .B(n343), .Y(n313) );
  INVX1 U364 ( .A(n313), .Y(n314) );
  OR2X2 U365 ( .A(n383), .B(n195), .Y(n315) );
  INVX1 U366 ( .A(n315), .Y(n316) );
  OR2X2 U367 ( .A(n194), .B(n144), .Y(n317) );
  INVX1 U368 ( .A(n317), .Y(n318) );
  INVX1 U369 ( .A(n457), .Y(n319) );
  AND2X2 U370 ( .A(\B<14> ), .B(n553), .Y(n320) );
  INVX1 U371 ( .A(n320), .Y(n321) );
  OR2X2 U372 ( .A(n28), .B(\Out<9> ), .Y(n322) );
  INVX1 U373 ( .A(n322), .Y(n323) );
  AND2X2 U374 ( .A(n578), .B(n577), .Y(n324) );
  INVX1 U375 ( .A(n324), .Y(n325) );
  INVX1 U376 ( .A(n496), .Y(n326) );
  INVX1 U377 ( .A(n326), .Y(n327) );
  INVX1 U378 ( .A(n49), .Y(n328) );
  INVX1 U379 ( .A(n52), .Y(n329) );
  AND2X2 U380 ( .A(n375), .B(n581), .Y(n330) );
  INVX1 U381 ( .A(n330), .Y(n331) );
  INVX1 U382 ( .A(n470), .Y(n332) );
  AND2X2 U383 ( .A(n407), .B(\A<6> ), .Y(n333) );
  INVX1 U384 ( .A(n333), .Y(n334) );
  INVX1 U385 ( .A(n336), .Y(n335) );
  BUFX2 U386 ( .A(n469), .Y(n336) );
  INVX1 U387 ( .A(n53), .Y(n337) );
  INVX1 U388 ( .A(n53), .Y(n338) );
  INVX1 U389 ( .A(n51), .Y(n339) );
  INVX1 U390 ( .A(n51), .Y(n340) );
  INVX1 U391 ( .A(n54), .Y(n341) );
  INVX1 U392 ( .A(n54), .Y(n342) );
  INVX1 U393 ( .A(n54), .Y(n343) );
  INVX1 U394 ( .A(n512), .Y(n344) );
  INVX1 U395 ( .A(n344), .Y(n345) );
  INVX1 U396 ( .A(n344), .Y(n346) );
  NAND3X1 U397 ( .A(n328), .B(n347), .C(n580), .Y(n398) );
  INVX1 U398 ( .A(n206), .Y(n347) );
  XOR2X1 U399 ( .A(n397), .B(n619), .Y(n348) );
  INVX1 U400 ( .A(n348), .Y(n558) );
  INVX2 U401 ( .A(n410), .Y(n349) );
  INVX1 U402 ( .A(n410), .Y(n605) );
  INVX1 U403 ( .A(n369), .Y(n350) );
  INVX1 U404 ( .A(\B<1> ), .Y(n351) );
  INVX1 U405 ( .A(n351), .Y(n352) );
  INVX1 U406 ( .A(n617), .Y(n353) );
  INVX2 U407 ( .A(n506), .Y(n617) );
  INVX1 U408 ( .A(n215), .Y(n354) );
  INVX1 U409 ( .A(\sum<3> ), .Y(n490) );
  INVX1 U410 ( .A(\B<7> ), .Y(n356) );
  INVX1 U411 ( .A(n356), .Y(n357) );
  INVX1 U412 ( .A(n237), .Y(n359) );
  INVX1 U413 ( .A(n604), .Y(n360) );
  XNOR2X1 U414 ( .A(\B<7> ), .B(n358), .Y(n418) );
  INVX1 U415 ( .A(n13), .Y(n362) );
  XNOR2X1 U416 ( .A(n404), .B(\A<15> ), .Y(n363) );
  BUFX2 U417 ( .A(\B<2> ), .Y(n364) );
  INVX2 U418 ( .A(n422), .Y(n608) );
  BUFX2 U419 ( .A(n613), .Y(n365) );
  INVX2 U420 ( .A(n3), .Y(n366) );
  INVX1 U421 ( .A(n415), .Y(\A_inv<0> ) );
  INVX1 U422 ( .A(n367), .Y(n368) );
  INVX2 U423 ( .A(n472), .Y(n369) );
  INVX1 U424 ( .A(n472), .Y(n616) );
  INVX1 U425 ( .A(\B<11> ), .Y(n370) );
  INVX1 U426 ( .A(n237), .Y(n371) );
  INVX1 U427 ( .A(\B<11> ), .Y(n372) );
  INVX1 U428 ( .A(n372), .Y(n373) );
  BUFX2 U429 ( .A(\Out<3> ), .Y(n374) );
  INVX1 U430 ( .A(n569), .Y(n375) );
  BUFX2 U431 ( .A(n615), .Y(n376) );
  INVX1 U432 ( .A(\B<10> ), .Y(n378) );
  OR2X2 U433 ( .A(n135), .B(n492), .Y(\Out<3> ) );
  INVX1 U434 ( .A(n411), .Y(n381) );
  INVX1 U435 ( .A(n411), .Y(n382) );
  XOR2X1 U436 ( .A(\B<6> ), .B(n403), .Y(n612) );
  OR2X2 U437 ( .A(n395), .B(n394), .Y(n383) );
  INVX1 U438 ( .A(\A<3> ), .Y(n384) );
  INVX1 U439 ( .A(\A<3> ), .Y(n386) );
  INVX1 U440 ( .A(n363), .Y(n606) );
  XNOR2X1 U441 ( .A(\B<15> ), .B(n367), .Y(n387) );
  XNOR2X1 U442 ( .A(\B<15> ), .B(n379), .Y(n388) );
  INVX4 U443 ( .A(n421), .Y(n609) );
  INVX1 U444 ( .A(n201), .Y(n584) );
  AND2X2 U445 ( .A(n76), .B(n389), .Y(n478) );
  INVX1 U446 ( .A(n477), .Y(n390) );
  NAND3X1 U447 ( .A(n218), .B(n334), .C(n478), .Y(n391) );
  INVX4 U448 ( .A(n409), .Y(n619) );
  INVX1 U449 ( .A(n607), .Y(n392) );
  INVX1 U450 ( .A(n392), .Y(n393) );
  AND2X2 U451 ( .A(n592), .B(\sum<14> ), .Y(n395) );
  INVX1 U452 ( .A(n443), .Y(n394) );
  INVX1 U453 ( .A(n7), .Y(n427) );
  INVX4 U454 ( .A(n424), .Y(n598) );
  BUFX2 U455 ( .A(Cout), .Y(n396) );
  INVX1 U456 ( .A(\sum<5> ), .Y(n450) );
  BUFX2 U457 ( .A(n16), .Y(n397) );
  INVX1 U458 ( .A(n18), .Y(n542) );
  INVX1 U459 ( .A(\B<14> ), .Y(n549) );
  INVX1 U460 ( .A(\B<9> ), .Y(n537) );
  INVX1 U461 ( .A(\B<15> ), .Y(n517) );
  INVX1 U462 ( .A(n8), .Y(n548) );
  INVX1 U463 ( .A(\B<6> ), .Y(n518) );
  INVX1 U464 ( .A(n400), .Y(n497) );
  INVX1 U465 ( .A(\B<8> ), .Y(n532) );
  INVX1 U466 ( .A(n58), .Y(n408) );
  XOR2X1 U467 ( .A(n404), .B(\A<10> ), .Y(n400) );
  INVX4 U468 ( .A(n423), .Y(n607) );
  INVX1 U469 ( .A(\Op<2> ), .Y(n569) );
  OR2X2 U470 ( .A(n195), .B(n203), .Y(\Out<11> ) );
  BUFX4 U471 ( .A(n591), .Y(n401) );
  INVX4 U472 ( .A(n337), .Y(n592) );
  INVX4 U473 ( .A(n339), .Y(n586) );
  BUFX4 U474 ( .A(n406), .Y(n407) );
  XNOR2X1 U475 ( .A(\A<14> ), .B(n404), .Y(n437) );
  XNOR2X1 U476 ( .A(\A<13> ), .B(n371), .Y(n409) );
  XNOR2X1 U477 ( .A(\A<12> ), .B(n359), .Y(n459) );
  INVX2 U478 ( .A(n459), .Y(n618) );
  XNOR2X1 U479 ( .A(\A<11> ), .B(n404), .Y(n506) );
  XNOR2X1 U480 ( .A(\A<9> ), .B(n404), .Y(n472) );
  XNOR2X1 U481 ( .A(\A<7> ), .B(n404), .Y(n410) );
  XNOR2X1 U482 ( .A(n404), .B(\A<6> ), .Y(n453) );
  XNOR2X1 U483 ( .A(n404), .B(\A<5> ), .Y(n411) );
  XNOR2X1 U484 ( .A(\A<4> ), .B(n404), .Y(n412) );
  XNOR2X1 U485 ( .A(n30), .B(\A<2> ), .Y(n413) );
  XNOR2X1 U486 ( .A(n30), .B(\A<1> ), .Y(n414) );
  XNOR2X1 U487 ( .A(n405), .B(\A<0> ), .Y(n415) );
  XNOR2X1 U488 ( .A(\B<14> ), .B(n234), .Y(n416) );
  INVX2 U489 ( .A(n416), .Y(n615) );
  XNOR2X1 U490 ( .A(\B<9> ), .B(n379), .Y(n614) );
  XNOR2X1 U491 ( .A(n15), .B(n239), .Y(n419) );
  XNOR2X1 U492 ( .A(\B<4> ), .B(n358), .Y(n420) );
  INVX2 U493 ( .A(n420), .Y(n610) );
  XNOR2X1 U494 ( .A(\B<3> ), .B(n403), .Y(n421) );
  XNOR2X1 U495 ( .A(n364), .B(n403), .Y(n422) );
  XNOR2X1 U496 ( .A(\B<0> ), .B(invB), .Y(n423) );
  XNOR2X1 U497 ( .A(n385), .B(n368), .Y(n424) );
  NOR3X1 U498 ( .A(n230), .B(n406), .C(n232), .Y(n591) );
  XNOR2X1 U499 ( .A(n388), .B(n606), .Y(n561) );
  INVX2 U500 ( .A(n406), .Y(n429) );
  NAND3X1 U501 ( .A(\Op<3> ), .B(n429), .C(n425), .Y(n583) );
  OR2X2 U502 ( .A(n201), .B(n375), .Y(n426) );
  INVX2 U503 ( .A(n426), .Y(n435) );
  NAND3X1 U504 ( .A(\Op<1> ), .B(n435), .C(n427), .Y(n588) );
  NAND3X1 U505 ( .A(n7), .B(n435), .C(n428), .Y(n512) );
  AND2X2 U506 ( .A(n407), .B(\A<0> ), .Y(n430) );
  AOI21X1 U507 ( .A(\B<15> ), .B(n52), .C(n430), .Y(n431) );
  OAI21X1 U508 ( .A(n345), .B(n533), .C(n252), .Y(n432) );
  AOI21X1 U509 ( .A(n388), .B(n170), .C(n432), .Y(n433) );
  OAI21X1 U510 ( .A(n561), .B(n402), .C(n101), .Y(n434) );
  AOI21X1 U511 ( .A(\shift_out<15> ), .B(n401), .C(n434), .Y(n436) );
  OR2X2 U512 ( .A(n7), .B(\Op<1> ), .Y(n555) );
  XNOR2X1 U513 ( .A(n615), .B(n620), .Y(n560) );
  AND2X2 U514 ( .A(n407), .B(\A<1> ), .Y(n438) );
  AOI21X1 U515 ( .A(\B<14> ), .B(n52), .C(n438), .Y(n439) );
  OAI21X1 U516 ( .A(n345), .B(n531), .C(n253), .Y(n440) );
  AOI21X1 U517 ( .A(n376), .B(n172), .C(n440), .Y(n441) );
  OAI21X1 U518 ( .A(n560), .B(n402), .C(n102), .Y(n442) );
  AOI21X1 U519 ( .A(\shift_out<14> ), .B(n401), .C(n442), .Y(n443) );
  INVX2 U520 ( .A(n402), .Y(n508) );
  XNOR2X1 U521 ( .A(n598), .B(n399), .Y(n574) );
  NAND3X1 U522 ( .A(n586), .B(n399), .C(n598), .Y(n444) );
  AOI21X1 U523 ( .A(n508), .B(n445), .C(n151), .Y(n446) );
  NAND3X1 U524 ( .A(n165), .B(n309), .C(n56), .Y(n447) );
  AOI21X1 U525 ( .A(n401), .B(\shift_out<1> ), .C(n282), .Y(n448) );
  XNOR2X1 U526 ( .A(n611), .B(n382), .Y(n571) );
  AOI21X1 U527 ( .A(n406), .B(\A<10> ), .C(n153), .Y(n449) );
  OAI21X1 U528 ( .A(n338), .B(n450), .C(n254), .Y(n452) );
  NAND3X1 U529 ( .A(n586), .B(n611), .C(n381), .Y(n451) );
  XNOR2X1 U530 ( .A(n240), .B(n234), .Y(n455) );
  XNOR2X1 U531 ( .A(n455), .B(n360), .Y(n578) );
  AOI22X1 U532 ( .A(n508), .B(n454), .C(n592), .D(\sum<6> ), .Y(n458) );
  NAND3X1 U533 ( .A(n604), .B(n586), .C(n612), .Y(n456) );
  AOI21X1 U534 ( .A(n401), .B(\shift_out<6> ), .C(n284), .Y(n457) );
  AND2X2 U535 ( .A(\A<4> ), .B(n344), .Y(n460) );
  AOI21X1 U536 ( .A(n17), .B(n303), .C(n460), .Y(n463) );
  AOI22X1 U537 ( .A(n18), .B(n52), .C(n401), .D(\shift_out<12> ), .Y(n462) );
  XNOR2X1 U538 ( .A(n17), .B(n618), .Y(n559) );
  OAI21X1 U539 ( .A(n559), .B(n402), .C(n111), .Y(n461) );
  AOI22X1 U540 ( .A(n508), .B(n348), .C(n592), .D(\sum<13> ), .Y(n466) );
  NAND3X1 U541 ( .A(n619), .B(n586), .C(n397), .Y(n464) );
  OAI21X1 U542 ( .A(n346), .B(n519), .C(n103), .Y(n465) );
  NAND3X1 U543 ( .A(n297), .B(n214), .C(n212), .Y(\Out<13> ) );
  AOI22X1 U544 ( .A(\B<8> ), .B(n52), .C(\shift_out<8> ), .D(n401), .Y(n471)
         );
  XNOR2X1 U545 ( .A(n242), .B(n215), .Y(n565) );
  OAI21X1 U546 ( .A(n565), .B(n402), .C(n260), .Y(n467) );
  AOI21X1 U547 ( .A(\sum<8> ), .B(n592), .C(n467), .Y(n470) );
  AND2X2 U548 ( .A(\A<0> ), .B(n344), .Y(n468) );
  AOI21X1 U549 ( .A(n243), .B(n305), .C(n468), .Y(n469) );
  XNOR2X1 U550 ( .A(\B<9> ), .B(n358), .Y(n474) );
  XNOR2X1 U551 ( .A(n474), .B(n350), .Y(n564) );
  INVX2 U552 ( .A(n564), .Y(n473) );
  AOI22X1 U553 ( .A(n508), .B(n473), .C(n592), .D(\sum<9> ), .Y(n479) );
  NAND3X1 U554 ( .A(n616), .B(n586), .C(n475), .Y(n476) );
  OAI21X1 U555 ( .A(n346), .B(n523), .C(n104), .Y(n477) );
  INVX2 U556 ( .A(\sum<4> ), .Y(n481) );
  XNOR2X1 U557 ( .A(n610), .B(n244), .Y(n570) );
  AOI21X1 U558 ( .A(n406), .B(\A<11> ), .C(n155), .Y(n480) );
  OAI21X1 U559 ( .A(n338), .B(n481), .C(n255), .Y(n484) );
  NAND3X1 U560 ( .A(n586), .B(n610), .C(n244), .Y(n482) );
  XNOR2X1 U561 ( .A(n608), .B(n355), .Y(n572) );
  NAND3X1 U562 ( .A(n608), .B(n586), .C(n355), .Y(n485) );
  AOI21X1 U563 ( .A(\B<2> ), .B(n343), .C(n157), .Y(n486) );
  OAI21X1 U564 ( .A(n572), .B(n402), .C(n105), .Y(n487) );
  AOI21X1 U565 ( .A(\sum<2> ), .B(n592), .C(n487), .Y(n488) );
  XNOR2X1 U566 ( .A(n609), .B(n601), .Y(n573) );
  AOI21X1 U567 ( .A(n406), .B(\A<12> ), .C(n159), .Y(n489) );
  OAI21X1 U568 ( .A(n338), .B(n490), .C(n256), .Y(n492) );
  NAND3X1 U569 ( .A(n586), .B(n601), .C(n609), .Y(n491) );
  XNOR2X1 U570 ( .A(n613), .B(n349), .Y(n577) );
  NAND3X1 U571 ( .A(n349), .B(n586), .C(n365), .Y(n493) );
  AOI21X1 U572 ( .A(n357), .B(n341), .C(n161), .Y(n494) );
  OAI21X1 U573 ( .A(n577), .B(n402), .C(n106), .Y(n495) );
  AOI21X1 U574 ( .A(\shift_out<7> ), .B(n401), .C(n495), .Y(n496) );
  XNOR2X1 U575 ( .A(n29), .B(n233), .Y(n498) );
  XNOR2X1 U576 ( .A(n498), .B(n497), .Y(n562) );
  INVX2 U577 ( .A(n498), .Y(n502) );
  AND2X2 U578 ( .A(n407), .B(\A<5> ), .Y(n499) );
  AOI21X1 U579 ( .A(n29), .B(n52), .C(n499), .Y(n500) );
  OAI21X1 U580 ( .A(n346), .B(n521), .C(n257), .Y(n501) );
  AOI21X1 U581 ( .A(n60), .B(n502), .C(n501), .Y(n503) );
  OAI21X1 U582 ( .A(n562), .B(n402), .C(n107), .Y(n504) );
  AOI21X1 U583 ( .A(\shift_out<10> ), .B(n401), .C(n504), .Y(n505) );
  NAND3X1 U584 ( .A(n11), .B(n316), .C(n167), .Y(n597) );
  XNOR2X1 U585 ( .A(n509), .B(n353), .Y(n563) );
  INVX2 U586 ( .A(n563), .Y(n507) );
  AOI22X1 U587 ( .A(n508), .B(n507), .C(\shift_out<11> ), .D(n401), .Y(n515)
         );
  INVX2 U588 ( .A(n509), .Y(n510) );
  NAND3X1 U589 ( .A(n617), .B(n586), .C(n510), .Y(n511) );
  OAI21X1 U590 ( .A(n345), .B(n525), .C(n108), .Y(n513) );
  AOI21X1 U591 ( .A(n373), .B(n52), .C(n513), .Y(n514) );
  AOI21X1 U592 ( .A(\B<15> ), .B(n516), .C(n222), .Y(n557) );
  AOI21X1 U593 ( .A(n518), .B(\A<6> ), .C(n163), .Y(n530) );
  AOI22X1 U594 ( .A(\B<4> ), .B(n520), .C(\B<5> ), .D(n519), .Y(n529) );
  AOI22X1 U595 ( .A(n352), .B(n523), .C(\B<0> ), .D(n522), .Y(n524) );
  AOI21X1 U596 ( .A(n526), .B(\A<4> ), .C(n286), .Y(n527) );
  OAI21X1 U597 ( .A(n307), .B(n180), .C(n223), .Y(n528) );
  AOI22X1 U598 ( .A(\B<7> ), .B(n533), .C(\B<6> ), .D(n531), .Y(n535) );
  OAI21X1 U599 ( .A(n533), .B(n357), .C(n113), .Y(n534) );
  AOI21X1 U600 ( .A(n300), .B(n174), .C(n534), .Y(n540) );
  INVX2 U601 ( .A(\A<8> ), .Y(n536) );
  OAI21X1 U602 ( .A(\A<9> ), .B(n537), .C(n262), .Y(n539) );
  AOI21X1 U603 ( .A(n537), .B(\A<9> ), .C(n66), .Y(n538) );
  OAI21X1 U604 ( .A(n175), .B(n539), .C(n258), .Y(n546) );
  AOI22X1 U605 ( .A(n373), .B(n543), .C(n29), .D(n541), .Y(n545) );
  OAI21X1 U606 ( .A(n543), .B(n373), .C(n264), .Y(n544) );
  AOI21X1 U607 ( .A(n546), .B(n301), .C(n544), .Y(n552) );
  OAI21X1 U608 ( .A(\A<13> ), .B(n548), .C(n68), .Y(n551) );
  AOI22X1 U609 ( .A(\A<14> ), .B(n549), .C(n548), .D(\A<13> ), .Y(n550) );
  OAI21X1 U610 ( .A(n176), .B(n551), .C(n251), .Y(n554) );
  AND2X2 U611 ( .A(n375), .B(n555), .Y(n556) );
  AND2X2 U612 ( .A(n561), .B(n560), .Y(n568) );
  INVX2 U613 ( .A(n562), .Y(n567) );
  NAND3X1 U614 ( .A(n565), .B(n564), .C(n563), .Y(n566) );
  XNOR2X1 U615 ( .A(n393), .B(n366), .Y(n589) );
  AND2X2 U616 ( .A(n589), .B(n7), .Y(n576) );
  AND2X2 U617 ( .A(n573), .B(n572), .Y(n575) );
  NAND3X1 U618 ( .A(n576), .B(n575), .C(n574), .Y(n579) );
  NOR3X1 U619 ( .A(n184), .B(n188), .C(n325), .Y(n580) );
  NAND3X1 U620 ( .A(n164), .B(n331), .C(n582), .Y(n585) );
  NAND3X1 U621 ( .A(n586), .B(n366), .C(n607), .Y(n587) );
  OAI21X1 U622 ( .A(n589), .B(n402), .C(n109), .Y(n590) );
  AOI21X1 U623 ( .A(n235), .B(n341), .C(n590), .Y(n594) );
  AOI22X1 U624 ( .A(\sum<0> ), .B(n592), .C(n401), .D(\shift_out<0> ), .Y(n593) );
  NOR3X1 U625 ( .A(n203), .B(n228), .C(n186), .Y(n595) );
  NAND3X1 U626 ( .A(n323), .B(n318), .C(n595), .Y(n596) );
  NOR3X1 U627 ( .A(n191), .B(n183), .C(n196), .Y(zero) );
  NOR2X1 U628 ( .A(n331), .B(n281), .Y(Ofl) );
  OR2X2 U629 ( .A(n148), .B(n199), .Y(\Out<0> ) );
endmodule


module adder_1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , 
        \A<9> , \A<8> , \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , 
        \A<0> }), .B({\B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , 
        \B<9> , \B<8> , \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , 
        \B<0> }), Cin, Overflow, Cout, .Sum({\Sum<15> , \Sum<14> , \Sum<13> , 
        \Sum<12> , \Sum<11> , \Sum<10> , \Sum<9> , \Sum<8> , \Sum<7> , 
        \Sum<6> , \Sum<5> , \Sum<4> , \Sum<3> , \Sum<2> , \Sum<1> , \Sum<0> })
 );
  input \A<15> , \A<14> , \A<13> , \A<12> , \A<11> , \A<10> , \A<9> , \A<8> ,
         \A<7> , \A<6> , \A<5> , \A<4> , \A<3> , \A<2> , \A<1> , \A<0> ,
         \B<15> , \B<14> , \B<13> , \B<12> , \B<11> , \B<10> , \B<9> , \B<8> ,
         \B<7> , \B<6> , \B<5> , \B<4> , \B<3> , \B<2> , \B<1> , \B<0> , Cin;
  output Overflow, Cout, \Sum<15> , \Sum<14> , \Sum<13> , \Sum<12> , \Sum<11> ,
         \Sum<10> , \Sum<9> , \Sum<8> , \Sum<7> , \Sum<6> , \Sum<5> , \Sum<4> ,
         \Sum<3> , \Sum<2> , \Sum<1> , \Sum<0> ;
  wire   c12, p12, g12, c8, p8, g8, c4, p4, g4, p0, g0, n2;

  FAX1 U1 ( .A(\B<15> ), .B(\A<15> ), .C(n2), .YC(), .YS(Overflow) );
  XOR2X1 U2 ( .A(\Sum<15> ), .B(Cout), .Y(n2) );
  cla_4_7 add1 ( .A({\A<15> , \A<14> , \A<13> , \A<12> }), .B({\B<15> , 
        \B<14> , \B<13> , \B<12> }), .Cin(c12), .p(p12), .g(g12), .S({
        \Sum<15> , \Sum<14> , \Sum<13> , \Sum<12> }), .Cout() );
  cla_4_6 add2 ( .A({\A<11> , \A<10> , \A<9> , \A<8> }), .B({\B<11> , \B<10> , 
        \B<9> , \B<8> }), .Cin(c8), .p(p8), .g(g8), .S({\Sum<11> , \Sum<10> , 
        \Sum<9> , \Sum<8> }), .Cout() );
  cla_4_5 add3 ( .A({\A<7> , \A<6> , \A<5> , \A<4> }), .B({\B<7> , \B<6> , 
        \B<5> , \B<4> }), .Cin(c4), .p(p4), .g(g4), .S({\Sum<7> , \Sum<6> , 
        \Sum<5> , \Sum<4> }), .Cout() );
  cla_4_4 add4 ( .A({\A<3> , \A<2> , \A<1> , \A<0> }), .B({\B<3> , \B<2> , 
        \B<1> , \B<0> }), .Cin(Cin), .p(p0), .g(g0), .S({\Sum<3> , \Sum<2> , 
        \Sum<1> , \Sum<0> }), .Cout() );
  groupcla_13 cla ( .p({p12, p8, p4, p0}), .g({g12, g8, g4, g0}), .Cin(Cin), 
        .c({Cout, c12, c8, c4}), .pg(), .gg() );
endmodule


module memory2c_0 ( .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), .addr({
        \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , 
        \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), enable, wr, createdump, 
        clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<15> , \addr<14> ,
         \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> ,
         \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , enable, wr, createdump, clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N177, N178, N179, N180, N181, N182, \mem<0><7> , \mem<0><6> ,
         \mem<0><5> , \mem<0><4> , \mem<0><3> , \mem<0><2> , \mem<0><1> ,
         \mem<0><0> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><7> ,
         \mem<2><6> , \mem<2><5> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><7> , \mem<3><6> , \mem<3><5> ,
         \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> , \mem<3><0> ,
         \mem<4><7> , \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> ,
         \mem<4><2> , \mem<4><1> , \mem<4><0> , \mem<5><7> , \mem<5><6> ,
         \mem<5><5> , \mem<5><4> , \mem<5><3> , \mem<5><2> , \mem<5><1> ,
         \mem<5><0> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><7> ,
         \mem<7><6> , \mem<7><5> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><7> , \mem<8><6> , \mem<8><5> ,
         \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> , \mem<8><0> ,
         \mem<9><7> , \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> ,
         \mem<9><2> , \mem<9><1> , \mem<9><0> , \mem<10><7> , \mem<10><6> ,
         \mem<10><5> , \mem<10><4> , \mem<10><3> , \mem<10><2> , \mem<10><1> ,
         \mem<10><0> , \mem<11><7> , \mem<11><6> , \mem<11><5> , \mem<11><4> ,
         \mem<11><3> , \mem<11><2> , \mem<11><1> , \mem<11><0> , \mem<12><7> ,
         \mem<12><6> , \mem<12><5> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><7> , \mem<13><6> , \mem<13><5> ,
         \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> , \mem<13><0> ,
         \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> , \mem<14><3> ,
         \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><7> ,
         \mem<17><6> , \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><7> , \mem<18><6> , \mem<18><5> ,
         \mem<18><4> , \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> ,
         \mem<19><7> , \mem<19><6> , \mem<19><5> , \mem<19><4> , \mem<19><3> ,
         \mem<19><2> , \mem<19><1> , \mem<19><0> , \mem<20><7> , \mem<20><6> ,
         \mem<20><5> , \mem<20><4> , \mem<20><3> , \mem<20><2> , \mem<20><1> ,
         \mem<20><0> , \mem<21><7> , \mem<21><6> , \mem<21><5> , \mem<21><4> ,
         \mem<21><3> , \mem<21><2> , \mem<21><1> , \mem<21><0> , \mem<22><7> ,
         \mem<22><6> , \mem<22><5> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><7> , \mem<23><6> , \mem<23><5> ,
         \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> , \mem<23><0> ,
         \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> , \mem<24><3> ,
         \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><7> ,
         \mem<27><6> , \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><7> , \mem<28><6> , \mem<28><5> ,
         \mem<28><4> , \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> ,
         \mem<29><7> , \mem<29><6> , \mem<29><5> , \mem<29><4> , \mem<29><3> ,
         \mem<29><2> , \mem<29><1> , \mem<29><0> , \mem<30><7> , \mem<30><6> ,
         \mem<30><5> , \mem<30><4> , \mem<30><3> , \mem<30><2> , \mem<30><1> ,
         \mem<30><0> , \mem<31><7> , \mem<31><6> , \mem<31><5> , \mem<31><4> ,
         \mem<31><3> , \mem<31><2> , \mem<31><1> , \mem<31><0> , \mem<32><7> ,
         \mem<32><6> , \mem<32><5> , \mem<32><4> , \mem<32><3> , \mem<32><2> ,
         \mem<32><1> , \mem<32><0> , \mem<33><7> , \mem<33><6> , \mem<33><5> ,
         \mem<33><4> , \mem<33><3> , \mem<33><2> , \mem<33><1> , \mem<33><0> ,
         \mem<34><7> , \mem<34><6> , \mem<34><5> , \mem<34><4> , \mem<34><3> ,
         \mem<34><2> , \mem<34><1> , \mem<34><0> , \mem<35><7> , \mem<35><6> ,
         \mem<35><5> , \mem<35><4> , \mem<35><3> , \mem<35><2> , \mem<35><1> ,
         \mem<35><0> , \mem<36><7> , \mem<36><6> , \mem<36><5> , \mem<36><4> ,
         \mem<36><3> , \mem<36><2> , \mem<36><1> , \mem<36><0> , \mem<37><7> ,
         \mem<37><6> , \mem<37><5> , \mem<37><4> , \mem<37><3> , \mem<37><2> ,
         \mem<37><1> , \mem<37><0> , \mem<38><7> , \mem<38><6> , \mem<38><5> ,
         \mem<38><4> , \mem<38><3> , \mem<38><2> , \mem<38><1> , \mem<38><0> ,
         \mem<39><7> , \mem<39><6> , \mem<39><5> , \mem<39><4> , \mem<39><3> ,
         \mem<39><2> , \mem<39><1> , \mem<39><0> , \mem<40><7> , \mem<40><6> ,
         \mem<40><5> , \mem<40><4> , \mem<40><3> , \mem<40><2> , \mem<40><1> ,
         \mem<40><0> , \mem<41><7> , \mem<41><6> , \mem<41><5> , \mem<41><4> ,
         \mem<41><3> , \mem<41><2> , \mem<41><1> , \mem<41><0> , \mem<42><7> ,
         \mem<42><6> , \mem<42><5> , \mem<42><4> , \mem<42><3> , \mem<42><2> ,
         \mem<42><1> , \mem<42><0> , \mem<43><7> , \mem<43><6> , \mem<43><5> ,
         \mem<43><4> , \mem<43><3> , \mem<43><2> , \mem<43><1> , \mem<43><0> ,
         \mem<44><7> , \mem<44><6> , \mem<44><5> , \mem<44><4> , \mem<44><3> ,
         \mem<44><2> , \mem<44><1> , \mem<44><0> , \mem<45><7> , \mem<45><6> ,
         \mem<45><5> , \mem<45><4> , \mem<45><3> , \mem<45><2> , \mem<45><1> ,
         \mem<45><0> , \mem<46><7> , \mem<46><6> , \mem<46><5> , \mem<46><4> ,
         \mem<46><3> , \mem<46><2> , \mem<46><1> , \mem<46><0> , \mem<47><7> ,
         \mem<47><6> , \mem<47><5> , \mem<47><4> , \mem<47><3> , \mem<47><2> ,
         \mem<47><1> , \mem<47><0> , \mem<48><7> , \mem<48><6> , \mem<48><5> ,
         \mem<48><4> , \mem<48><3> , \mem<48><2> , \mem<48><1> , \mem<48><0> ,
         \mem<49><7> , \mem<49><6> , \mem<49><5> , \mem<49><4> , \mem<49><3> ,
         \mem<49><2> , \mem<49><1> , \mem<49><0> , \mem<50><7> , \mem<50><6> ,
         \mem<50><5> , \mem<50><4> , \mem<50><3> , \mem<50><2> , \mem<50><1> ,
         \mem<50><0> , \mem<51><7> , \mem<51><6> , \mem<51><5> , \mem<51><4> ,
         \mem<51><3> , \mem<51><2> , \mem<51><1> , \mem<51><0> , \mem<52><7> ,
         \mem<52><6> , \mem<52><5> , \mem<52><4> , \mem<52><3> , \mem<52><2> ,
         \mem<52><1> , \mem<52><0> , \mem<53><7> , \mem<53><6> , \mem<53><5> ,
         \mem<53><4> , \mem<53><3> , \mem<53><2> , \mem<53><1> , \mem<53><0> ,
         \mem<54><7> , \mem<54><6> , \mem<54><5> , \mem<54><4> , \mem<54><3> ,
         \mem<54><2> , \mem<54><1> , \mem<54><0> , \mem<55><7> , \mem<55><6> ,
         \mem<55><5> , \mem<55><4> , \mem<55><3> , \mem<55><2> , \mem<55><1> ,
         \mem<55><0> , \mem<56><7> , \mem<56><6> , \mem<56><5> , \mem<56><4> ,
         \mem<56><3> , \mem<56><2> , \mem<56><1> , \mem<56><0> , \mem<57><7> ,
         \mem<57><6> , \mem<57><5> , \mem<57><4> , \mem<57><3> , \mem<57><2> ,
         \mem<57><1> , \mem<57><0> , \mem<58><7> , \mem<58><6> , \mem<58><5> ,
         \mem<58><4> , \mem<58><3> , \mem<58><2> , \mem<58><1> , \mem<58><0> ,
         \mem<59><7> , \mem<59><6> , \mem<59><5> , \mem<59><4> , \mem<59><3> ,
         \mem<59><2> , \mem<59><1> , \mem<59><0> , \mem<60><7> , \mem<60><6> ,
         \mem<60><5> , \mem<60><4> , \mem<60><3> , \mem<60><2> , \mem<60><1> ,
         \mem<60><0> , \mem<61><7> , \mem<61><6> , \mem<61><5> , \mem<61><4> ,
         \mem<61><3> , \mem<61><2> , \mem<61><1> , \mem<61><0> , \mem<62><7> ,
         \mem<62><6> , \mem<62><5> , \mem<62><4> , \mem<62><3> , \mem<62><2> ,
         \mem<62><1> , \mem<62><0> , \mem<63><7> , \mem<63><6> , \mem<63><5> ,
         \mem<63><4> , \mem<63><3> , \mem<63><2> , \mem<63><1> , \mem<63><0> ,
         N185, N186, N187, N188, N189, N190, N191, N192, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n568, n569, n571, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989;
  assign N177 = \addr<0> ;
  assign N178 = \addr<1> ;
  assign N179 = \addr<2> ;
  assign N180 = \addr<3> ;
  assign N181 = \addr<4> ;
  assign N182 = \addr<5> ;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n6478), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n6479), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n6480), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n6481), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n6482), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n6483), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n6484), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n6485), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n6486), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n6487), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n6488), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n6489), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n6490), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n6491), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n6492), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n6493), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n6494), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n6495), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n6496), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n6497), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n6498), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n6499), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n6500), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n6501), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n6502), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n6503), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n6504), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n6505), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n6506), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n6507), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n6508), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n6509), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n6510), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n6511), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n6512), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n6513), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n6514), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n6515), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n6516), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n6517), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n6518), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n6519), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n6520), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n6521), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n6522), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n6523), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n6524), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n6525), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n6526), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n6527), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n6528), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n6529), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n6530), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n6531), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n6532), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n6533), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n6534), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n6535), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n6536), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n6537), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n6538), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n6539), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n6540), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n6541), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n6542), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n6543), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n6544), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n6545), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n6546), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n6547), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n6548), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n6549), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n6550), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n6551), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n6552), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n6553), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n6554), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n6555), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n6556), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n6557), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n6558), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n6559), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n6560), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n6561), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n6562), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n6563), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n6564), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n6565), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n6566), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n6567), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n6568), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n6569), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n6570), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n6571), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n6572), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n6573), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n6574), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n6575), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n6576), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n6577), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n6578), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n6579), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n6580), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n6581), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n6582), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n6583), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n6584), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n6585), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n6586), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n6587), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n6588), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n6589), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n6590), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n6591), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n6592), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n6593), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n6594), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n6595), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n6596), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n6597), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n6598), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n6599), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n6600), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n6601), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n6602), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n6603), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n6604), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n6605), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n6606), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n6607), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n6608), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n6609), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n6610), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n6611), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n6612), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n6613), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n6614), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n6615), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n6616), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n6617), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n6618), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n6619), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n6620), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n6621), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n6622), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n6623), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n6624), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n6625), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n6626), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n6627), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n6628), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n6629), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n6630), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n6631), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n6632), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n6633), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n6634), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n6635), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n6636), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n6637), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n6638), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n6639), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n6640), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n6641), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n6642), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n6643), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n6644), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n6645), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n6646), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n6647), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n6648), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n6649), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n6650), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n6651), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n6652), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n6653), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n6654), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n6655), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n6656), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n6657), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n6658), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n6659), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n6660), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n6661), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n6662), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n6663), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n6664), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n6665), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n6666), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n6667), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n6668), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n6669), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n6670), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n6671), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n6672), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n6673), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n6674), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n6675), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n6676), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n6677), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n6678), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n6679), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n6680), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n6681), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n6682), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n6683), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n6684), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n6685), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n6686), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n6687), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n6688), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n6689), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n6690), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n6691), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n6692), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n6693), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n6694), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n6695), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n6696), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n6697), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n6698), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n6699), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n6700), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n6701), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n6702), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n6703), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n6704), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n6705), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n6706), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n6707), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n6708), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n6709), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n6710), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n6711), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n6712), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n6713), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n6714), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n6715), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n6716), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n6717), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n6718), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n6719), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n6720), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n6721), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n6722), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n6723), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n6724), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n6725), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n6726), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n6727), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n6728), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n6729), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n6730), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n6731), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n6732), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n6733), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n6734), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n6735), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n6736), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n6737), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n6738), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n6739), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n6740), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n6741), .CLK(clk), .Q(\mem<32><0> ) );
  DFFPOSX1 \mem_reg<33><7>  ( .D(n6742), .CLK(clk), .Q(\mem<33><7> ) );
  DFFPOSX1 \mem_reg<33><6>  ( .D(n6743), .CLK(clk), .Q(\mem<33><6> ) );
  DFFPOSX1 \mem_reg<33><5>  ( .D(n6744), .CLK(clk), .Q(\mem<33><5> ) );
  DFFPOSX1 \mem_reg<33><4>  ( .D(n6745), .CLK(clk), .Q(\mem<33><4> ) );
  DFFPOSX1 \mem_reg<33><3>  ( .D(n6746), .CLK(clk), .Q(\mem<33><3> ) );
  DFFPOSX1 \mem_reg<33><2>  ( .D(n6747), .CLK(clk), .Q(\mem<33><2> ) );
  DFFPOSX1 \mem_reg<33><1>  ( .D(n6748), .CLK(clk), .Q(\mem<33><1> ) );
  DFFPOSX1 \mem_reg<33><0>  ( .D(n6749), .CLK(clk), .Q(\mem<33><0> ) );
  DFFPOSX1 \mem_reg<34><7>  ( .D(n6750), .CLK(clk), .Q(\mem<34><7> ) );
  DFFPOSX1 \mem_reg<34><6>  ( .D(n6751), .CLK(clk), .Q(\mem<34><6> ) );
  DFFPOSX1 \mem_reg<34><5>  ( .D(n6752), .CLK(clk), .Q(\mem<34><5> ) );
  DFFPOSX1 \mem_reg<34><4>  ( .D(n6753), .CLK(clk), .Q(\mem<34><4> ) );
  DFFPOSX1 \mem_reg<34><3>  ( .D(n6754), .CLK(clk), .Q(\mem<34><3> ) );
  DFFPOSX1 \mem_reg<34><2>  ( .D(n6755), .CLK(clk), .Q(\mem<34><2> ) );
  DFFPOSX1 \mem_reg<34><1>  ( .D(n6756), .CLK(clk), .Q(\mem<34><1> ) );
  DFFPOSX1 \mem_reg<34><0>  ( .D(n6757), .CLK(clk), .Q(\mem<34><0> ) );
  DFFPOSX1 \mem_reg<35><7>  ( .D(n6758), .CLK(clk), .Q(\mem<35><7> ) );
  DFFPOSX1 \mem_reg<35><6>  ( .D(n6759), .CLK(clk), .Q(\mem<35><6> ) );
  DFFPOSX1 \mem_reg<35><5>  ( .D(n6760), .CLK(clk), .Q(\mem<35><5> ) );
  DFFPOSX1 \mem_reg<35><4>  ( .D(n6761), .CLK(clk), .Q(\mem<35><4> ) );
  DFFPOSX1 \mem_reg<35><3>  ( .D(n6762), .CLK(clk), .Q(\mem<35><3> ) );
  DFFPOSX1 \mem_reg<35><2>  ( .D(n6763), .CLK(clk), .Q(\mem<35><2> ) );
  DFFPOSX1 \mem_reg<35><1>  ( .D(n6764), .CLK(clk), .Q(\mem<35><1> ) );
  DFFPOSX1 \mem_reg<35><0>  ( .D(n6765), .CLK(clk), .Q(\mem<35><0> ) );
  DFFPOSX1 \mem_reg<36><7>  ( .D(n6766), .CLK(clk), .Q(\mem<36><7> ) );
  DFFPOSX1 \mem_reg<36><6>  ( .D(n6767), .CLK(clk), .Q(\mem<36><6> ) );
  DFFPOSX1 \mem_reg<36><5>  ( .D(n6768), .CLK(clk), .Q(\mem<36><5> ) );
  DFFPOSX1 \mem_reg<36><4>  ( .D(n6769), .CLK(clk), .Q(\mem<36><4> ) );
  DFFPOSX1 \mem_reg<36><3>  ( .D(n6770), .CLK(clk), .Q(\mem<36><3> ) );
  DFFPOSX1 \mem_reg<36><2>  ( .D(n6771), .CLK(clk), .Q(\mem<36><2> ) );
  DFFPOSX1 \mem_reg<36><1>  ( .D(n6772), .CLK(clk), .Q(\mem<36><1> ) );
  DFFPOSX1 \mem_reg<36><0>  ( .D(n6773), .CLK(clk), .Q(\mem<36><0> ) );
  DFFPOSX1 \mem_reg<37><7>  ( .D(n6774), .CLK(clk), .Q(\mem<37><7> ) );
  DFFPOSX1 \mem_reg<37><6>  ( .D(n6775), .CLK(clk), .Q(\mem<37><6> ) );
  DFFPOSX1 \mem_reg<37><5>  ( .D(n6776), .CLK(clk), .Q(\mem<37><5> ) );
  DFFPOSX1 \mem_reg<37><4>  ( .D(n6777), .CLK(clk), .Q(\mem<37><4> ) );
  DFFPOSX1 \mem_reg<37><3>  ( .D(n6778), .CLK(clk), .Q(\mem<37><3> ) );
  DFFPOSX1 \mem_reg<37><2>  ( .D(n6779), .CLK(clk), .Q(\mem<37><2> ) );
  DFFPOSX1 \mem_reg<37><1>  ( .D(n6780), .CLK(clk), .Q(\mem<37><1> ) );
  DFFPOSX1 \mem_reg<37><0>  ( .D(n6781), .CLK(clk), .Q(\mem<37><0> ) );
  DFFPOSX1 \mem_reg<38><7>  ( .D(n6782), .CLK(clk), .Q(\mem<38><7> ) );
  DFFPOSX1 \mem_reg<38><6>  ( .D(n6783), .CLK(clk), .Q(\mem<38><6> ) );
  DFFPOSX1 \mem_reg<38><5>  ( .D(n6784), .CLK(clk), .Q(\mem<38><5> ) );
  DFFPOSX1 \mem_reg<38><4>  ( .D(n6785), .CLK(clk), .Q(\mem<38><4> ) );
  DFFPOSX1 \mem_reg<38><3>  ( .D(n6786), .CLK(clk), .Q(\mem<38><3> ) );
  DFFPOSX1 \mem_reg<38><2>  ( .D(n6787), .CLK(clk), .Q(\mem<38><2> ) );
  DFFPOSX1 \mem_reg<38><1>  ( .D(n6788), .CLK(clk), .Q(\mem<38><1> ) );
  DFFPOSX1 \mem_reg<38><0>  ( .D(n6789), .CLK(clk), .Q(\mem<38><0> ) );
  DFFPOSX1 \mem_reg<39><7>  ( .D(n6790), .CLK(clk), .Q(\mem<39><7> ) );
  DFFPOSX1 \mem_reg<39><6>  ( .D(n6791), .CLK(clk), .Q(\mem<39><6> ) );
  DFFPOSX1 \mem_reg<39><5>  ( .D(n6792), .CLK(clk), .Q(\mem<39><5> ) );
  DFFPOSX1 \mem_reg<39><4>  ( .D(n6793), .CLK(clk), .Q(\mem<39><4> ) );
  DFFPOSX1 \mem_reg<39><3>  ( .D(n6794), .CLK(clk), .Q(\mem<39><3> ) );
  DFFPOSX1 \mem_reg<39><2>  ( .D(n6795), .CLK(clk), .Q(\mem<39><2> ) );
  DFFPOSX1 \mem_reg<39><1>  ( .D(n6796), .CLK(clk), .Q(\mem<39><1> ) );
  DFFPOSX1 \mem_reg<39><0>  ( .D(n6797), .CLK(clk), .Q(\mem<39><0> ) );
  DFFPOSX1 \mem_reg<40><7>  ( .D(n6798), .CLK(clk), .Q(\mem<40><7> ) );
  DFFPOSX1 \mem_reg<40><6>  ( .D(n6799), .CLK(clk), .Q(\mem<40><6> ) );
  DFFPOSX1 \mem_reg<40><5>  ( .D(n6800), .CLK(clk), .Q(\mem<40><5> ) );
  DFFPOSX1 \mem_reg<40><4>  ( .D(n6801), .CLK(clk), .Q(\mem<40><4> ) );
  DFFPOSX1 \mem_reg<40><3>  ( .D(n6802), .CLK(clk), .Q(\mem<40><3> ) );
  DFFPOSX1 \mem_reg<40><2>  ( .D(n6803), .CLK(clk), .Q(\mem<40><2> ) );
  DFFPOSX1 \mem_reg<40><1>  ( .D(n6804), .CLK(clk), .Q(\mem<40><1> ) );
  DFFPOSX1 \mem_reg<40><0>  ( .D(n6805), .CLK(clk), .Q(\mem<40><0> ) );
  DFFPOSX1 \mem_reg<41><7>  ( .D(n6806), .CLK(clk), .Q(\mem<41><7> ) );
  DFFPOSX1 \mem_reg<41><6>  ( .D(n6807), .CLK(clk), .Q(\mem<41><6> ) );
  DFFPOSX1 \mem_reg<41><5>  ( .D(n6808), .CLK(clk), .Q(\mem<41><5> ) );
  DFFPOSX1 \mem_reg<41><4>  ( .D(n6809), .CLK(clk), .Q(\mem<41><4> ) );
  DFFPOSX1 \mem_reg<41><3>  ( .D(n6810), .CLK(clk), .Q(\mem<41><3> ) );
  DFFPOSX1 \mem_reg<41><2>  ( .D(n6811), .CLK(clk), .Q(\mem<41><2> ) );
  DFFPOSX1 \mem_reg<41><1>  ( .D(n6812), .CLK(clk), .Q(\mem<41><1> ) );
  DFFPOSX1 \mem_reg<41><0>  ( .D(n6813), .CLK(clk), .Q(\mem<41><0> ) );
  DFFPOSX1 \mem_reg<42><7>  ( .D(n6814), .CLK(clk), .Q(\mem<42><7> ) );
  DFFPOSX1 \mem_reg<42><6>  ( .D(n6815), .CLK(clk), .Q(\mem<42><6> ) );
  DFFPOSX1 \mem_reg<42><5>  ( .D(n6816), .CLK(clk), .Q(\mem<42><5> ) );
  DFFPOSX1 \mem_reg<42><4>  ( .D(n6817), .CLK(clk), .Q(\mem<42><4> ) );
  DFFPOSX1 \mem_reg<42><3>  ( .D(n6818), .CLK(clk), .Q(\mem<42><3> ) );
  DFFPOSX1 \mem_reg<42><2>  ( .D(n6819), .CLK(clk), .Q(\mem<42><2> ) );
  DFFPOSX1 \mem_reg<42><1>  ( .D(n6820), .CLK(clk), .Q(\mem<42><1> ) );
  DFFPOSX1 \mem_reg<42><0>  ( .D(n6821), .CLK(clk), .Q(\mem<42><0> ) );
  DFFPOSX1 \mem_reg<43><7>  ( .D(n6822), .CLK(clk), .Q(\mem<43><7> ) );
  DFFPOSX1 \mem_reg<43><6>  ( .D(n6823), .CLK(clk), .Q(\mem<43><6> ) );
  DFFPOSX1 \mem_reg<43><5>  ( .D(n6824), .CLK(clk), .Q(\mem<43><5> ) );
  DFFPOSX1 \mem_reg<43><4>  ( .D(n6825), .CLK(clk), .Q(\mem<43><4> ) );
  DFFPOSX1 \mem_reg<43><3>  ( .D(n6826), .CLK(clk), .Q(\mem<43><3> ) );
  DFFPOSX1 \mem_reg<43><2>  ( .D(n6827), .CLK(clk), .Q(\mem<43><2> ) );
  DFFPOSX1 \mem_reg<43><1>  ( .D(n6828), .CLK(clk), .Q(\mem<43><1> ) );
  DFFPOSX1 \mem_reg<43><0>  ( .D(n6829), .CLK(clk), .Q(\mem<43><0> ) );
  DFFPOSX1 \mem_reg<44><7>  ( .D(n6830), .CLK(clk), .Q(\mem<44><7> ) );
  DFFPOSX1 \mem_reg<44><6>  ( .D(n6831), .CLK(clk), .Q(\mem<44><6> ) );
  DFFPOSX1 \mem_reg<44><5>  ( .D(n6832), .CLK(clk), .Q(\mem<44><5> ) );
  DFFPOSX1 \mem_reg<44><4>  ( .D(n6833), .CLK(clk), .Q(\mem<44><4> ) );
  DFFPOSX1 \mem_reg<44><3>  ( .D(n6834), .CLK(clk), .Q(\mem<44><3> ) );
  DFFPOSX1 \mem_reg<44><2>  ( .D(n6835), .CLK(clk), .Q(\mem<44><2> ) );
  DFFPOSX1 \mem_reg<44><1>  ( .D(n6836), .CLK(clk), .Q(\mem<44><1> ) );
  DFFPOSX1 \mem_reg<44><0>  ( .D(n6837), .CLK(clk), .Q(\mem<44><0> ) );
  DFFPOSX1 \mem_reg<45><7>  ( .D(n6838), .CLK(clk), .Q(\mem<45><7> ) );
  DFFPOSX1 \mem_reg<45><6>  ( .D(n6839), .CLK(clk), .Q(\mem<45><6> ) );
  DFFPOSX1 \mem_reg<45><5>  ( .D(n6840), .CLK(clk), .Q(\mem<45><5> ) );
  DFFPOSX1 \mem_reg<45><4>  ( .D(n6841), .CLK(clk), .Q(\mem<45><4> ) );
  DFFPOSX1 \mem_reg<45><3>  ( .D(n6842), .CLK(clk), .Q(\mem<45><3> ) );
  DFFPOSX1 \mem_reg<45><2>  ( .D(n6843), .CLK(clk), .Q(\mem<45><2> ) );
  DFFPOSX1 \mem_reg<45><1>  ( .D(n6844), .CLK(clk), .Q(\mem<45><1> ) );
  DFFPOSX1 \mem_reg<45><0>  ( .D(n6845), .CLK(clk), .Q(\mem<45><0> ) );
  DFFPOSX1 \mem_reg<46><7>  ( .D(n6846), .CLK(clk), .Q(\mem<46><7> ) );
  DFFPOSX1 \mem_reg<46><6>  ( .D(n6847), .CLK(clk), .Q(\mem<46><6> ) );
  DFFPOSX1 \mem_reg<46><5>  ( .D(n6848), .CLK(clk), .Q(\mem<46><5> ) );
  DFFPOSX1 \mem_reg<46><4>  ( .D(n6849), .CLK(clk), .Q(\mem<46><4> ) );
  DFFPOSX1 \mem_reg<46><3>  ( .D(n6850), .CLK(clk), .Q(\mem<46><3> ) );
  DFFPOSX1 \mem_reg<46><2>  ( .D(n6851), .CLK(clk), .Q(\mem<46><2> ) );
  DFFPOSX1 \mem_reg<46><1>  ( .D(n6852), .CLK(clk), .Q(\mem<46><1> ) );
  DFFPOSX1 \mem_reg<46><0>  ( .D(n6853), .CLK(clk), .Q(\mem<46><0> ) );
  DFFPOSX1 \mem_reg<47><7>  ( .D(n6854), .CLK(clk), .Q(\mem<47><7> ) );
  DFFPOSX1 \mem_reg<47><6>  ( .D(n6855), .CLK(clk), .Q(\mem<47><6> ) );
  DFFPOSX1 \mem_reg<47><5>  ( .D(n6856), .CLK(clk), .Q(\mem<47><5> ) );
  DFFPOSX1 \mem_reg<47><4>  ( .D(n6857), .CLK(clk), .Q(\mem<47><4> ) );
  DFFPOSX1 \mem_reg<47><3>  ( .D(n6858), .CLK(clk), .Q(\mem<47><3> ) );
  DFFPOSX1 \mem_reg<47><2>  ( .D(n6859), .CLK(clk), .Q(\mem<47><2> ) );
  DFFPOSX1 \mem_reg<47><1>  ( .D(n6860), .CLK(clk), .Q(\mem<47><1> ) );
  DFFPOSX1 \mem_reg<47><0>  ( .D(n6861), .CLK(clk), .Q(\mem<47><0> ) );
  DFFPOSX1 \mem_reg<48><7>  ( .D(n6862), .CLK(clk), .Q(\mem<48><7> ) );
  DFFPOSX1 \mem_reg<48><6>  ( .D(n6863), .CLK(clk), .Q(\mem<48><6> ) );
  DFFPOSX1 \mem_reg<48><5>  ( .D(n6864), .CLK(clk), .Q(\mem<48><5> ) );
  DFFPOSX1 \mem_reg<48><4>  ( .D(n6865), .CLK(clk), .Q(\mem<48><4> ) );
  DFFPOSX1 \mem_reg<48><3>  ( .D(n6866), .CLK(clk), .Q(\mem<48><3> ) );
  DFFPOSX1 \mem_reg<48><2>  ( .D(n6867), .CLK(clk), .Q(\mem<48><2> ) );
  DFFPOSX1 \mem_reg<48><1>  ( .D(n6868), .CLK(clk), .Q(\mem<48><1> ) );
  DFFPOSX1 \mem_reg<48><0>  ( .D(n6869), .CLK(clk), .Q(\mem<48><0> ) );
  DFFPOSX1 \mem_reg<49><7>  ( .D(n6870), .CLK(clk), .Q(\mem<49><7> ) );
  DFFPOSX1 \mem_reg<49><6>  ( .D(n6871), .CLK(clk), .Q(\mem<49><6> ) );
  DFFPOSX1 \mem_reg<49><5>  ( .D(n6872), .CLK(clk), .Q(\mem<49><5> ) );
  DFFPOSX1 \mem_reg<49><4>  ( .D(n6873), .CLK(clk), .Q(\mem<49><4> ) );
  DFFPOSX1 \mem_reg<49><3>  ( .D(n6874), .CLK(clk), .Q(\mem<49><3> ) );
  DFFPOSX1 \mem_reg<49><2>  ( .D(n6875), .CLK(clk), .Q(\mem<49><2> ) );
  DFFPOSX1 \mem_reg<49><1>  ( .D(n6876), .CLK(clk), .Q(\mem<49><1> ) );
  DFFPOSX1 \mem_reg<49><0>  ( .D(n6877), .CLK(clk), .Q(\mem<49><0> ) );
  DFFPOSX1 \mem_reg<50><7>  ( .D(n6878), .CLK(clk), .Q(\mem<50><7> ) );
  DFFPOSX1 \mem_reg<50><6>  ( .D(n6879), .CLK(clk), .Q(\mem<50><6> ) );
  DFFPOSX1 \mem_reg<50><5>  ( .D(n6880), .CLK(clk), .Q(\mem<50><5> ) );
  DFFPOSX1 \mem_reg<50><4>  ( .D(n6881), .CLK(clk), .Q(\mem<50><4> ) );
  DFFPOSX1 \mem_reg<50><3>  ( .D(n6882), .CLK(clk), .Q(\mem<50><3> ) );
  DFFPOSX1 \mem_reg<50><2>  ( .D(n6883), .CLK(clk), .Q(\mem<50><2> ) );
  DFFPOSX1 \mem_reg<50><1>  ( .D(n6884), .CLK(clk), .Q(\mem<50><1> ) );
  DFFPOSX1 \mem_reg<50><0>  ( .D(n6885), .CLK(clk), .Q(\mem<50><0> ) );
  DFFPOSX1 \mem_reg<51><7>  ( .D(n6886), .CLK(clk), .Q(\mem<51><7> ) );
  DFFPOSX1 \mem_reg<51><6>  ( .D(n6887), .CLK(clk), .Q(\mem<51><6> ) );
  DFFPOSX1 \mem_reg<51><5>  ( .D(n6888), .CLK(clk), .Q(\mem<51><5> ) );
  DFFPOSX1 \mem_reg<51><4>  ( .D(n6889), .CLK(clk), .Q(\mem<51><4> ) );
  DFFPOSX1 \mem_reg<51><3>  ( .D(n6890), .CLK(clk), .Q(\mem<51><3> ) );
  DFFPOSX1 \mem_reg<51><2>  ( .D(n6891), .CLK(clk), .Q(\mem<51><2> ) );
  DFFPOSX1 \mem_reg<51><1>  ( .D(n6892), .CLK(clk), .Q(\mem<51><1> ) );
  DFFPOSX1 \mem_reg<51><0>  ( .D(n6893), .CLK(clk), .Q(\mem<51><0> ) );
  DFFPOSX1 \mem_reg<52><7>  ( .D(n6894), .CLK(clk), .Q(\mem<52><7> ) );
  DFFPOSX1 \mem_reg<52><6>  ( .D(n6895), .CLK(clk), .Q(\mem<52><6> ) );
  DFFPOSX1 \mem_reg<52><5>  ( .D(n6896), .CLK(clk), .Q(\mem<52><5> ) );
  DFFPOSX1 \mem_reg<52><4>  ( .D(n6897), .CLK(clk), .Q(\mem<52><4> ) );
  DFFPOSX1 \mem_reg<52><3>  ( .D(n6898), .CLK(clk), .Q(\mem<52><3> ) );
  DFFPOSX1 \mem_reg<52><2>  ( .D(n6899), .CLK(clk), .Q(\mem<52><2> ) );
  DFFPOSX1 \mem_reg<52><1>  ( .D(n6900), .CLK(clk), .Q(\mem<52><1> ) );
  DFFPOSX1 \mem_reg<52><0>  ( .D(n6901), .CLK(clk), .Q(\mem<52><0> ) );
  DFFPOSX1 \mem_reg<53><7>  ( .D(n6902), .CLK(clk), .Q(\mem<53><7> ) );
  DFFPOSX1 \mem_reg<53><6>  ( .D(n6903), .CLK(clk), .Q(\mem<53><6> ) );
  DFFPOSX1 \mem_reg<53><5>  ( .D(n6904), .CLK(clk), .Q(\mem<53><5> ) );
  DFFPOSX1 \mem_reg<53><4>  ( .D(n6905), .CLK(clk), .Q(\mem<53><4> ) );
  DFFPOSX1 \mem_reg<53><3>  ( .D(n6906), .CLK(clk), .Q(\mem<53><3> ) );
  DFFPOSX1 \mem_reg<53><2>  ( .D(n6907), .CLK(clk), .Q(\mem<53><2> ) );
  DFFPOSX1 \mem_reg<53><1>  ( .D(n6908), .CLK(clk), .Q(\mem<53><1> ) );
  DFFPOSX1 \mem_reg<53><0>  ( .D(n6909), .CLK(clk), .Q(\mem<53><0> ) );
  DFFPOSX1 \mem_reg<54><7>  ( .D(n6910), .CLK(clk), .Q(\mem<54><7> ) );
  DFFPOSX1 \mem_reg<54><6>  ( .D(n6911), .CLK(clk), .Q(\mem<54><6> ) );
  DFFPOSX1 \mem_reg<54><5>  ( .D(n6912), .CLK(clk), .Q(\mem<54><5> ) );
  DFFPOSX1 \mem_reg<54><4>  ( .D(n6913), .CLK(clk), .Q(\mem<54><4> ) );
  DFFPOSX1 \mem_reg<54><3>  ( .D(n6914), .CLK(clk), .Q(\mem<54><3> ) );
  DFFPOSX1 \mem_reg<54><2>  ( .D(n6915), .CLK(clk), .Q(\mem<54><2> ) );
  DFFPOSX1 \mem_reg<54><1>  ( .D(n6916), .CLK(clk), .Q(\mem<54><1> ) );
  DFFPOSX1 \mem_reg<54><0>  ( .D(n6917), .CLK(clk), .Q(\mem<54><0> ) );
  DFFPOSX1 \mem_reg<55><7>  ( .D(n6918), .CLK(clk), .Q(\mem<55><7> ) );
  DFFPOSX1 \mem_reg<55><6>  ( .D(n6919), .CLK(clk), .Q(\mem<55><6> ) );
  DFFPOSX1 \mem_reg<55><5>  ( .D(n6920), .CLK(clk), .Q(\mem<55><5> ) );
  DFFPOSX1 \mem_reg<55><4>  ( .D(n6921), .CLK(clk), .Q(\mem<55><4> ) );
  DFFPOSX1 \mem_reg<55><3>  ( .D(n6922), .CLK(clk), .Q(\mem<55><3> ) );
  DFFPOSX1 \mem_reg<55><2>  ( .D(n6923), .CLK(clk), .Q(\mem<55><2> ) );
  DFFPOSX1 \mem_reg<55><1>  ( .D(n6924), .CLK(clk), .Q(\mem<55><1> ) );
  DFFPOSX1 \mem_reg<55><0>  ( .D(n6925), .CLK(clk), .Q(\mem<55><0> ) );
  DFFPOSX1 \mem_reg<56><7>  ( .D(n6926), .CLK(clk), .Q(\mem<56><7> ) );
  DFFPOSX1 \mem_reg<56><6>  ( .D(n6927), .CLK(clk), .Q(\mem<56><6> ) );
  DFFPOSX1 \mem_reg<56><5>  ( .D(n6928), .CLK(clk), .Q(\mem<56><5> ) );
  DFFPOSX1 \mem_reg<56><4>  ( .D(n6929), .CLK(clk), .Q(\mem<56><4> ) );
  DFFPOSX1 \mem_reg<56><3>  ( .D(n6930), .CLK(clk), .Q(\mem<56><3> ) );
  DFFPOSX1 \mem_reg<56><2>  ( .D(n6931), .CLK(clk), .Q(\mem<56><2> ) );
  DFFPOSX1 \mem_reg<56><1>  ( .D(n6932), .CLK(clk), .Q(\mem<56><1> ) );
  DFFPOSX1 \mem_reg<56><0>  ( .D(n6933), .CLK(clk), .Q(\mem<56><0> ) );
  DFFPOSX1 \mem_reg<57><7>  ( .D(n6934), .CLK(clk), .Q(\mem<57><7> ) );
  DFFPOSX1 \mem_reg<57><6>  ( .D(n6935), .CLK(clk), .Q(\mem<57><6> ) );
  DFFPOSX1 \mem_reg<57><5>  ( .D(n6936), .CLK(clk), .Q(\mem<57><5> ) );
  DFFPOSX1 \mem_reg<57><4>  ( .D(n6937), .CLK(clk), .Q(\mem<57><4> ) );
  DFFPOSX1 \mem_reg<57><3>  ( .D(n6938), .CLK(clk), .Q(\mem<57><3> ) );
  DFFPOSX1 \mem_reg<57><2>  ( .D(n6939), .CLK(clk), .Q(\mem<57><2> ) );
  DFFPOSX1 \mem_reg<57><1>  ( .D(n6940), .CLK(clk), .Q(\mem<57><1> ) );
  DFFPOSX1 \mem_reg<57><0>  ( .D(n6941), .CLK(clk), .Q(\mem<57><0> ) );
  DFFPOSX1 \mem_reg<58><7>  ( .D(n6942), .CLK(clk), .Q(\mem<58><7> ) );
  DFFPOSX1 \mem_reg<58><6>  ( .D(n6943), .CLK(clk), .Q(\mem<58><6> ) );
  DFFPOSX1 \mem_reg<58><5>  ( .D(n6944), .CLK(clk), .Q(\mem<58><5> ) );
  DFFPOSX1 \mem_reg<58><4>  ( .D(n6945), .CLK(clk), .Q(\mem<58><4> ) );
  DFFPOSX1 \mem_reg<58><3>  ( .D(n6946), .CLK(clk), .Q(\mem<58><3> ) );
  DFFPOSX1 \mem_reg<58><2>  ( .D(n6947), .CLK(clk), .Q(\mem<58><2> ) );
  DFFPOSX1 \mem_reg<58><1>  ( .D(n6948), .CLK(clk), .Q(\mem<58><1> ) );
  DFFPOSX1 \mem_reg<58><0>  ( .D(n6949), .CLK(clk), .Q(\mem<58><0> ) );
  DFFPOSX1 \mem_reg<59><7>  ( .D(n6950), .CLK(clk), .Q(\mem<59><7> ) );
  DFFPOSX1 \mem_reg<59><6>  ( .D(n6951), .CLK(clk), .Q(\mem<59><6> ) );
  DFFPOSX1 \mem_reg<59><5>  ( .D(n6952), .CLK(clk), .Q(\mem<59><5> ) );
  DFFPOSX1 \mem_reg<59><4>  ( .D(n6953), .CLK(clk), .Q(\mem<59><4> ) );
  DFFPOSX1 \mem_reg<59><3>  ( .D(n6954), .CLK(clk), .Q(\mem<59><3> ) );
  DFFPOSX1 \mem_reg<59><2>  ( .D(n6955), .CLK(clk), .Q(\mem<59><2> ) );
  DFFPOSX1 \mem_reg<59><1>  ( .D(n6956), .CLK(clk), .Q(\mem<59><1> ) );
  DFFPOSX1 \mem_reg<59><0>  ( .D(n6957), .CLK(clk), .Q(\mem<59><0> ) );
  DFFPOSX1 \mem_reg<60><7>  ( .D(n6958), .CLK(clk), .Q(\mem<60><7> ) );
  DFFPOSX1 \mem_reg<60><6>  ( .D(n6959), .CLK(clk), .Q(\mem<60><6> ) );
  DFFPOSX1 \mem_reg<60><5>  ( .D(n6960), .CLK(clk), .Q(\mem<60><5> ) );
  DFFPOSX1 \mem_reg<60><4>  ( .D(n6961), .CLK(clk), .Q(\mem<60><4> ) );
  DFFPOSX1 \mem_reg<60><3>  ( .D(n6962), .CLK(clk), .Q(\mem<60><3> ) );
  DFFPOSX1 \mem_reg<60><2>  ( .D(n6963), .CLK(clk), .Q(\mem<60><2> ) );
  DFFPOSX1 \mem_reg<60><1>  ( .D(n6964), .CLK(clk), .Q(\mem<60><1> ) );
  DFFPOSX1 \mem_reg<60><0>  ( .D(n6965), .CLK(clk), .Q(\mem<60><0> ) );
  DFFPOSX1 \mem_reg<61><7>  ( .D(n6966), .CLK(clk), .Q(\mem<61><7> ) );
  DFFPOSX1 \mem_reg<61><6>  ( .D(n6967), .CLK(clk), .Q(\mem<61><6> ) );
  DFFPOSX1 \mem_reg<61><5>  ( .D(n6968), .CLK(clk), .Q(\mem<61><5> ) );
  DFFPOSX1 \mem_reg<61><4>  ( .D(n6969), .CLK(clk), .Q(\mem<61><4> ) );
  DFFPOSX1 \mem_reg<61><3>  ( .D(n6970), .CLK(clk), .Q(\mem<61><3> ) );
  DFFPOSX1 \mem_reg<61><2>  ( .D(n6971), .CLK(clk), .Q(\mem<61><2> ) );
  DFFPOSX1 \mem_reg<61><1>  ( .D(n6972), .CLK(clk), .Q(\mem<61><1> ) );
  DFFPOSX1 \mem_reg<61><0>  ( .D(n6973), .CLK(clk), .Q(\mem<61><0> ) );
  DFFPOSX1 \mem_reg<62><7>  ( .D(n6974), .CLK(clk), .Q(\mem<62><7> ) );
  DFFPOSX1 \mem_reg<62><6>  ( .D(n6975), .CLK(clk), .Q(\mem<62><6> ) );
  DFFPOSX1 \mem_reg<62><5>  ( .D(n6976), .CLK(clk), .Q(\mem<62><5> ) );
  DFFPOSX1 \mem_reg<62><4>  ( .D(n6977), .CLK(clk), .Q(\mem<62><4> ) );
  DFFPOSX1 \mem_reg<62><3>  ( .D(n6978), .CLK(clk), .Q(\mem<62><3> ) );
  DFFPOSX1 \mem_reg<62><2>  ( .D(n6979), .CLK(clk), .Q(\mem<62><2> ) );
  DFFPOSX1 \mem_reg<62><1>  ( .D(n6980), .CLK(clk), .Q(\mem<62><1> ) );
  DFFPOSX1 \mem_reg<62><0>  ( .D(n6981), .CLK(clk), .Q(\mem<62><0> ) );
  DFFPOSX1 \mem_reg<63><7>  ( .D(n6982), .CLK(clk), .Q(\mem<63><7> ) );
  DFFPOSX1 \mem_reg<63><6>  ( .D(n6983), .CLK(clk), .Q(\mem<63><6> ) );
  DFFPOSX1 \mem_reg<63><5>  ( .D(n6984), .CLK(clk), .Q(\mem<63><5> ) );
  DFFPOSX1 \mem_reg<63><4>  ( .D(n6985), .CLK(clk), .Q(\mem<63><4> ) );
  DFFPOSX1 \mem_reg<63><3>  ( .D(n6986), .CLK(clk), .Q(\mem<63><3> ) );
  DFFPOSX1 \mem_reg<63><2>  ( .D(n6987), .CLK(clk), .Q(\mem<63><2> ) );
  DFFPOSX1 \mem_reg<63><1>  ( .D(n6988), .CLK(clk), .Q(\mem<63><1> ) );
  DFFPOSX1 \mem_reg<63><0>  ( .D(n6989), .CLK(clk), .Q(\mem<63><0> ) );
  INVX2 U3 ( .A(N177), .Y(n1) );
  AND2X2 U4 ( .A(n1), .B(n5216), .Y(n2) );
  AND2X2 U5 ( .A(n3928), .B(n3), .Y(n1541) );
  AND2X2 U6 ( .A(n4949), .B(n92), .Y(n3) );
  AND2X2 U7 ( .A(n92), .B(\data_in<1> ), .Y(n4) );
  MUX2X1 U8 ( .B(n6461), .A(n6462), .S(n3911), .Y(n6485) );
  AND2X2 U9 ( .A(n92), .B(n672), .Y(n5) );
  AND2X2 U10 ( .A(n5750), .B(n4949), .Y(n6) );
  INVX2 U11 ( .A(n4948), .Y(n4949) );
  INVX1 U12 ( .A(n27), .Y(n7) );
  AND2X2 U13 ( .A(n130), .B(n837), .Y(n8) );
  AND2X2 U14 ( .A(n812), .B(n5119), .Y(n9) );
  AND2X2 U15 ( .A(n227), .B(n896), .Y(n10) );
  AND2X2 U16 ( .A(n220), .B(n896), .Y(n11) );
  AND2X2 U17 ( .A(n5140), .B(n765), .Y(n12) );
  AND2X2 U18 ( .A(n131), .B(n740), .Y(n13) );
  AND2X2 U19 ( .A(n5735), .B(n713), .Y(n14) );
  INVX1 U20 ( .A(n6427), .Y(n15) );
  INVX1 U21 ( .A(n409), .Y(n16) );
  AND2X2 U22 ( .A(n217), .B(n873), .Y(n17) );
  AND2X2 U23 ( .A(n224), .B(n873), .Y(n18) );
  AND2X2 U24 ( .A(n5726), .B(n6457), .Y(n19) );
  AND2X2 U25 ( .A(n3681), .B(n6457), .Y(n20) );
  INVX1 U26 ( .A(n5687), .Y(n3934) );
  INVX1 U27 ( .A(n168), .Y(n5186) );
  INVX2 U28 ( .A(n564), .Y(n5181) );
  INVX2 U29 ( .A(n879), .Y(n880) );
  AND2X2 U30 ( .A(n4940), .B(n833), .Y(n21) );
  INVX1 U31 ( .A(n102), .Y(n22) );
  INVX2 U32 ( .A(n5076), .Y(n6426) );
  INVX1 U33 ( .A(n3960), .Y(n3957) );
  INVX1 U34 ( .A(n408), .Y(n23) );
  AND2X2 U35 ( .A(n3678), .B(n6457), .Y(n24) );
  INVX4 U36 ( .A(n5716), .Y(n6457) );
  INVX2 U37 ( .A(n3947), .Y(n5179) );
  INVX2 U38 ( .A(n3965), .Y(n3992) );
  INVX1 U39 ( .A(n31), .Y(n25) );
  INVX1 U40 ( .A(N180), .Y(n5759) );
  INVX1 U41 ( .A(n5713), .Y(n26) );
  INVX1 U42 ( .A(n5713), .Y(n27) );
  INVX1 U43 ( .A(n3656), .Y(n28) );
  INVX1 U44 ( .A(n557), .Y(n29) );
  INVX1 U45 ( .A(n56), .Y(n30) );
  INVX1 U46 ( .A(n5180), .Y(n31) );
  INVX1 U47 ( .A(n31), .Y(n32) );
  INVX1 U48 ( .A(N179), .Y(n5180) );
  INVX4 U49 ( .A(n564), .Y(n33) );
  INVX1 U50 ( .A(n564), .Y(n6459) );
  OR2X1 U51 ( .A(n1694), .B(n473), .Y(n472) );
  INVX1 U52 ( .A(n5758), .Y(n5757) );
  INVX2 U53 ( .A(n5653), .Y(n5209) );
  INVX2 U54 ( .A(n5655), .Y(n5217) );
  INVX2 U55 ( .A(n5650), .Y(n5657) );
  INVX2 U56 ( .A(N178), .Y(n5704) );
  INVX8 U57 ( .A(n5704), .Y(n5673) );
  INVX4 U58 ( .A(n5091), .Y(n3948) );
  INVX2 U59 ( .A(n872), .Y(n5052) );
  INVX2 U60 ( .A(n826), .Y(n827) );
  OR2X2 U61 ( .A(n3916), .B(n171), .Y(n34) );
  INVX4 U62 ( .A(n4963), .Y(n4964) );
  INVX2 U63 ( .A(n765), .Y(n5009) );
  INVX2 U64 ( .A(n5190), .Y(n3989) );
  INVX1 U65 ( .A(\mem<11><5> ), .Y(n5169) );
  INVX1 U66 ( .A(n104), .Y(n79) );
  INVX1 U67 ( .A(\mem<21><4> ), .Y(n6125) );
  INVX1 U68 ( .A(\mem<49><4> ), .Y(n6133) );
  INVX1 U69 ( .A(\mem<33><4> ), .Y(n6116) );
  INVX1 U70 ( .A(\mem<37><4> ), .Y(n6117) );
  INVX1 U71 ( .A(\mem<40><4> ), .Y(n6120) );
  INVX1 U72 ( .A(\mem<58><0> ), .Y(n5779) );
  INVX1 U73 ( .A(\mem<9><1> ), .Y(n5874) );
  INVX1 U74 ( .A(\mem<53><1> ), .Y(n5906) );
  INVX1 U75 ( .A(\mem<1><4> ), .Y(n6150) );
  INVX1 U76 ( .A(\mem<1><0> ), .Y(n5838) );
  INVX1 U77 ( .A(\mem<1><6> ), .Y(n6302) );
  INVX1 U78 ( .A(\mem<9><3> ), .Y(n6031) );
  INVX1 U79 ( .A(\mem<13><3> ), .Y(n6032) );
  INVX1 U80 ( .A(\mem<16><3> ), .Y(n6035) );
  INVX1 U81 ( .A(\mem<37><3> ), .Y(n6040) );
  INVX1 U82 ( .A(\mem<33><3> ), .Y(n6039) );
  INVX1 U83 ( .A(\mem<40><3> ), .Y(n6043) );
  INVX1 U84 ( .A(\mem<1><3> ), .Y(n6072) );
  INVX1 U85 ( .A(\mem<46><1> ), .Y(n5928) );
  INVX1 U86 ( .A(\mem<48><1> ), .Y(n5926) );
  INVX1 U87 ( .A(\mem<41><1> ), .Y(n5931) );
  INVX1 U88 ( .A(\mem<32><2> ), .Y(n5946) );
  INVX1 U89 ( .A(\mem<28><2> ), .Y(n5944) );
  INVX1 U90 ( .A(\mem<1><2> ), .Y(n6001) );
  INVX1 U91 ( .A(\mem<12><5> ), .Y(n6174) );
  INVX1 U92 ( .A(\mem<13><5> ), .Y(n6178) );
  INVX1 U93 ( .A(\mem<16><5> ), .Y(n6181) );
  INVX1 U94 ( .A(\mem<17><5> ), .Y(n6198) );
  INVX1 U95 ( .A(\mem<1><7> ), .Y(n6382) );
  AND2X1 U96 ( .A(n5427), .B(n5196), .Y(n4145) );
  INVX1 U97 ( .A(\mem<1><5> ), .Y(n6223) );
  INVX1 U98 ( .A(\mem<5><5> ), .Y(n6225) );
  INVX1 U99 ( .A(\mem<6><5> ), .Y(n6220) );
  INVX1 U100 ( .A(\mem<16><4> ), .Y(n6109) );
  INVX1 U101 ( .A(\mem<13><4> ), .Y(n6106) );
  INVX1 U102 ( .A(\mem<9><4> ), .Y(n6105) );
  INVX1 U103 ( .A(\mem<35><3> ), .Y(n3916) );
  INVX1 U104 ( .A(\mem<28><4> ), .Y(n6096) );
  INVX1 U105 ( .A(\mem<32><4> ), .Y(n6098) );
  INVX1 U106 ( .A(\mem<20><4> ), .Y(n6122) );
  INVX1 U107 ( .A(\mem<17><4> ), .Y(n6124) );
  INVX1 U108 ( .A(\mem<18><4> ), .Y(n207) );
  INVX1 U109 ( .A(\mem<24><4> ), .Y(n6128) );
  INVX1 U110 ( .A(\mem<53><4> ), .Y(n6134) );
  INVX1 U111 ( .A(\mem<56><4> ), .Y(n6137) );
  INVX1 U112 ( .A(\mem<52><4> ), .Y(n6130) );
  INVX1 U113 ( .A(\mem<36><4> ), .Y(n6113) );
  INVX1 U114 ( .A(\mem<12><4> ), .Y(n6103) );
  INVX1 U115 ( .A(\mem<34><4> ), .Y(n214) );
  INVX1 U116 ( .A(\mem<33><0> ), .Y(n5799) );
  INVX1 U117 ( .A(\mem<40><0> ), .Y(n5803) );
  INVX1 U118 ( .A(\mem<37><0> ), .Y(n5800) );
  INVX1 U119 ( .A(\mem<9><0> ), .Y(n5788) );
  INVX1 U120 ( .A(\mem<16><0> ), .Y(n5792) );
  INVX1 U121 ( .A(\mem<13><0> ), .Y(n5789) );
  INVX1 U122 ( .A(\mem<24><0> ), .Y(n5814) );
  INVX1 U123 ( .A(\mem<17><0> ), .Y(n5810) );
  INVX1 U124 ( .A(\mem<21><0> ), .Y(n5811) );
  INVX1 U125 ( .A(\mem<56><0> ), .Y(n5825) );
  INVX1 U126 ( .A(\mem<53><0> ), .Y(n5822) );
  INVX1 U127 ( .A(\mem<49><0> ), .Y(n5821) );
  INVX1 U128 ( .A(\mem<32><0> ), .Y(n5767) );
  INVX1 U129 ( .A(\mem<28><0> ), .Y(n5764) );
  INVX1 U130 ( .A(\mem<59><0> ), .Y(n5782) );
  INVX1 U131 ( .A(\mem<62><0> ), .Y(n5777) );
  INVX1 U132 ( .A(\mem<24><6> ), .Y(n6278) );
  INVX1 U133 ( .A(\mem<21><6> ), .Y(n6275) );
  INVX1 U134 ( .A(\mem<17><6> ), .Y(n6274) );
  INVX1 U135 ( .A(\mem<53><6> ), .Y(n6286) );
  INVX1 U136 ( .A(\mem<56><6> ), .Y(n6289) );
  INVX1 U137 ( .A(\mem<49><6> ), .Y(n6285) );
  INVX1 U138 ( .A(\mem<16><6> ), .Y(n6259) );
  INVX1 U139 ( .A(\mem<9><6> ), .Y(n6255) );
  INVX1 U140 ( .A(\mem<13><6> ), .Y(n6256) );
  INVX1 U141 ( .A(\mem<40><6> ), .Y(n6269) );
  INVX1 U142 ( .A(\mem<37><6> ), .Y(n6266) );
  INVX1 U143 ( .A(\mem<33><6> ), .Y(n6265) );
  INVX1 U144 ( .A(\mem<32><6> ), .Y(n6249) );
  INVX1 U145 ( .A(\mem<28><6> ), .Y(n6247) );
  INVX1 U146 ( .A(\mem<40><1> ), .Y(n5888) );
  INVX1 U147 ( .A(\mem<33><1> ), .Y(n5884) );
  INVX1 U148 ( .A(\mem<37><1> ), .Y(n5885) );
  INVX1 U149 ( .A(\mem<12><1> ), .Y(n5871) );
  INVX1 U150 ( .A(\mem<16><1> ), .Y(n5878) );
  INVX1 U151 ( .A(\mem<13><1> ), .Y(n5875) );
  INVX1 U152 ( .A(\mem<21><1> ), .Y(n5896) );
  INVX1 U153 ( .A(\mem<24><1> ), .Y(n5899) );
  INVX1 U154 ( .A(\mem<17><1> ), .Y(n5895) );
  INVX1 U155 ( .A(\mem<56><1> ), .Y(n5909) );
  INVX1 U156 ( .A(\mem<49><1> ), .Y(n5905) );
  INVX1 U157 ( .A(\mem<45><1> ), .Y(n5932) );
  INVX1 U158 ( .A(\mem<21><3> ), .Y(n6049) );
  INVX1 U159 ( .A(\mem<24><3> ), .Y(n6052) );
  INVX1 U160 ( .A(\mem<17><3> ), .Y(n6048) );
  INVX1 U161 ( .A(\mem<53><3> ), .Y(n6060) );
  INVX1 U162 ( .A(\mem<56><3> ), .Y(n6063) );
  INVX1 U163 ( .A(\mem<49><3> ), .Y(n6059) );
  INVX1 U164 ( .A(\mem<45><4> ), .Y(n6160) );
  INVX1 U165 ( .A(\mem<41><4> ), .Y(n6159) );
  INVX1 U166 ( .A(\mem<48><4> ), .Y(n6154) );
  INVX1 U167 ( .A(\mem<46><4> ), .Y(n6156) );
  INVX1 U168 ( .A(\mem<8><4> ), .Y(n6144) );
  INVX1 U169 ( .A(\mem<6><4> ), .Y(n6146) );
  INVX1 U170 ( .A(\mem<5><4> ), .Y(n6151) );
  INVX1 U171 ( .A(\mem<9><5> ), .Y(n6177) );
  INVX1 U172 ( .A(n97), .Y(n5277) );
  INVX1 U173 ( .A(\mem<63><1> ), .Y(n99) );
  INVX1 U174 ( .A(\mem<62><1> ), .Y(n98) );
  INVX1 U175 ( .A(\mem<41><0> ), .Y(n5851) );
  INVX1 U176 ( .A(\mem<45><0> ), .Y(n5853) );
  INVX1 U177 ( .A(\mem<48><0> ), .Y(n5845) );
  INVX1 U178 ( .A(\mem<46><0> ), .Y(n5847) );
  INVX1 U179 ( .A(\mem<8><0> ), .Y(n5833) );
  INVX1 U180 ( .A(\mem<6><0> ), .Y(n5834) );
  INVX1 U181 ( .A(\mem<5><0> ), .Y(n5840) );
  INVX1 U182 ( .A(\mem<36><0> ), .Y(n5796) );
  INVX1 U183 ( .A(\mem<12><0> ), .Y(n5786) );
  INVX1 U184 ( .A(\mem<52><0> ), .Y(n5818) );
  INVX1 U185 ( .A(\mem<20><0> ), .Y(n5808) );
  INVX1 U186 ( .A(\mem<41><6> ), .Y(n6313) );
  INVX1 U187 ( .A(\mem<45><6> ), .Y(n6315) );
  INVX1 U188 ( .A(\mem<48><6> ), .Y(n6307) );
  INVX1 U189 ( .A(\mem<46><6> ), .Y(n6309) );
  INVX1 U190 ( .A(\mem<8><6> ), .Y(n6296) );
  INVX1 U191 ( .A(\mem<6><6> ), .Y(n6298) );
  INVX1 U192 ( .A(\mem<5><6> ), .Y(n6304) );
  INVX1 U193 ( .A(\mem<52><6> ), .Y(n6282) );
  INVX1 U194 ( .A(\mem<36><6> ), .Y(n6263) );
  INVX1 U195 ( .A(\mem<12><6> ), .Y(n6253) );
  INVX1 U196 ( .A(\mem<36><1> ), .Y(n5882) );
  INVX1 U197 ( .A(\mem<20><1> ), .Y(n5892) );
  INVX1 U198 ( .A(\mem<32><1> ), .Y(n5866) );
  INVX1 U199 ( .A(\mem<28><1> ), .Y(n5864) );
  INVX1 U200 ( .A(\mem<8><1> ), .Y(n5915) );
  INVX1 U201 ( .A(\mem<6><1> ), .Y(n5917) );
  INVX1 U202 ( .A(\mem<5><1> ), .Y(n5923) );
  INVX1 U203 ( .A(\mem<13><2> ), .Y(n5955) );
  INVX1 U204 ( .A(\mem<16><2> ), .Y(n5958) );
  INVX1 U205 ( .A(\mem<9><2> ), .Y(n5953) );
  INVX1 U206 ( .A(\mem<40><2> ), .Y(n5968) );
  INVX1 U207 ( .A(\mem<33><2> ), .Y(n5964) );
  INVX1 U208 ( .A(\mem<37><2> ), .Y(n5965) );
  INVX1 U209 ( .A(\mem<21><2> ), .Y(n5975) );
  INVX1 U210 ( .A(\mem<24><2> ), .Y(n5978) );
  INVX1 U211 ( .A(\mem<17><2> ), .Y(n5974) );
  INVX1 U212 ( .A(\mem<56><2> ), .Y(n5989) );
  INVX1 U213 ( .A(\mem<53><2> ), .Y(n5986) );
  INVX1 U214 ( .A(\mem<49><2> ), .Y(n5985) );
  INVX1 U215 ( .A(\mem<10><3> ), .Y(n84) );
  INVX1 U216 ( .A(\mem<12><3> ), .Y(n6028) );
  INVX1 U217 ( .A(\mem<34><3> ), .Y(n405) );
  INVX1 U218 ( .A(\mem<36><3> ), .Y(n6037) );
  INVX1 U219 ( .A(\mem<20><3> ), .Y(n6045) );
  INVX1 U220 ( .A(\mem<52><3> ), .Y(n6056) );
  INVX1 U221 ( .A(\mem<32><3> ), .Y(n6023) );
  INVX1 U222 ( .A(\mem<28><3> ), .Y(n6021) );
  INVX1 U223 ( .A(\mem<45><3> ), .Y(n6084) );
  INVX1 U224 ( .A(\mem<46><3> ), .Y(n6079) );
  INVX1 U225 ( .A(\mem<48><3> ), .Y(n6077) );
  INVX1 U226 ( .A(\mem<8><3> ), .Y(n6069) );
  INVX1 U227 ( .A(\mem<5><3> ), .Y(n6074) );
  INVX1 U228 ( .A(\mem<40><5> ), .Y(n6192) );
  INVX1 U229 ( .A(\mem<33><5> ), .Y(n6188) );
  INVX1 U230 ( .A(\mem<37><5> ), .Y(n6189) );
  INVX1 U231 ( .A(\mem<24><5> ), .Y(n6202) );
  INVX1 U232 ( .A(\mem<20><5> ), .Y(n6196) );
  INVX1 U233 ( .A(\mem<56><5> ), .Y(n6212) );
  INVX1 U234 ( .A(\mem<49><5> ), .Y(n6208) );
  INVX1 U235 ( .A(\mem<53><5> ), .Y(n6209) );
  INVX1 U236 ( .A(\mem<8><5> ), .Y(n6218) );
  INVX1 U237 ( .A(\mem<17><7> ), .Y(n6354) );
  INVX1 U238 ( .A(\mem<24><7> ), .Y(n6358) );
  INVX1 U239 ( .A(\mem<21><7> ), .Y(n6355) );
  INVX1 U240 ( .A(\mem<53><7> ), .Y(n6366) );
  INVX1 U241 ( .A(\mem<56><7> ), .Y(n6369) );
  INVX1 U242 ( .A(\mem<49><7> ), .Y(n6365) );
  INVX1 U243 ( .A(\mem<16><7> ), .Y(n6338) );
  INVX1 U244 ( .A(\mem<9><7> ), .Y(n6334) );
  INVX1 U245 ( .A(\mem<13><7> ), .Y(n6335) );
  INVX1 U246 ( .A(\mem<33><7> ), .Y(n6344) );
  INVX1 U247 ( .A(\mem<40><7> ), .Y(n6348) );
  INVX1 U248 ( .A(\mem<37><7> ), .Y(n6345) );
  INVX1 U249 ( .A(\mem<32><7> ), .Y(n6328) );
  INVX1 U250 ( .A(\mem<28><7> ), .Y(n6326) );
  INVX1 U251 ( .A(\mem<58><3> ), .Y(n5197) );
  INVX1 U252 ( .A(n5667), .Y(n94) );
  INVX1 U253 ( .A(n5667), .Y(n3969) );
  AND2X1 U254 ( .A(n1122), .B(n1099), .Y(n637) );
  INVX1 U255 ( .A(\mem<36><2> ), .Y(n5962) );
  INVX1 U256 ( .A(\mem<12><2> ), .Y(n5951) );
  INVX1 U257 ( .A(\mem<52><2> ), .Y(n5982) );
  INVX1 U258 ( .A(\mem<20><2> ), .Y(n5972) );
  AND2X1 U259 ( .A(n639), .B(n640), .Y(n916) );
  INVX1 U260 ( .A(\mem<41><2> ), .Y(n6012) );
  INVX1 U261 ( .A(\mem<45><2> ), .Y(n6013) );
  INVX1 U262 ( .A(\mem<48><2> ), .Y(n6006) );
  INVX1 U263 ( .A(\mem<46><2> ), .Y(n6008) );
  INVX1 U264 ( .A(\mem<6><2> ), .Y(n5997) );
  INVX1 U265 ( .A(\mem<8><2> ), .Y(n5996) );
  INVX1 U266 ( .A(\mem<5><2> ), .Y(n6003) );
  AND2X1 U267 ( .A(n935), .B(n496), .Y(n1675) );
  INVX1 U268 ( .A(\mem<36><5> ), .Y(n6185) );
  INVX1 U269 ( .A(n27), .Y(n204) );
  INVX1 U270 ( .A(\mem<21><5> ), .Y(n6199) );
  INVX1 U271 ( .A(\mem<52><5> ), .Y(n6206) );
  INVX1 U272 ( .A(\mem<32><5> ), .Y(n6169) );
  INVX1 U273 ( .A(\mem<28><5> ), .Y(n6167) );
  INVX1 U274 ( .A(\mem<41><5> ), .Y(n6234) );
  INVX1 U275 ( .A(\mem<45><5> ), .Y(n6235) );
  INVX1 U276 ( .A(\mem<48><5> ), .Y(n6228) );
  INVX1 U277 ( .A(\mem<46><5> ), .Y(n6230) );
  INVX1 U278 ( .A(\mem<41><7> ), .Y(n6392) );
  INVX1 U279 ( .A(\mem<45><7> ), .Y(n6394) );
  INVX1 U280 ( .A(\mem<48><7> ), .Y(n6386) );
  INVX1 U281 ( .A(\mem<46><7> ), .Y(n6388) );
  INVX1 U282 ( .A(\mem<8><7> ), .Y(n6376) );
  INVX1 U283 ( .A(\mem<6><7> ), .Y(n6378) );
  INVX1 U284 ( .A(\mem<5><7> ), .Y(n6383) );
  INVX1 U285 ( .A(\mem<52><7> ), .Y(n6362) );
  INVX1 U286 ( .A(\mem<20><7> ), .Y(n6352) );
  INVX1 U287 ( .A(\mem<36><7> ), .Y(n6342) );
  INVX1 U288 ( .A(\mem<12><7> ), .Y(n6332) );
  INVX1 U289 ( .A(n5670), .Y(n5158) );
  INVX1 U290 ( .A(n5669), .Y(n3974) );
  INVX1 U291 ( .A(rst), .Y(n5760) );
  AND2X1 U292 ( .A(n5439), .B(n3948), .Y(n3739) );
  AND2X1 U293 ( .A(n937), .B(n966), .Y(n1687) );
  AND2X1 U294 ( .A(n5379), .B(n3917), .Y(n3723) );
  AND2X1 U295 ( .A(n5631), .B(n5185), .Y(n4133) );
  INVX1 U296 ( .A(\data_in<8> ), .Y(n6461) );
  INVX1 U297 ( .A(\mem<0><0> ), .Y(n6462) );
  INVX1 U298 ( .A(\data_in<9> ), .Y(n6463) );
  INVX1 U299 ( .A(\mem<0><1> ), .Y(n6464) );
  INVX1 U300 ( .A(\data_in<10> ), .Y(n6465) );
  INVX1 U301 ( .A(\mem<0><2> ), .Y(n6466) );
  INVX1 U302 ( .A(\data_in<11> ), .Y(n6467) );
  INVX1 U303 ( .A(\mem<0><3> ), .Y(n6468) );
  INVX1 U304 ( .A(\data_in<12> ), .Y(n6469) );
  INVX1 U305 ( .A(\mem<0><4> ), .Y(n6470) );
  INVX1 U306 ( .A(\data_in<13> ), .Y(n6471) );
  INVX1 U307 ( .A(\mem<0><5> ), .Y(n6472) );
  INVX1 U308 ( .A(\data_in<14> ), .Y(n6473) );
  INVX1 U309 ( .A(\mem<0><6> ), .Y(n6474) );
  INVX1 U310 ( .A(\data_in<15> ), .Y(n6475) );
  INVX1 U311 ( .A(\mem<0><7> ), .Y(n6476) );
  INVX1 U312 ( .A(n5187), .Y(n5742) );
  INVX8 U313 ( .A(n5648), .Y(n5649) );
  INVX8 U314 ( .A(n81), .Y(n5686) );
  INVX1 U315 ( .A(n5649), .Y(n72) );
  AND2X1 U316 ( .A(n6173), .B(n4112), .Y(n596) );
  INVX1 U317 ( .A(n5649), .Y(n71) );
  AND2X2 U318 ( .A(\mem<57><1> ), .B(n5753), .Y(n35) );
  AND2X2 U319 ( .A(\mem<57><3> ), .B(n5753), .Y(n36) );
  AND2X2 U320 ( .A(\mem<57><5> ), .B(n5753), .Y(n37) );
  INVX4 U321 ( .A(n88), .Y(n5750) );
  AND2X2 U322 ( .A(\mem<59><1> ), .B(n185), .Y(n38) );
  AND2X2 U323 ( .A(\mem<59><3> ), .B(n184), .Y(n39) );
  AND2X2 U324 ( .A(\mem<59><5> ), .B(n190), .Y(n40) );
  AND2X2 U325 ( .A(\mem<62><3> ), .B(n5732), .Y(n41) );
  AND2X2 U326 ( .A(\mem<62><5> ), .B(n5732), .Y(n42) );
  INVX1 U327 ( .A(\mem<41><3> ), .Y(n6083) );
  INVX2 U328 ( .A(n5738), .Y(n5736) );
  MUX2X1 U329 ( .B(n6473), .A(n6474), .S(n3911), .Y(n6479) );
  AND2X2 U330 ( .A(n678), .B(n133), .Y(n43) );
  AND2X2 U331 ( .A(n161), .B(n837), .Y(n44) );
  INVX1 U332 ( .A(n46), .Y(n45) );
  INVX1 U333 ( .A(n5713), .Y(n46) );
  INVX2 U334 ( .A(n904), .Y(n47) );
  AND2X2 U335 ( .A(n812), .B(n5120), .Y(n48) );
  AND2X2 U336 ( .A(n5728), .B(n783), .Y(n49) );
  INVX1 U337 ( .A(n63), .Y(n50) );
  AND2X2 U338 ( .A(n162), .B(n740), .Y(n51) );
  AND2X2 U339 ( .A(n5732), .B(n713), .Y(n52) );
  INVX4 U340 ( .A(n5733), .Y(n5732) );
  AND2X2 U341 ( .A(n223), .B(n696), .Y(n53) );
  INVX2 U342 ( .A(n3684), .Y(n223) );
  INVX1 U343 ( .A(n3656), .Y(n54) );
  INVX1 U344 ( .A(n3656), .Y(n61) );
  INVX1 U345 ( .A(n5708), .Y(n55) );
  INVX1 U346 ( .A(n6429), .Y(n56) );
  INVX1 U347 ( .A(n869), .Y(n57) );
  INVX1 U348 ( .A(n6400), .Y(n58) );
  INVX1 U349 ( .A(n6400), .Y(n59) );
  INVX1 U350 ( .A(n691), .Y(n60) );
  INVX1 U351 ( .A(n3656), .Y(n68) );
  INVX1 U352 ( .A(n26), .Y(n62) );
  INVX1 U353 ( .A(n903), .Y(n63) );
  MUX2X1 U354 ( .B(n5500), .A(n5499), .S(n5659), .Y(n5498) );
  AND2X2 U355 ( .A(n5121), .B(n765), .Y(n64) );
  MUX2X1 U356 ( .B(n5567), .A(n5570), .S(n5209), .Y(n5581) );
  MUX2X1 U357 ( .B(n5446), .A(n5445), .S(n5659), .Y(n5444) );
  INVX1 U358 ( .A(n5807), .Y(n65) );
  INVX1 U359 ( .A(n16), .Y(n66) );
  INVX1 U360 ( .A(n876), .Y(n67) );
  MUX2X1 U361 ( .B(n5611), .A(n5610), .S(n5658), .Y(n5609) );
  MUX2X1 U362 ( .B(n523), .A(n600), .S(n5649), .Y(n5246) );
  INVX2 U363 ( .A(n3656), .Y(n3657) );
  MUX2X1 U364 ( .B(n498), .A(n5523), .S(n5649), .Y(n5522) );
  INVX2 U365 ( .A(n5649), .Y(n5212) );
  MUX2X1 U366 ( .B(n603), .A(n5440), .S(n5648), .Y(n5439) );
  INVX1 U367 ( .A(n5156), .Y(n6424) );
  INVX1 U368 ( .A(n897), .Y(n69) );
  INVX1 U369 ( .A(n4939), .Y(n70) );
  MUX2X1 U370 ( .B(n588), .A(n519), .S(n5150), .Y(N185) );
  MUX2X1 U371 ( .B(n583), .A(n612), .S(n71), .Y(n5593) );
  MUX2X1 U372 ( .B(n601), .A(n5274), .S(n72), .Y(n5273) );
  INVX1 U373 ( .A(n5205), .Y(n73) );
  MUX2X1 U374 ( .B(n528), .A(n5353), .S(n5212), .Y(n5352) );
  INVX1 U375 ( .A(n833), .Y(n74) );
  MUX2X1 U376 ( .B(\mem<15><3> ), .A(\mem<14><3> ), .S(n5678), .Y(n5414) );
  INVX1 U377 ( .A(n694), .Y(n75) );
  INVX4 U378 ( .A(n5697), .Y(n5688) );
  MUX2X1 U379 ( .B(n5400), .A(n5399), .S(n5660), .Y(n5398) );
  INVX8 U380 ( .A(n5678), .Y(n5694) );
  INVX2 U381 ( .A(n22), .Y(n76) );
  INVX1 U382 ( .A(n6427), .Y(n5708) );
  INVX1 U383 ( .A(n102), .Y(n6427) );
  INVX2 U384 ( .A(n5113), .Y(n78) );
  MUX2X1 U385 ( .B(n608), .A(n5385), .S(n5660), .Y(n5384) );
  INVX4 U386 ( .A(n616), .Y(n77) );
  INVX2 U387 ( .A(n616), .Y(n205) );
  INVX2 U388 ( .A(n5698), .Y(n5675) );
  INVX1 U389 ( .A(n5160), .Y(n3959) );
  INVX1 U390 ( .A(n408), .Y(n80) );
  INVX1 U391 ( .A(n5220), .Y(n5151) );
  INVX1 U392 ( .A(n80), .Y(n6439) );
  INVX2 U393 ( .A(n3965), .Y(n81) );
  INVX1 U394 ( .A(n5145), .Y(n82) );
  INVX2 U395 ( .A(n5718), .Y(n92) );
  OAI21X1 U396 ( .A(n84), .B(n5119), .C(n85), .Y(n83) );
  OR2X2 U397 ( .A(n5723), .B(n6035), .Y(n85) );
  INVX1 U398 ( .A(n3660), .Y(n86) );
  INVX4 U399 ( .A(n3658), .Y(n3660) );
  INVX2 U400 ( .A(n5754), .Y(n87) );
  INVX1 U401 ( .A(n5754), .Y(n88) );
  INVX1 U402 ( .A(n5754), .Y(n5752) );
  AND2X2 U403 ( .A(n5219), .B(\mem<52><1> ), .Y(n5903) );
  INVX1 U404 ( .A(n5719), .Y(n103) );
  MUX2X1 U405 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n93), .Y(n5320) );
  INVX1 U406 ( .A(n1), .Y(n89) );
  NOR3X1 U407 ( .A(n1152), .B(\addr<7> ), .C(n3034), .Y(n90) );
  INVX1 U408 ( .A(n3991), .Y(n91) );
  INVX1 U409 ( .A(n3940), .Y(n93) );
  MUX2X1 U410 ( .B(n5417), .A(n5416), .S(n94), .Y(n5415) );
  INVX1 U411 ( .A(n103), .Y(n95) );
  BUFX2 U412 ( .A(n29), .Y(n96) );
  MUX2X1 U413 ( .B(n99), .A(n98), .S(n5679), .Y(n97) );
  INVX1 U414 ( .A(n5157), .Y(n100) );
  INVX1 U415 ( .A(n5752), .Y(n101) );
  MUX2X1 U416 ( .B(n610), .A(n5425), .S(n5648), .Y(n5424) );
  INVX2 U417 ( .A(N180), .Y(n5648) );
  NOR3X1 U418 ( .A(n3926), .B(n4221), .C(n5082), .Y(n102) );
  INVX1 U419 ( .A(n205), .Y(n104) );
  INVX1 U420 ( .A(n104), .Y(n105) );
  INVX1 U421 ( .A(n5677), .Y(n106) );
  INVX4 U422 ( .A(n3993), .Y(n5677) );
  INVX1 U423 ( .A(N177), .Y(n107) );
  INVX1 U424 ( .A(n517), .Y(n108) );
  AND2X2 U425 ( .A(n168), .B(n623), .Y(n109) );
  INVX1 U426 ( .A(n5746), .Y(n110) );
  INVX1 U427 ( .A(n5746), .Y(n111) );
  INVX1 U428 ( .A(n110), .Y(n112) );
  INVX1 U429 ( .A(n110), .Y(n113) );
  INVX1 U430 ( .A(n111), .Y(n114) );
  INVX1 U431 ( .A(n111), .Y(n115) );
  INVX1 U432 ( .A(n3943), .Y(n116) );
  INVX1 U433 ( .A(n116), .Y(n117) );
  INVX1 U434 ( .A(n116), .Y(n118) );
  INVX1 U435 ( .A(n156), .Y(n119) );
  INVX1 U436 ( .A(n116), .Y(n120) );
  INVX1 U437 ( .A(n5745), .Y(n121) );
  INVX1 U438 ( .A(n5745), .Y(n122) );
  INVX1 U439 ( .A(n121), .Y(n123) );
  INVX1 U440 ( .A(n121), .Y(n124) );
  INVX1 U441 ( .A(n122), .Y(n125) );
  INVX1 U442 ( .A(n122), .Y(n126) );
  INVX1 U443 ( .A(n5743), .Y(n127) );
  INVX1 U444 ( .A(n3944), .Y(n128) );
  INVX1 U445 ( .A(n122), .Y(n129) );
  INVX1 U446 ( .A(n127), .Y(n130) );
  INVX1 U447 ( .A(n127), .Y(n131) );
  INVX1 U448 ( .A(n148), .Y(n132) );
  INVX1 U449 ( .A(n150), .Y(n133) );
  INVX1 U450 ( .A(n132), .Y(n134) );
  INVX1 U451 ( .A(n132), .Y(n135) );
  INVX1 U452 ( .A(n122), .Y(n136) );
  INVX1 U453 ( .A(n158), .Y(n137) );
  INVX1 U454 ( .A(n158), .Y(n138) );
  INVX1 U455 ( .A(n156), .Y(n139) );
  INVX1 U456 ( .A(n5744), .Y(n140) );
  INVX1 U457 ( .A(n160), .Y(n141) );
  INVX1 U458 ( .A(n140), .Y(n142) );
  INVX1 U459 ( .A(n140), .Y(n143) );
  INVX1 U460 ( .A(n109), .Y(n144) );
  INVX1 U461 ( .A(n109), .Y(n145) );
  INVX1 U462 ( .A(n109), .Y(n146) );
  INVX1 U463 ( .A(n109), .Y(n147) );
  INVX1 U464 ( .A(n109), .Y(n148) );
  INVX1 U465 ( .A(n144), .Y(n149) );
  INVX1 U466 ( .A(n144), .Y(n150) );
  INVX1 U467 ( .A(n145), .Y(n151) );
  INVX1 U468 ( .A(n145), .Y(n152) );
  INVX1 U469 ( .A(n146), .Y(n153) );
  INVX1 U470 ( .A(n146), .Y(n154) );
  INVX1 U471 ( .A(n147), .Y(n155) );
  INVX1 U472 ( .A(n147), .Y(n156) );
  INVX1 U473 ( .A(n148), .Y(n157) );
  INVX1 U474 ( .A(n148), .Y(n158) );
  INVX1 U475 ( .A(n5219), .Y(n159) );
  INVX1 U476 ( .A(n159), .Y(n160) );
  INVX1 U477 ( .A(n159), .Y(n161) );
  INVX1 U478 ( .A(n146), .Y(n162) );
  INVX1 U479 ( .A(n5745), .Y(n163) );
  INVX1 U480 ( .A(n159), .Y(n164) );
  INVX1 U481 ( .A(n3943), .Y(n3944) );
  INVX1 U482 ( .A(n5219), .Y(n5745) );
  INVX1 U483 ( .A(n3944), .Y(n5743) );
  INVX1 U484 ( .A(n155), .Y(n5744) );
  INVX1 U485 ( .A(n3654), .Y(n165) );
  INVX1 U486 ( .A(n165), .Y(n166) );
  INVX1 U487 ( .A(n5679), .Y(n167) );
  INVX2 U488 ( .A(n5755), .Y(n5679) );
  MUX2X1 U489 ( .B(n530), .A(n5312), .S(n5212), .Y(n5311) );
  MUX2X1 U490 ( .B(n526), .A(n5303), .S(n5662), .Y(n5302) );
  INVX2 U491 ( .A(n3658), .Y(n3659) );
  INVX1 U492 ( .A(n3992), .Y(n168) );
  INVX1 U493 ( .A(n6454), .Y(n169) );
  INVX1 U494 ( .A(n6454), .Y(n170) );
  INVX1 U495 ( .A(n169), .Y(n171) );
  INVX1 U496 ( .A(n177), .Y(n172) );
  INVX1 U497 ( .A(n5747), .Y(n173) );
  INVX1 U498 ( .A(n172), .Y(n174) );
  INVX1 U499 ( .A(n173), .Y(n175) );
  INVX1 U500 ( .A(n170), .Y(n176) );
  INVX1 U501 ( .A(n170), .Y(n177) );
  INVX1 U502 ( .A(n5174), .Y(n178) );
  INVX1 U503 ( .A(n5174), .Y(n179) );
  INVX1 U504 ( .A(n2), .Y(n180) );
  INVX1 U505 ( .A(n5174), .Y(n181) );
  INVX1 U506 ( .A(n2), .Y(n182) );
  INVX1 U507 ( .A(n178), .Y(n183) );
  INVX1 U508 ( .A(n178), .Y(n184) );
  INVX1 U509 ( .A(n178), .Y(n185) );
  INVX1 U510 ( .A(n179), .Y(n186) );
  INVX1 U511 ( .A(n179), .Y(n187) );
  INVX1 U512 ( .A(n179), .Y(n188) );
  INVX1 U513 ( .A(n180), .Y(n189) );
  INVX1 U514 ( .A(n181), .Y(n190) );
  INVX1 U515 ( .A(n5747), .Y(n191) );
  INVX1 U516 ( .A(n171), .Y(n192) );
  INVX1 U517 ( .A(n182), .Y(n193) );
  INVX1 U518 ( .A(n180), .Y(n194) );
  INVX1 U519 ( .A(n180), .Y(n195) );
  INVX1 U520 ( .A(n180), .Y(n196) );
  INVX1 U521 ( .A(n181), .Y(n197) );
  INVX1 U522 ( .A(n181), .Y(n198) );
  INVX1 U523 ( .A(n181), .Y(n199) );
  INVX1 U524 ( .A(n182), .Y(n200) );
  INVX1 U525 ( .A(n182), .Y(n201) );
  INVX1 U526 ( .A(n182), .Y(n202) );
  INVX1 U527 ( .A(n182), .Y(n203) );
  INVX1 U528 ( .A(n2), .Y(n6454) );
  INVX1 U529 ( .A(n5125), .Y(n5133) );
  INVX2 U530 ( .A(n5677), .Y(n5690) );
  INVX1 U531 ( .A(n616), .Y(n617) );
  OAI21X1 U532 ( .A(n207), .B(n5119), .C(n208), .Y(n206) );
  OR2X2 U533 ( .A(n5722), .B(n6128), .Y(n208) );
  INVX2 U534 ( .A(n5152), .Y(n3947) );
  INVX1 U535 ( .A(n5713), .Y(n209) );
  INVX1 U536 ( .A(n209), .Y(n210) );
  INVX1 U537 ( .A(n5699), .Y(n211) );
  INVX1 U538 ( .A(n5699), .Y(n5701) );
  INVX1 U539 ( .A(n5123), .Y(n5128) );
  INVX1 U540 ( .A(n5124), .Y(n5129) );
  INVX8 U541 ( .A(n5725), .Y(n5722) );
  INVX1 U542 ( .A(n5133), .Y(n215) );
  INVX1 U543 ( .A(n3994), .Y(n5153) );
  INVX1 U544 ( .A(n497), .Y(n212) );
  INVX1 U545 ( .A(n5154), .Y(n3965) );
  OR2X2 U546 ( .A(n1699), .B(n479), .Y(n478) );
  OAI21X1 U547 ( .A(n214), .B(n215), .C(n216), .Y(n213) );
  OR2X2 U548 ( .A(n5722), .B(n6120), .Y(n216) );
  INVX1 U549 ( .A(n5135), .Y(n5141) );
  INVX4 U550 ( .A(n548), .Y(n549) );
  INVX4 U551 ( .A(n228), .Y(n5678) );
  INVX1 U552 ( .A(n165), .Y(n5138) );
  INVX1 U553 ( .A(N177), .Y(n5154) );
  INVX4 U554 ( .A(n3660), .Y(n5719) );
  INVX8 U555 ( .A(n3660), .Y(n5717) );
  INVX4 U556 ( .A(N181), .Y(n5843) );
  INVX1 U557 ( .A(n33), .Y(n5182) );
  INVX1 U558 ( .A(n78), .Y(n5178) );
  INVX1 U559 ( .A(n3685), .Y(n217) );
  INVX1 U560 ( .A(n3685), .Y(n218) );
  INVX1 U561 ( .A(n5729), .Y(n219) );
  INVX1 U562 ( .A(n5729), .Y(n220) );
  INVX1 U563 ( .A(n5728), .Y(n221) );
  INVX1 U564 ( .A(n5728), .Y(n222) );
  INVX1 U565 ( .A(n3684), .Y(n224) );
  INVX1 U566 ( .A(n3684), .Y(n225) );
  INVX1 U567 ( .A(n3684), .Y(n226) );
  INVX1 U568 ( .A(n3684), .Y(n227) );
  INVX1 U569 ( .A(n1), .Y(n228) );
  INVX1 U570 ( .A(n217), .Y(n5729) );
  INVX1 U571 ( .A(n217), .Y(n5728) );
  INVX1 U572 ( .A(n5152), .Y(n5190) );
  INVX1 U573 ( .A(N177), .Y(n5756) );
  INVX1 U574 ( .A(n4938), .Y(n229) );
  INVX1 U575 ( .A(n4938), .Y(n230) );
  BUFX2 U576 ( .A(n4938), .Y(n231) );
  BUFX2 U577 ( .A(n4938), .Y(n232) );
  BUFX2 U578 ( .A(n4938), .Y(n233) );
  INVX1 U579 ( .A(n231), .Y(n234) );
  INVX1 U580 ( .A(n231), .Y(n235) );
  INVX1 U581 ( .A(n231), .Y(n236) );
  INVX1 U582 ( .A(n231), .Y(n237) );
  INVX1 U583 ( .A(n232), .Y(n238) );
  INVX1 U584 ( .A(n232), .Y(n239) );
  INVX1 U585 ( .A(n232), .Y(n240) );
  INVX1 U586 ( .A(n232), .Y(n241) );
  INVX1 U587 ( .A(n229), .Y(n242) );
  INVX1 U588 ( .A(n229), .Y(n243) );
  INVX1 U589 ( .A(n229), .Y(n244) );
  INVX1 U590 ( .A(n242), .Y(n245) );
  INVX1 U591 ( .A(n242), .Y(n246) );
  INVX1 U592 ( .A(n242), .Y(n247) );
  INVX1 U593 ( .A(n243), .Y(n248) );
  INVX1 U594 ( .A(n243), .Y(n249) );
  INVX1 U595 ( .A(n243), .Y(n250) );
  INVX1 U596 ( .A(n244), .Y(n251) );
  INVX1 U597 ( .A(n244), .Y(n252) );
  INVX1 U598 ( .A(n244), .Y(n253) );
  INVX1 U599 ( .A(n230), .Y(n254) );
  INVX1 U600 ( .A(n230), .Y(n255) );
  INVX1 U601 ( .A(n230), .Y(n256) );
  INVX1 U602 ( .A(n254), .Y(n257) );
  INVX1 U603 ( .A(n254), .Y(n258) );
  INVX1 U604 ( .A(n254), .Y(n259) );
  INVX1 U605 ( .A(n255), .Y(n260) );
  INVX1 U606 ( .A(n255), .Y(n261) );
  INVX1 U607 ( .A(n256), .Y(n262) );
  INVX1 U608 ( .A(n256), .Y(n263) );
  INVX1 U609 ( .A(n5180), .Y(n264) );
  INVX2 U610 ( .A(n5650), .Y(n5656) );
  AND2X2 U611 ( .A(\mem<15><1> ), .B(n205), .Y(n265) );
  INVX1 U612 ( .A(n265), .Y(n266) );
  AND2X2 U613 ( .A(n205), .B(\mem<15><3> ), .Y(n267) );
  INVX1 U614 ( .A(n267), .Y(n268) );
  AND2X2 U615 ( .A(\mem<35><7> ), .B(n201), .Y(n269) );
  INVX1 U616 ( .A(n269), .Y(n270) );
  AND2X2 U617 ( .A(\mem<56><0> ), .B(n4984), .Y(n271) );
  INVX1 U618 ( .A(n271), .Y(n272) );
  AND2X2 U619 ( .A(\mem<56><1> ), .B(n4985), .Y(n273) );
  INVX1 U620 ( .A(n273), .Y(n274) );
  AND2X2 U621 ( .A(\mem<56><3> ), .B(n4985), .Y(n275) );
  INVX1 U622 ( .A(n275), .Y(n276) );
  AND2X2 U623 ( .A(\mem<56><4> ), .B(n4984), .Y(n277) );
  INVX1 U624 ( .A(n277), .Y(n278) );
  AND2X2 U625 ( .A(\mem<56><6> ), .B(n4984), .Y(n279) );
  INVX1 U626 ( .A(n279), .Y(n280) );
  AND2X2 U627 ( .A(\mem<56><7> ), .B(n4985), .Y(n281) );
  INVX1 U628 ( .A(n281), .Y(n282) );
  AND2X2 U629 ( .A(\mem<48><3> ), .B(n6402), .Y(n283) );
  INVX1 U630 ( .A(n283), .Y(n284) );
  AND2X2 U631 ( .A(\mem<48><4> ), .B(n6402), .Y(n285) );
  INVX1 U632 ( .A(n285), .Y(n286) );
  AND2X2 U633 ( .A(\mem<48><5> ), .B(n6402), .Y(n287) );
  INVX1 U634 ( .A(n287), .Y(n288) );
  AND2X2 U635 ( .A(\mem<48><6> ), .B(n6402), .Y(n289) );
  INVX1 U636 ( .A(n289), .Y(n290) );
  AND2X2 U637 ( .A(\mem<48><7> ), .B(n6402), .Y(n291) );
  INVX1 U638 ( .A(n291), .Y(n292) );
  AND2X2 U639 ( .A(\mem<41><0> ), .B(n5010), .Y(n293) );
  INVX1 U640 ( .A(n293), .Y(n294) );
  AND2X2 U641 ( .A(\mem<41><1> ), .B(n5010), .Y(n295) );
  INVX1 U642 ( .A(n295), .Y(n296) );
  AND2X2 U643 ( .A(\mem<41><3> ), .B(n5011), .Y(n297) );
  INVX1 U644 ( .A(n297), .Y(n298) );
  AND2X2 U645 ( .A(\mem<41><4> ), .B(n5011), .Y(n299) );
  INVX1 U646 ( .A(n299), .Y(n300) );
  AND2X2 U647 ( .A(\mem<41><6> ), .B(n5011), .Y(n301) );
  INVX1 U648 ( .A(n301), .Y(n302) );
  AND2X2 U649 ( .A(\mem<41><7> ), .B(n5010), .Y(n303) );
  INVX1 U650 ( .A(n303), .Y(n304) );
  AND2X2 U651 ( .A(\mem<34><2> ), .B(n5022), .Y(n305) );
  INVX1 U652 ( .A(n305), .Y(n306) );
  AND2X2 U653 ( .A(\mem<34><5> ), .B(n5023), .Y(n307) );
  INVX1 U654 ( .A(n307), .Y(n308) );
  AND2X2 U655 ( .A(\mem<10><0> ), .B(n5060), .Y(n309) );
  INVX1 U656 ( .A(n309), .Y(n310) );
  AND2X2 U657 ( .A(\mem<10><1> ), .B(n5060), .Y(n311) );
  INVX1 U658 ( .A(n311), .Y(n312) );
  AND2X2 U659 ( .A(\mem<10><2> ), .B(n5060), .Y(n313) );
  INVX1 U660 ( .A(n313), .Y(n314) );
  AND2X2 U661 ( .A(\mem<10><4> ), .B(n5060), .Y(n315) );
  INVX1 U662 ( .A(n315), .Y(n316) );
  AND2X2 U663 ( .A(\mem<10><5> ), .B(n5060), .Y(n317) );
  INVX1 U664 ( .A(n317), .Y(n318) );
  AND2X2 U665 ( .A(\mem<10><6> ), .B(n5060), .Y(n319) );
  INVX1 U666 ( .A(n319), .Y(n320) );
  AND2X2 U667 ( .A(\mem<5><0> ), .B(n5065), .Y(n321) );
  INVX1 U668 ( .A(n321), .Y(n322) );
  AND2X2 U669 ( .A(\mem<5><1> ), .B(n5066), .Y(n323) );
  INVX1 U670 ( .A(n323), .Y(n324) );
  AND2X2 U671 ( .A(\mem<5><3> ), .B(n5066), .Y(n325) );
  INVX1 U672 ( .A(n325), .Y(n326) );
  AND2X2 U673 ( .A(\mem<5><4> ), .B(n5065), .Y(n327) );
  INVX1 U674 ( .A(n327), .Y(n328) );
  AND2X2 U675 ( .A(\mem<5><6> ), .B(n5065), .Y(n329) );
  INVX1 U676 ( .A(n329), .Y(n330) );
  AND2X2 U677 ( .A(\mem<5><7> ), .B(n5066), .Y(n331) );
  INVX1 U678 ( .A(n331), .Y(n332) );
  AND2X2 U679 ( .A(\mem<47><0> ), .B(n4998), .Y(n333) );
  INVX1 U680 ( .A(n333), .Y(n334) );
  AND2X2 U681 ( .A(\mem<47><1> ), .B(n4999), .Y(n335) );
  INVX1 U682 ( .A(n335), .Y(n336) );
  AND2X2 U683 ( .A(\mem<47><2> ), .B(n4998), .Y(n337) );
  INVX1 U684 ( .A(n337), .Y(n338) );
  AND2X2 U685 ( .A(\mem<47><3> ), .B(n4999), .Y(n339) );
  INVX1 U686 ( .A(n339), .Y(n340) );
  AND2X2 U687 ( .A(\mem<47><4> ), .B(n4998), .Y(n341) );
  INVX1 U688 ( .A(n341), .Y(n342) );
  AND2X2 U689 ( .A(\mem<47><5> ), .B(n4999), .Y(n343) );
  INVX1 U690 ( .A(n343), .Y(n344) );
  AND2X2 U691 ( .A(\mem<47><6> ), .B(n4998), .Y(n345) );
  INVX1 U692 ( .A(n345), .Y(n346) );
  AND2X2 U693 ( .A(\mem<47><7> ), .B(n4999), .Y(n347) );
  INVX1 U694 ( .A(n347), .Y(n348) );
  AND2X2 U695 ( .A(\mem<46><0> ), .B(n5000), .Y(n349) );
  INVX1 U696 ( .A(n349), .Y(n350) );
  AND2X2 U697 ( .A(\mem<46><1> ), .B(n5001), .Y(n351) );
  INVX1 U698 ( .A(n351), .Y(n352) );
  AND2X2 U699 ( .A(\mem<46><2> ), .B(n5000), .Y(n353) );
  INVX1 U700 ( .A(n353), .Y(n354) );
  AND2X2 U701 ( .A(\mem<46><3> ), .B(n5001), .Y(n355) );
  INVX1 U702 ( .A(n355), .Y(n356) );
  AND2X2 U703 ( .A(\mem<46><4> ), .B(n5000), .Y(n357) );
  INVX1 U704 ( .A(n357), .Y(n358) );
  AND2X2 U705 ( .A(\mem<46><5> ), .B(n5001), .Y(n359) );
  INVX1 U706 ( .A(n359), .Y(n360) );
  AND2X2 U707 ( .A(\mem<46><6> ), .B(n5000), .Y(n361) );
  INVX1 U708 ( .A(n361), .Y(n362) );
  AND2X2 U709 ( .A(\mem<46><7> ), .B(n5001), .Y(n363) );
  INVX1 U710 ( .A(n363), .Y(n364) );
  AND2X2 U711 ( .A(\mem<43><1> ), .B(n5007), .Y(n365) );
  INVX1 U712 ( .A(n365), .Y(n366) );
  AND2X2 U713 ( .A(\mem<43><3> ), .B(n5007), .Y(n367) );
  INVX1 U714 ( .A(n367), .Y(n368) );
  AND2X2 U715 ( .A(\mem<43><4> ), .B(n5006), .Y(n369) );
  INVX1 U716 ( .A(n369), .Y(n370) );
  AND2X2 U717 ( .A(\mem<43><6> ), .B(n5006), .Y(n371) );
  INVX1 U718 ( .A(n371), .Y(n372) );
  AND2X2 U719 ( .A(\mem<43><7> ), .B(n5007), .Y(n373) );
  INVX1 U720 ( .A(n373), .Y(n374) );
  AND2X2 U721 ( .A(\mem<41><2> ), .B(n5011), .Y(n375) );
  INVX1 U722 ( .A(n375), .Y(n376) );
  AND2X2 U723 ( .A(\mem<41><5> ), .B(n5010), .Y(n377) );
  INVX1 U724 ( .A(n377), .Y(n378) );
  AND2X2 U725 ( .A(\mem<34><0> ), .B(n5022), .Y(n379) );
  INVX1 U726 ( .A(n379), .Y(n380) );
  AND2X2 U727 ( .A(\mem<34><1> ), .B(n5022), .Y(n381) );
  INVX1 U728 ( .A(n381), .Y(n382) );
  AND2X2 U729 ( .A(\mem<34><3> ), .B(n5022), .Y(n383) );
  INVX1 U730 ( .A(n383), .Y(n384) );
  AND2X2 U731 ( .A(\mem<34><4> ), .B(n5023), .Y(n385) );
  INVX1 U732 ( .A(n385), .Y(n386) );
  AND2X2 U733 ( .A(\mem<34><6> ), .B(n5023), .Y(n387) );
  INVX1 U734 ( .A(n387), .Y(n388) );
  AND2X2 U735 ( .A(\mem<34><7> ), .B(n5023), .Y(n389) );
  INVX1 U736 ( .A(n389), .Y(n390) );
  AND2X2 U737 ( .A(\mem<35><0> ), .B(n5020), .Y(n391) );
  INVX1 U738 ( .A(n391), .Y(n392) );
  AND2X2 U739 ( .A(\mem<35><1> ), .B(n5020), .Y(n393) );
  INVX1 U740 ( .A(n393), .Y(n394) );
  AND2X2 U741 ( .A(\mem<35><3> ), .B(n5021), .Y(n395) );
  INVX1 U742 ( .A(n395), .Y(n396) );
  AND2X2 U743 ( .A(\mem<35><4> ), .B(n5021), .Y(n397) );
  INVX1 U744 ( .A(n397), .Y(n398) );
  AND2X2 U745 ( .A(\mem<35><6> ), .B(n5021), .Y(n399) );
  INVX1 U746 ( .A(n399), .Y(n400) );
  AND2X2 U747 ( .A(\mem<35><7> ), .B(n5020), .Y(n401) );
  INVX1 U748 ( .A(n401), .Y(n402) );
  INVX2 U749 ( .A(n3964), .Y(n5697) );
  INVX1 U750 ( .A(n5651), .Y(n5652) );
  INVX4 U751 ( .A(n5651), .Y(n5654) );
  INVX1 U752 ( .A(n5652), .Y(n3949) );
  INVX1 U753 ( .A(n5654), .Y(n3956) );
  INVX1 U754 ( .A(n5123), .Y(n5126) );
  AND2X2 U755 ( .A(n4162), .B(n6027), .Y(n597) );
  INVX1 U756 ( .A(n5756), .Y(n5113) );
  INVX1 U757 ( .A(n5125), .Y(n5132) );
  INVX1 U758 ( .A(n5132), .Y(n406) );
  NOR3X1 U759 ( .A(n1152), .B(\addr<7> ), .C(n3034), .Y(n403) );
  INVX1 U760 ( .A(\addr<7> ), .Y(n5772) );
  OAI21X1 U761 ( .A(n405), .B(n406), .C(n407), .Y(n404) );
  OR2X2 U762 ( .A(n5723), .B(n6043), .Y(n407) );
  INVX1 U763 ( .A(N179), .Y(n5758) );
  OR2X2 U764 ( .A(n100), .B(n3661), .Y(n408) );
  INVX1 U765 ( .A(n408), .Y(n409) );
  OR2X2 U766 ( .A(n413), .B(n411), .Y(n410) );
  OR2X2 U767 ( .A(n4251), .B(n412), .Y(n411) );
  INVX1 U768 ( .A(n5827), .Y(n412) );
  INVX1 U769 ( .A(n5828), .Y(n413) );
  OR2X2 U770 ( .A(n35), .B(n415), .Y(n414) );
  OR2X2 U771 ( .A(n4177), .B(n38), .Y(n415) );
  OR2X2 U772 ( .A(n419), .B(n417), .Y(n416) );
  OR2X2 U773 ( .A(n418), .B(n3850), .Y(n417) );
  INVX1 U774 ( .A(n5890), .Y(n418) );
  INVX1 U775 ( .A(n5891), .Y(n419) );
  OR2X2 U776 ( .A(n423), .B(n421), .Y(n420) );
  OR2X2 U777 ( .A(n422), .B(n3851), .Y(n421) );
  INVX1 U778 ( .A(n5970), .Y(n422) );
  INVX1 U779 ( .A(n5971), .Y(n423) );
  OR2X2 U780 ( .A(n36), .B(n425), .Y(n424) );
  OR2X2 U781 ( .A(n4180), .B(n39), .Y(n425) );
  OR2X2 U782 ( .A(n428), .B(n427), .Y(n426) );
  OR2X2 U783 ( .A(n4225), .B(n404), .Y(n427) );
  INVX1 U784 ( .A(n6044), .Y(n428) );
  OR2X2 U785 ( .A(n431), .B(n430), .Y(n429) );
  OR2X2 U786 ( .A(n4037), .B(n213), .Y(n430) );
  INVX1 U787 ( .A(n6121), .Y(n431) );
  OR2X2 U788 ( .A(n37), .B(n433), .Y(n432) );
  OR2X2 U789 ( .A(n4184), .B(n40), .Y(n433) );
  OR2X2 U790 ( .A(n437), .B(n435), .Y(n434) );
  OR2X2 U791 ( .A(n4038), .B(n436), .Y(n435) );
  INVX1 U792 ( .A(n6194), .Y(n436) );
  INVX1 U793 ( .A(n6195), .Y(n437) );
  OR2X2 U794 ( .A(n441), .B(n439), .Y(n438) );
  OR2X2 U795 ( .A(n440), .B(n3853), .Y(n439) );
  INVX1 U796 ( .A(n6214), .Y(n440) );
  INVX1 U797 ( .A(n6215), .Y(n441) );
  OR2X2 U798 ( .A(n445), .B(n443), .Y(n442) );
  OR2X2 U799 ( .A(n444), .B(n3855), .Y(n443) );
  INVX1 U800 ( .A(n6271), .Y(n444) );
  INVX1 U801 ( .A(n6272), .Y(n445) );
  OR2X2 U802 ( .A(n449), .B(n447), .Y(n446) );
  OR2X2 U803 ( .A(n4233), .B(n448), .Y(n447) );
  INVX1 U804 ( .A(n6350), .Y(n448) );
  INVX1 U805 ( .A(n6351), .Y(n449) );
  OR2X2 U806 ( .A(n453), .B(n451), .Y(n450) );
  OR2X2 U807 ( .A(n4234), .B(n452), .Y(n451) );
  INVX1 U808 ( .A(n6371), .Y(n452) );
  INVX1 U809 ( .A(n6372), .Y(n453) );
  OR2X2 U810 ( .A(n1659), .B(n455), .Y(n454) );
  OR2X2 U811 ( .A(n1658), .B(n3849), .Y(n455) );
  OR2X2 U812 ( .A(n1661), .B(n457), .Y(n456) );
  OR2X2 U813 ( .A(n1660), .B(n1707), .Y(n457) );
  OR2X2 U814 ( .A(n1663), .B(n459), .Y(n458) );
  OR2X2 U815 ( .A(n3031), .B(n1662), .Y(n459) );
  OR2X2 U816 ( .A(n1665), .B(n461), .Y(n460) );
  OR2X2 U817 ( .A(n1664), .B(n1709), .Y(n461) );
  OR2X2 U818 ( .A(n1667), .B(n463), .Y(n462) );
  OR2X2 U819 ( .A(n3036), .B(n1666), .Y(n463) );
  OR2X2 U820 ( .A(n1668), .B(n465), .Y(n464) );
  OR2X2 U821 ( .A(n649), .B(n206), .Y(n465) );
  OR2X2 U822 ( .A(n654), .B(n467), .Y(n466) );
  OR2X2 U823 ( .A(n1669), .B(n1670), .Y(n467) );
  OR2X2 U824 ( .A(n1672), .B(n469), .Y(n468) );
  OR2X2 U825 ( .A(n1671), .B(n1710), .Y(n469) );
  OR2X2 U826 ( .A(n1674), .B(n471), .Y(n470) );
  OR2X2 U827 ( .A(n1673), .B(n3857), .Y(n471) );
  OR2X2 U828 ( .A(n4036), .B(n1693), .Y(n473) );
  OR2X2 U829 ( .A(n1696), .B(n475), .Y(n474) );
  OR2X2 U830 ( .A(n1695), .B(n1708), .Y(n475) );
  OR2X2 U831 ( .A(n1697), .B(n477), .Y(n476) );
  OR2X2 U832 ( .A(n3035), .B(n83), .Y(n477) );
  OR2X2 U833 ( .A(n1698), .B(n3852), .Y(n479) );
  OR2X2 U834 ( .A(n1701), .B(n481), .Y(n480) );
  OR2X2 U835 ( .A(n1700), .B(n3854), .Y(n481) );
  OR2X2 U836 ( .A(n1703), .B(n483), .Y(n482) );
  OR2X2 U837 ( .A(n1702), .B(n3856), .Y(n483) );
  OR2X2 U838 ( .A(n4181), .B(n485), .Y(n484) );
  OR2X2 U839 ( .A(n3007), .B(n41), .Y(n485) );
  OR2X2 U840 ( .A(n4185), .B(n487), .Y(n486) );
  OR2X2 U841 ( .A(n3008), .B(n42), .Y(n487) );
  OR2X2 U842 ( .A(n3016), .B(n489), .Y(n488) );
  OR2X2 U843 ( .A(n4222), .B(n3015), .Y(n489) );
  OR2X2 U844 ( .A(n3018), .B(n491), .Y(n490) );
  OR2X2 U845 ( .A(n3017), .B(n641), .Y(n491) );
  OR2X2 U846 ( .A(n3020), .B(n493), .Y(n492) );
  OR2X2 U847 ( .A(n3019), .B(n644), .Y(n493) );
  OR2X2 U848 ( .A(n3022), .B(n495), .Y(n494) );
  OR2X2 U849 ( .A(n4232), .B(n3021), .Y(n495) );
  AND2X2 U850 ( .A(n6184), .B(n6183), .Y(n496) );
  OR2X2 U851 ( .A(n1142), .B(n5184), .Y(n497) );
  AND2X2 U852 ( .A(n3722), .B(n3688), .Y(n498) );
  AND2X2 U853 ( .A(n3724), .B(n3690), .Y(n499) );
  AND2X2 U854 ( .A(n3726), .B(n3692), .Y(n500) );
  AND2X2 U855 ( .A(n3728), .B(n3694), .Y(n501) );
  AND2X2 U856 ( .A(n3921), .B(n3922), .Y(n502) );
  AND2X2 U857 ( .A(n3924), .B(n3923), .Y(n503) );
  AND2X2 U858 ( .A(n3929), .B(n3930), .Y(n504) );
  AND2X2 U859 ( .A(n3696), .B(n3730), .Y(n505) );
  AND2X2 U860 ( .A(n3732), .B(n3698), .Y(n506) );
  AND2X2 U861 ( .A(n3734), .B(n3700), .Y(n507) );
  AND2X2 U862 ( .A(n3932), .B(n3933), .Y(n508) );
  AND2X2 U863 ( .A(n3937), .B(n3936), .Y(n509) );
  AND2X2 U864 ( .A(n3938), .B(n3939), .Y(n510) );
  AND2X2 U865 ( .A(n3941), .B(n3942), .Y(n511) );
  AND2X2 U866 ( .A(n3946), .B(n3945), .Y(n512) );
  AND2X2 U867 ( .A(n3736), .B(n3702), .Y(n513) );
  AND2X2 U868 ( .A(n3738), .B(n3704), .Y(n514) );
  AND2X2 U869 ( .A(n3740), .B(n3706), .Y(n515) );
  AND2X2 U870 ( .A(n3950), .B(n3951), .Y(n516) );
  OR2X2 U871 ( .A(n5724), .B(n6402), .Y(n517) );
  AND2X2 U872 ( .A(n3952), .B(n3953), .Y(n518) );
  AND2X2 U873 ( .A(n3742), .B(n1081), .Y(n519) );
  AND2X2 U874 ( .A(n3744), .B(n3708), .Y(n520) );
  AND2X2 U875 ( .A(n3962), .B(n3963), .Y(n521) );
  AND2X2 U876 ( .A(n1114), .B(n3710), .Y(n522) );
  AND2X2 U877 ( .A(n3746), .B(n3712), .Y(n523) );
  AND2X2 U878 ( .A(n3976), .B(n3975), .Y(n524) );
  AND2X2 U879 ( .A(n3978), .B(n3977), .Y(n525) );
  AND2X2 U880 ( .A(n3979), .B(n3980), .Y(n526) );
  AND2X2 U881 ( .A(n3748), .B(n1083), .Y(n527) );
  AND2X2 U882 ( .A(n3750), .B(n3714), .Y(n528) );
  AND2X2 U883 ( .A(n3752), .B(n1085), .Y(n529) );
  AND2X2 U884 ( .A(n3754), .B(n1087), .Y(n530) );
  AND2X2 U885 ( .A(n3987), .B(n3986), .Y(n531) );
  AND2X2 U886 ( .A(n3756), .B(n3716), .Y(n532) );
  AND2X2 U887 ( .A(n663), .B(n662), .Y(n533) );
  INVX1 U888 ( .A(n533), .Y(n534) );
  AND2X2 U889 ( .A(n3758), .B(n3718), .Y(n535) );
  AND2X2 U890 ( .A(n3998), .B(n3999), .Y(n536) );
  AND2X2 U891 ( .A(n5861), .B(n5860), .Y(n537) );
  OR2X2 U892 ( .A(n5772), .B(n539), .Y(n538) );
  OR2X2 U893 ( .A(n4165), .B(n4166), .Y(n539) );
  AND2X2 U894 ( .A(n541), .B(n1107), .Y(n540) );
  AND2X2 U895 ( .A(n6320), .B(n4164), .Y(n541) );
  AND2X2 U896 ( .A(n5940), .B(n5939), .Y(n542) );
  AND2X2 U897 ( .A(n6092), .B(n6091), .Y(n543) );
  AND2X2 U898 ( .A(n6241), .B(n545), .Y(n544) );
  AND2X2 U899 ( .A(n6243), .B(n6242), .Y(n545) );
  AND2X2 U900 ( .A(n6321), .B(n547), .Y(n546) );
  AND2X2 U901 ( .A(n6323), .B(n6322), .Y(n547) );
  OR2X2 U902 ( .A(n626), .B(n550), .Y(n548) );
  OR2X2 U903 ( .A(n627), .B(n605), .Y(n550) );
  OR2X2 U904 ( .A(N181), .B(n5073), .Y(n551) );
  OR2X2 U905 ( .A(N181), .B(n5074), .Y(n552) );
  AND2X2 U906 ( .A(n1111), .B(n1078), .Y(n553) );
  AND2X2 U907 ( .A(n1077), .B(n1110), .Y(n554) );
  OR2X2 U908 ( .A(N181), .B(n5078), .Y(n555) );
  OR2X2 U909 ( .A(N181), .B(n5079), .Y(n556) );
  OR2X2 U910 ( .A(n5080), .B(n3663), .Y(n557) );
  OR2X2 U911 ( .A(n5081), .B(n5086), .Y(n558) );
  OR2X2 U912 ( .A(N181), .B(n5083), .Y(n559) );
  OR2X2 U913 ( .A(n5084), .B(n5085), .Y(n560) );
  OR2X2 U914 ( .A(n5086), .B(n5087), .Y(n561) );
  OR2X2 U915 ( .A(N181), .B(n5088), .Y(n562) );
  AND2X2 U916 ( .A(n62), .B(n4959), .Y(n563) );
  OR2X2 U917 ( .A(n5089), .B(n633), .Y(n564) );
  OR2X2 U918 ( .A(n5090), .B(n5091), .Y(n565) );
  OR2X2 U919 ( .A(n5096), .B(n4945), .Y(n566) );
  INVX1 U920 ( .A(n566), .Y(\data_out<15> ) );
  OR2X2 U921 ( .A(n5098), .B(n5086), .Y(n568) );
  OR2X2 U922 ( .A(n5104), .B(n4945), .Y(n569) );
  INVX1 U923 ( .A(n569), .Y(\data_out<12> ) );
  OR2X2 U924 ( .A(n5105), .B(n4945), .Y(n571) );
  INVX1 U925 ( .A(n571), .Y(\data_out<10> ) );
  OR2X2 U926 ( .A(n5112), .B(n5091), .Y(n573) );
  AND2X2 U927 ( .A(n4116), .B(n4088), .Y(n574) );
  AND2X2 U928 ( .A(n5161), .B(n5162), .Y(n575) );
  AND2X2 U929 ( .A(n1118), .B(n4118), .Y(n576) );
  AND2X2 U930 ( .A(n4120), .B(n4122), .Y(n577) );
  AND2X2 U931 ( .A(n5166), .B(n5167), .Y(n578) );
  AND2X2 U932 ( .A(n4124), .B(n4126), .Y(n579) );
  AND2X2 U933 ( .A(n1120), .B(n76), .Y(n580) );
  INVX1 U934 ( .A(n580), .Y(n581) );
  AND2X2 U935 ( .A(n5172), .B(n5171), .Y(n582) );
  AND2X2 U936 ( .A(n4130), .B(n4128), .Y(n583) );
  AND2X2 U937 ( .A(n551), .B(n561), .Y(n584) );
  AND2X2 U938 ( .A(n4132), .B(n4090), .Y(n585) );
  AND2X2 U939 ( .A(n4092), .B(n1089), .Y(n586) );
  AND2X2 U940 ( .A(n3760), .B(n1091), .Y(n587) );
  AND2X2 U941 ( .A(n1093), .B(n4134), .Y(n588) );
  AND2X2 U942 ( .A(n552), .B(n560), .Y(n589) );
  OR2X2 U943 ( .A(N178), .B(n25), .Y(n590) );
  INVX1 U944 ( .A(n590), .Y(n591) );
  AND2X2 U945 ( .A(n5911), .B(n5912), .Y(n592) );
  AND2X2 U946 ( .A(n6139), .B(n6140), .Y(n593) );
  AND2X2 U947 ( .A(n593), .B(n4110), .Y(n594) );
  INVX1 U948 ( .A(n594), .Y(n595) );
  AND2X2 U949 ( .A(n4136), .B(n1095), .Y(n598) );
  AND2X2 U950 ( .A(n555), .B(n568), .Y(n599) );
  AND2X2 U951 ( .A(n4138), .B(n4140), .Y(n600) );
  AND2X2 U952 ( .A(n4142), .B(n4094), .Y(n601) );
  AND2X2 U953 ( .A(n5870), .B(n4160), .Y(n602) );
  AND2X2 U954 ( .A(n4144), .B(n4146), .Y(n603) );
  AND2X2 U955 ( .A(n4148), .B(n4096), .Y(n604) );
  OR2X2 U956 ( .A(n5724), .B(n3925), .Y(n605) );
  AND2X2 U957 ( .A(n5199), .B(n5198), .Y(n606) );
  AND2X2 U958 ( .A(n558), .B(n559), .Y(n607) );
  AND2X2 U959 ( .A(n5200), .B(n5201), .Y(n608) );
  AND2X2 U960 ( .A(n5202), .B(n5203), .Y(n609) );
  AND2X2 U961 ( .A(n4150), .B(n4098), .Y(n610) );
  AND2X2 U962 ( .A(n4152), .B(n4100), .Y(n611) );
  AND2X2 U963 ( .A(n4154), .B(n4102), .Y(n612) );
  AND2X2 U964 ( .A(n5210), .B(n5211), .Y(n613) );
  AND2X2 U965 ( .A(n565), .B(n562), .Y(n614) );
  AND2X2 U966 ( .A(n4156), .B(n4104), .Y(n615) );
  OR2X2 U967 ( .A(n89), .B(n1143), .Y(n616) );
  AND2X2 U968 ( .A(n5214), .B(n5213), .Y(n618) );
  AND2X2 U969 ( .A(n4158), .B(n1097), .Y(n619) );
  AND2X2 U970 ( .A(n573), .B(n556), .Y(n620) );
  OR2X2 U971 ( .A(\addr<6> ), .B(\addr<8> ), .Y(n621) );
  OR2X2 U972 ( .A(n5757), .B(n5704), .Y(n622) );
  INVX1 U973 ( .A(n622), .Y(n623) );
  OR2X2 U974 ( .A(n1134), .B(n1145), .Y(n624) );
  INVX1 U975 ( .A(n624), .Y(n625) );
  OR2X2 U976 ( .A(n538), .B(n4942), .Y(n626) );
  OR2X2 U977 ( .A(n4167), .B(n1140), .Y(n627) );
  OR2X2 U978 ( .A(N182), .B(n5759), .Y(n628) );
  INVX1 U979 ( .A(n628), .Y(n629) );
  AND2X2 U980 ( .A(n5759), .B(n5151), .Y(n630) );
  AND2X2 U981 ( .A(n5832), .B(n5843), .Y(n631) );
  INVX1 U982 ( .A(n631), .Y(n632) );
  OR2X2 U983 ( .A(n632), .B(\addr<15> ), .Y(n633) );
  OR2X2 U984 ( .A(n4169), .B(\addr<15> ), .Y(n634) );
  AND2X2 U985 ( .A(n5863), .B(n5862), .Y(n635) );
  AND2X2 U986 ( .A(n5869), .B(n5868), .Y(n636) );
  INVX1 U987 ( .A(n637), .Y(n638) );
  AND2X2 U988 ( .A(n5943), .B(n5942), .Y(n639) );
  AND2X2 U989 ( .A(n5949), .B(n5948), .Y(n640) );
  OR2X2 U990 ( .A(n5988), .B(n5987), .Y(n641) );
  AND2X2 U991 ( .A(n6019), .B(n6020), .Y(n642) );
  AND2X2 U992 ( .A(n6026), .B(n6025), .Y(n643) );
  OR2X2 U993 ( .A(n6061), .B(n6062), .Y(n644) );
  AND2X2 U994 ( .A(n1124), .B(n1101), .Y(n645) );
  INVX1 U995 ( .A(n645), .Y(n646) );
  AND2X2 U996 ( .A(n6095), .B(n6094), .Y(n647) );
  AND2X2 U997 ( .A(n6101), .B(n6100), .Y(n648) );
  OR2X2 U998 ( .A(n6127), .B(n6126), .Y(n649) );
  AND2X2 U999 ( .A(n1126), .B(n3720), .Y(n650) );
  INVX1 U1000 ( .A(n650), .Y(n651) );
  AND2X2 U1001 ( .A(n6166), .B(n6165), .Y(n652) );
  AND2X2 U1002 ( .A(n6172), .B(n6171), .Y(n653) );
  OR2X2 U1003 ( .A(n6200), .B(n6201), .Y(n654) );
  AND2X2 U1004 ( .A(n1112), .B(n1079), .Y(n655) );
  AND2X2 U1005 ( .A(n1128), .B(n1103), .Y(n656) );
  INVX1 U1006 ( .A(n656), .Y(n657) );
  AND2X2 U1007 ( .A(n6246), .B(n6245), .Y(n658) );
  AND2X2 U1008 ( .A(n6252), .B(n6251), .Y(n659) );
  AND2X2 U1009 ( .A(n1130), .B(n1105), .Y(n660) );
  INVX1 U1010 ( .A(n660), .Y(n661) );
  AND2X2 U1011 ( .A(n6325), .B(n6324), .Y(n662) );
  AND2X2 U1012 ( .A(n6331), .B(n6330), .Y(n663) );
  AND2X2 U1013 ( .A(n1132), .B(n1109), .Y(n664) );
  INVX1 U1014 ( .A(n664), .Y(n665) );
  AND2X2 U1015 ( .A(n3928), .B(n4953), .Y(n666) );
  AND2X2 U1016 ( .A(n3928), .B(n4960), .Y(n667) );
  AND2X2 U1017 ( .A(n3927), .B(n4956), .Y(n668) );
  AND2X2 U1018 ( .A(n3928), .B(n4962), .Y(n669) );
  AND2X2 U1019 ( .A(n3927), .B(n4964), .Y(n670) );
  AND2X2 U1020 ( .A(n3927), .B(n4966), .Y(n671) );
  AND2X2 U1021 ( .A(n3928), .B(n4949), .Y(n672) );
  AND2X2 U1022 ( .A(n6401), .B(n6457), .Y(n673) );
  INVX1 U1023 ( .A(n673), .Y(n674) );
  AND2X2 U1024 ( .A(n5702), .B(n4954), .Y(n675) );
  AND2X2 U1025 ( .A(n5702), .B(n4958), .Y(n676) );
  AND2X2 U1026 ( .A(n5700), .B(n4956), .Y(n677) );
  AND2X2 U1027 ( .A(n5176), .B(n4962), .Y(n678) );
  AND2X2 U1028 ( .A(\data_in<0> ), .B(n1551), .Y(n679) );
  INVX1 U1029 ( .A(n679), .Y(n680) );
  AND2X2 U1030 ( .A(n1551), .B(\data_in<1> ), .Y(n681) );
  INVX1 U1031 ( .A(n681), .Y(n682) );
  AND2X2 U1032 ( .A(\data_in<3> ), .B(n1551), .Y(n683) );
  INVX1 U1033 ( .A(n683), .Y(n684) );
  AND2X2 U1034 ( .A(\data_in<4> ), .B(n1551), .Y(n685) );
  INVX1 U1035 ( .A(n685), .Y(n686) );
  AND2X2 U1036 ( .A(\data_in<6> ), .B(n1551), .Y(n687) );
  INVX1 U1037 ( .A(n687), .Y(n688) );
  AND2X2 U1038 ( .A(\data_in<7> ), .B(n1551), .Y(n689) );
  INVX1 U1039 ( .A(n689), .Y(n690) );
  AND2X2 U1040 ( .A(n5177), .B(n4964), .Y(n691) );
  AND2X2 U1041 ( .A(n5176), .B(n4966), .Y(n692) );
  AND2X2 U1042 ( .A(n5177), .B(n4949), .Y(n693) );
  AND2X2 U1043 ( .A(n54), .B(n5726), .Y(n694) );
  INVX1 U1044 ( .A(n694), .Y(n695) );
  AND2X2 U1045 ( .A(n28), .B(n4952), .Y(n696) );
  AND2X2 U1046 ( .A(\data_in<8> ), .B(n1561), .Y(n697) );
  INVX1 U1047 ( .A(n697), .Y(n698) );
  AND2X2 U1048 ( .A(\data_in<9> ), .B(n1561), .Y(n699) );
  INVX1 U1049 ( .A(n699), .Y(n700) );
  AND2X2 U1050 ( .A(\data_in<10> ), .B(n1561), .Y(n701) );
  INVX1 U1051 ( .A(n701), .Y(n702) );
  AND2X2 U1052 ( .A(\data_in<11> ), .B(n1561), .Y(n703) );
  INVX1 U1053 ( .A(n703), .Y(n704) );
  AND2X2 U1054 ( .A(\data_in<12> ), .B(n1561), .Y(n705) );
  INVX1 U1055 ( .A(n705), .Y(n706) );
  AND2X2 U1056 ( .A(\data_in<13> ), .B(n1561), .Y(n707) );
  INVX1 U1057 ( .A(n707), .Y(n708) );
  AND2X2 U1058 ( .A(n1561), .B(\data_in<14> ), .Y(n709) );
  INVX1 U1059 ( .A(n709), .Y(n710) );
  AND2X2 U1060 ( .A(\data_in<15> ), .B(n1561), .Y(n711) );
  INVX1 U1061 ( .A(n711), .Y(n712) );
  AND2X2 U1062 ( .A(n68), .B(n4959), .Y(n713) );
  AND2X2 U1063 ( .A(\data_in<8> ), .B(n1563), .Y(n714) );
  AND2X2 U1064 ( .A(\data_in<9> ), .B(n1563), .Y(n715) );
  AND2X2 U1065 ( .A(\data_in<10> ), .B(n14), .Y(n716) );
  INVX1 U1066 ( .A(n716), .Y(n717) );
  AND2X2 U1067 ( .A(\data_in<11> ), .B(n14), .Y(n718) );
  INVX1 U1068 ( .A(n718), .Y(n719) );
  AND2X2 U1069 ( .A(\data_in<12> ), .B(n1563), .Y(n720) );
  INVX1 U1070 ( .A(n720), .Y(n721) );
  AND2X2 U1071 ( .A(\data_in<13> ), .B(n1563), .Y(n722) );
  INVX1 U1072 ( .A(n722), .Y(n723) );
  AND2X2 U1073 ( .A(\data_in<14> ), .B(n14), .Y(n724) );
  INVX1 U1074 ( .A(n724), .Y(n725) );
  AND2X2 U1075 ( .A(\data_in<15> ), .B(n14), .Y(n726) );
  INVX1 U1076 ( .A(n726), .Y(n727) );
  AND2X2 U1077 ( .A(n28), .B(n4956), .Y(n728) );
  AND2X2 U1078 ( .A(\data_in<8> ), .B(n1565), .Y(n729) );
  AND2X2 U1079 ( .A(\data_in<9> ), .B(n1565), .Y(n730) );
  INVX1 U1080 ( .A(n730), .Y(n731) );
  AND2X2 U1081 ( .A(\data_in<11> ), .B(n1565), .Y(n732) );
  INVX1 U1082 ( .A(n732), .Y(n733) );
  AND2X2 U1083 ( .A(\data_in<12> ), .B(n1565), .Y(n734) );
  INVX1 U1084 ( .A(n734), .Y(n735) );
  AND2X2 U1085 ( .A(\data_in<14> ), .B(n1565), .Y(n736) );
  INVX1 U1086 ( .A(n736), .Y(n737) );
  AND2X2 U1087 ( .A(\data_in<15> ), .B(n1565), .Y(n738) );
  INVX1 U1088 ( .A(n738), .Y(n739) );
  AND2X2 U1089 ( .A(n61), .B(n4962), .Y(n740) );
  AND2X2 U1090 ( .A(\data_in<8> ), .B(n13), .Y(n741) );
  INVX1 U1091 ( .A(n741), .Y(n742) );
  AND2X2 U1092 ( .A(\data_in<9> ), .B(n1567), .Y(n743) );
  AND2X2 U1093 ( .A(\data_in<11> ), .B(n1567), .Y(n744) );
  INVX1 U1094 ( .A(n744), .Y(n745) );
  AND2X2 U1095 ( .A(\data_in<12> ), .B(n13), .Y(n746) );
  INVX1 U1096 ( .A(n746), .Y(n747) );
  AND2X2 U1097 ( .A(\data_in<14> ), .B(n13), .Y(n748) );
  INVX1 U1098 ( .A(n748), .Y(n749) );
  AND2X2 U1099 ( .A(\data_in<15> ), .B(n1567), .Y(n750) );
  INVX1 U1100 ( .A(n750), .Y(n751) );
  AND2X2 U1101 ( .A(n61), .B(n4964), .Y(n752) );
  AND2X2 U1102 ( .A(\data_in<8> ), .B(n1569), .Y(n753) );
  INVX1 U1103 ( .A(n753), .Y(n754) );
  AND2X2 U1104 ( .A(\data_in<9> ), .B(n1569), .Y(n755) );
  INVX1 U1105 ( .A(n755), .Y(n756) );
  AND2X2 U1106 ( .A(\data_in<11> ), .B(n1569), .Y(n757) );
  INVX1 U1107 ( .A(n757), .Y(n758) );
  AND2X2 U1108 ( .A(\data_in<12> ), .B(n1569), .Y(n759) );
  INVX1 U1109 ( .A(n759), .Y(n760) );
  AND2X2 U1110 ( .A(\data_in<14> ), .B(n1569), .Y(n761) );
  INVX1 U1111 ( .A(n761), .Y(n762) );
  AND2X2 U1112 ( .A(\data_in<15> ), .B(n1569), .Y(n763) );
  INVX1 U1113 ( .A(n763), .Y(n764) );
  AND2X2 U1114 ( .A(n54), .B(n4966), .Y(n765) );
  AND2X2 U1115 ( .A(\data_in<8> ), .B(n64), .Y(n766) );
  AND2X2 U1116 ( .A(\data_in<9> ), .B(n1571), .Y(n767) );
  INVX1 U1117 ( .A(n767), .Y(n768) );
  AND2X2 U1118 ( .A(\data_in<11> ), .B(n64), .Y(n769) );
  INVX1 U1119 ( .A(n769), .Y(n770) );
  AND2X2 U1120 ( .A(\data_in<12> ), .B(n64), .Y(n771) );
  INVX1 U1121 ( .A(n771), .Y(n772) );
  AND2X2 U1122 ( .A(\data_in<14> ), .B(n1571), .Y(n773) );
  INVX1 U1123 ( .A(n773), .Y(n774) );
  AND2X2 U1124 ( .A(\data_in<15> ), .B(n64), .Y(n775) );
  INVX1 U1125 ( .A(n775), .Y(n776) );
  AND2X2 U1126 ( .A(n68), .B(n4950), .Y(n777) );
  AND2X2 U1127 ( .A(\data_in<10> ), .B(n1573), .Y(n778) );
  INVX1 U1128 ( .A(n778), .Y(n779) );
  AND2X2 U1129 ( .A(\data_in<13> ), .B(n1573), .Y(n780) );
  INVX1 U1130 ( .A(n780), .Y(n781) );
  AND2X2 U1131 ( .A(n6423), .B(n6457), .Y(n782) );
  AND2X2 U1132 ( .A(n4946), .B(n4953), .Y(n783) );
  AND2X2 U1133 ( .A(\data_in<0> ), .B(n49), .Y(n784) );
  INVX1 U1134 ( .A(n784), .Y(n785) );
  AND2X2 U1135 ( .A(\data_in<8> ), .B(n1575), .Y(n786) );
  INVX1 U1136 ( .A(n786), .Y(n787) );
  AND2X2 U1137 ( .A(\data_in<1> ), .B(n49), .Y(n788) );
  INVX1 U1138 ( .A(n788), .Y(n789) );
  AND2X2 U1139 ( .A(\data_in<9> ), .B(n1575), .Y(n790) );
  INVX1 U1140 ( .A(n790), .Y(n791) );
  AND2X2 U1141 ( .A(\data_in<3> ), .B(n49), .Y(n792) );
  INVX1 U1142 ( .A(n792), .Y(n793) );
  AND2X2 U1143 ( .A(\data_in<11> ), .B(n1575), .Y(n794) );
  INVX1 U1144 ( .A(n794), .Y(n795) );
  AND2X2 U1145 ( .A(\data_in<4> ), .B(n49), .Y(n796) );
  INVX1 U1146 ( .A(n796), .Y(n797) );
  AND2X2 U1147 ( .A(\data_in<12> ), .B(n1575), .Y(n798) );
  INVX1 U1148 ( .A(n798), .Y(n799) );
  AND2X2 U1149 ( .A(\data_in<6> ), .B(n49), .Y(n800) );
  INVX1 U1150 ( .A(n800), .Y(n801) );
  AND2X2 U1151 ( .A(\data_in<14> ), .B(n1575), .Y(n802) );
  INVX1 U1152 ( .A(n802), .Y(n803) );
  AND2X2 U1153 ( .A(\data_in<7> ), .B(n49), .Y(n804) );
  INVX1 U1154 ( .A(n804), .Y(n805) );
  AND2X2 U1155 ( .A(\data_in<15> ), .B(n1575), .Y(n806) );
  INVX1 U1156 ( .A(n806), .Y(n807) );
  AND2X2 U1157 ( .A(n5156), .B(n4960), .Y(n808) );
  AND2X2 U1158 ( .A(n5156), .B(n4956), .Y(n809) );
  AND2X2 U1159 ( .A(n4962), .B(n5156), .Y(n810) );
  AND2X2 U1160 ( .A(n29), .B(n4964), .Y(n811) );
  AND2X2 U1161 ( .A(n4966), .B(n4946), .Y(n812) );
  AND2X2 U1162 ( .A(\data_in<8> ), .B(n1585), .Y(n813) );
  AND2X2 U1163 ( .A(\data_in<9> ), .B(n9), .Y(n814) );
  INVX1 U1164 ( .A(n814), .Y(n815) );
  AND2X2 U1165 ( .A(\data_in<11> ), .B(n1585), .Y(n816) );
  INVX1 U1166 ( .A(n816), .Y(n817) );
  AND2X2 U1167 ( .A(\data_in<12> ), .B(n1585), .Y(n818) );
  INVX1 U1168 ( .A(n818), .Y(n819) );
  AND2X2 U1169 ( .A(\data_in<14> ), .B(n9), .Y(n820) );
  INVX1 U1170 ( .A(n820), .Y(n821) );
  AND2X2 U1171 ( .A(\data_in<15> ), .B(n9), .Y(n822) );
  INVX1 U1172 ( .A(n822), .Y(n823) );
  AND2X2 U1173 ( .A(n5156), .B(n4949), .Y(n824) );
  AND2X2 U1174 ( .A(n4953), .B(n5708), .Y(n825) );
  AND2X2 U1175 ( .A(n15), .B(n4958), .Y(n826) );
  AND2X2 U1176 ( .A(n4956), .B(n3983), .Y(n828) );
  AND2X2 U1177 ( .A(n15), .B(n4962), .Y(n829) );
  AND2X2 U1178 ( .A(n4964), .B(n3981), .Y(n830) );
  AND2X2 U1179 ( .A(n4966), .B(n5708), .Y(n831) );
  AND2X2 U1180 ( .A(n4949), .B(n3983), .Y(n832) );
  AND2X2 U1181 ( .A(n6428), .B(n6457), .Y(n833) );
  AND2X2 U1182 ( .A(n5194), .B(n4954), .Y(n834) );
  AND2X2 U1183 ( .A(n5194), .B(n4958), .Y(n835) );
  AND2X2 U1184 ( .A(n5194), .B(n4956), .Y(n836) );
  AND2X2 U1185 ( .A(n5194), .B(n4962), .Y(n837) );
  AND2X2 U1186 ( .A(\data_in<0> ), .B(n44), .Y(n838) );
  INVX1 U1187 ( .A(n838), .Y(n839) );
  AND2X2 U1188 ( .A(\data_in<8> ), .B(n8), .Y(n840) );
  INVX1 U1189 ( .A(n840), .Y(n841) );
  AND2X2 U1190 ( .A(\data_in<1> ), .B(n1612), .Y(n842) );
  INVX1 U1191 ( .A(n842), .Y(n843) );
  AND2X2 U1192 ( .A(\data_in<9> ), .B(n8), .Y(n844) );
  AND2X2 U1193 ( .A(\data_in<2> ), .B(n1612), .Y(n845) );
  INVX1 U1194 ( .A(n845), .Y(n846) );
  AND2X2 U1195 ( .A(\data_in<10> ), .B(n8), .Y(n847) );
  INVX1 U1196 ( .A(n847), .Y(n848) );
  AND2X2 U1197 ( .A(\data_in<3> ), .B(n44), .Y(n849) );
  INVX1 U1198 ( .A(n849), .Y(n850) );
  AND2X2 U1199 ( .A(\data_in<11> ), .B(n1613), .Y(n851) );
  INVX1 U1200 ( .A(n851), .Y(n852) );
  AND2X2 U1201 ( .A(\data_in<4> ), .B(n44), .Y(n853) );
  INVX1 U1202 ( .A(n853), .Y(n854) );
  AND2X2 U1203 ( .A(\data_in<12> ), .B(n1613), .Y(n855) );
  INVX1 U1204 ( .A(n855), .Y(n856) );
  AND2X2 U1205 ( .A(\data_in<5> ), .B(n1612), .Y(n857) );
  INVX1 U1206 ( .A(n857), .Y(n858) );
  AND2X2 U1207 ( .A(\data_in<13> ), .B(n1613), .Y(n859) );
  INVX1 U1208 ( .A(n859), .Y(n860) );
  AND2X2 U1209 ( .A(\data_in<6> ), .B(n1612), .Y(n861) );
  INVX1 U1210 ( .A(n861), .Y(n862) );
  AND2X2 U1211 ( .A(\data_in<14> ), .B(n1613), .Y(n863) );
  INVX1 U1212 ( .A(n863), .Y(n864) );
  AND2X2 U1213 ( .A(\data_in<7> ), .B(n44), .Y(n865) );
  INVX1 U1214 ( .A(n865), .Y(n866) );
  AND2X2 U1215 ( .A(\data_in<15> ), .B(n8), .Y(n867) );
  INVX1 U1216 ( .A(n867), .Y(n868) );
  AND2X2 U1217 ( .A(n5194), .B(n4964), .Y(n869) );
  AND2X2 U1218 ( .A(n5194), .B(n4966), .Y(n870) );
  AND2X2 U1219 ( .A(n5194), .B(n4950), .Y(n871) );
  AND2X2 U1220 ( .A(n6430), .B(n6457), .Y(n872) );
  AND2X2 U1221 ( .A(n4952), .B(n66), .Y(n873) );
  AND2X2 U1222 ( .A(n5205), .B(n4956), .Y(n874) );
  AND2X2 U1223 ( .A(n5207), .B(n4962), .Y(n875) );
  AND2X2 U1224 ( .A(n5205), .B(n4964), .Y(n876) );
  AND2X2 U1225 ( .A(n4966), .B(n5207), .Y(n877) );
  AND2X2 U1226 ( .A(n66), .B(n4949), .Y(n878) );
  AND2X2 U1227 ( .A(n6440), .B(n6457), .Y(n879) );
  AND2X2 U1228 ( .A(\data_in<0> ), .B(n1634), .Y(n881) );
  INVX1 U1229 ( .A(n881), .Y(n882) );
  AND2X2 U1230 ( .A(\data_in<1> ), .B(n1634), .Y(n883) );
  AND2X2 U1231 ( .A(\data_in<2> ), .B(n1634), .Y(n884) );
  INVX1 U1232 ( .A(n884), .Y(n885) );
  AND2X2 U1233 ( .A(\data_in<3> ), .B(n1634), .Y(n886) );
  INVX1 U1234 ( .A(n886), .Y(n887) );
  AND2X2 U1235 ( .A(\data_in<4> ), .B(n1634), .Y(n888) );
  INVX1 U1236 ( .A(n888), .Y(n889) );
  AND2X2 U1237 ( .A(\data_in<5> ), .B(n1634), .Y(n890) );
  INVX1 U1238 ( .A(n890), .Y(n891) );
  AND2X2 U1239 ( .A(\data_in<6> ), .B(n1634), .Y(n892) );
  INVX1 U1240 ( .A(n892), .Y(n893) );
  AND2X2 U1241 ( .A(\data_in<7> ), .B(n1634), .Y(n894) );
  INVX1 U1242 ( .A(n894), .Y(n895) );
  AND2X2 U1243 ( .A(n5181), .B(n4952), .Y(n896) );
  AND2X2 U1244 ( .A(n33), .B(n4959), .Y(n897) );
  INVX1 U1245 ( .A(n897), .Y(n898) );
  AND2X2 U1246 ( .A(n33), .B(n4956), .Y(n899) );
  AND2X2 U1247 ( .A(n33), .B(n4962), .Y(n900) );
  AND2X2 U1248 ( .A(n5181), .B(n4964), .Y(n901) );
  AND2X2 U1249 ( .A(n33), .B(n4966), .Y(n902) );
  AND2X2 U1250 ( .A(n5181), .B(n4114), .Y(n903) );
  INVX1 U1251 ( .A(n903), .Y(n904) );
  BUFX2 U1252 ( .A(n6141), .Y(n905) );
  AND2X2 U1253 ( .A(n648), .B(n647), .Y(n906) );
  INVX1 U1254 ( .A(n906), .Y(n907) );
  AND2X2 U1255 ( .A(n1116), .B(n75), .Y(n908) );
  INVX1 U1256 ( .A(n908), .Y(n909) );
  AND2X2 U1257 ( .A(n546), .B(n540), .Y(n910) );
  INVX1 U1258 ( .A(n910), .Y(n911) );
  AND2X2 U1259 ( .A(n4216), .B(n544), .Y(n912) );
  INVX1 U1260 ( .A(n912), .Y(n913) );
  AND2X2 U1261 ( .A(n659), .B(n658), .Y(n914) );
  INVX1 U1262 ( .A(n914), .Y(n915) );
  INVX1 U1263 ( .A(n916), .Y(n917) );
  AND2X2 U1264 ( .A(n642), .B(n643), .Y(n918) );
  INVX1 U1265 ( .A(n918), .Y(n919) );
  OR2X2 U1266 ( .A(n5781), .B(n5780), .Y(n920) );
  INVX1 U1267 ( .A(n920), .Y(n921) );
  OR2X2 U1268 ( .A(\addr<15> ), .B(n4175), .Y(n922) );
  INVX1 U1269 ( .A(n922), .Y(n923) );
  OR2X2 U1270 ( .A(n5835), .B(n5836), .Y(n924) );
  INVX1 U1271 ( .A(n924), .Y(n925) );
  OR2X2 U1272 ( .A(n5849), .B(n5848), .Y(n926) );
  INVX1 U1273 ( .A(n926), .Y(n927) );
  OR2X2 U1274 ( .A(n5925), .B(n5924), .Y(n928) );
  INVX1 U1275 ( .A(n928), .Y(n929) );
  OR2X2 U1276 ( .A(n6010), .B(n6009), .Y(n930) );
  INVX1 U1277 ( .A(n930), .Y(n931) );
  OR2X2 U1278 ( .A(n6148), .B(n6147), .Y(n932) );
  INVX1 U1279 ( .A(n932), .Y(n933) );
  OR2X2 U1280 ( .A(n6179), .B(n6180), .Y(n934) );
  INVX1 U1281 ( .A(n934), .Y(n935) );
  OR2X2 U1282 ( .A(n6222), .B(n6221), .Y(n936) );
  INVX1 U1283 ( .A(n936), .Y(n937) );
  OR2X2 U1284 ( .A(n6300), .B(n6299), .Y(n938) );
  INVX1 U1285 ( .A(n938), .Y(n939) );
  OR2X2 U1286 ( .A(n6385), .B(n6384), .Y(n940) );
  INVX1 U1287 ( .A(n940), .Y(n941) );
  BUFX2 U1288 ( .A(n6142), .Y(n942) );
  AND2X2 U1289 ( .A(n635), .B(n636), .Y(n943) );
  INVX1 U1290 ( .A(n943), .Y(n944) );
  AND2X2 U1291 ( .A(\mem<31><3> ), .B(n225), .Y(n945) );
  INVX1 U1292 ( .A(n945), .Y(n946) );
  AND2X2 U1293 ( .A(\mem<31><1> ), .B(n223), .Y(n947) );
  INVX1 U1294 ( .A(n947), .Y(n948) );
  OR2X2 U1295 ( .A(\addr<13> ), .B(n621), .Y(n949) );
  INVX1 U1296 ( .A(n949), .Y(n950) );
  OR2X2 U1297 ( .A(n5842), .B(n5841), .Y(n951) );
  INVX1 U1298 ( .A(n951), .Y(n952) );
  OR2X2 U1299 ( .A(n5855), .B(n5854), .Y(n953) );
  INVX1 U1300 ( .A(n953), .Y(n954) );
  OR2X2 U1301 ( .A(n5919), .B(n5918), .Y(n955) );
  INVX1 U1302 ( .A(n955), .Y(n956) );
  OR2X2 U1303 ( .A(n6005), .B(n6004), .Y(n957) );
  INVX1 U1304 ( .A(n957), .Y(n958) );
  OR2X2 U1305 ( .A(n6015), .B(n6014), .Y(n959) );
  INVX1 U1306 ( .A(n959), .Y(n960) );
  OR2X2 U1307 ( .A(n6076), .B(n6075), .Y(n961) );
  INVX1 U1308 ( .A(n961), .Y(n962) );
  OR2X2 U1309 ( .A(n6153), .B(n6152), .Y(n963) );
  INVX1 U1310 ( .A(n963), .Y(n964) );
  OR2X2 U1311 ( .A(n6227), .B(n6226), .Y(n965) );
  INVX1 U1312 ( .A(n965), .Y(n966) );
  OR2X2 U1313 ( .A(n6306), .B(n6305), .Y(n967) );
  INVX1 U1314 ( .A(n967), .Y(n968) );
  OR2X2 U1315 ( .A(n6380), .B(n6379), .Y(n969) );
  INVX1 U1316 ( .A(n969), .Y(n970) );
  AND2X2 U1317 ( .A(\mem<11><0> ), .B(n194), .Y(n971) );
  INVX1 U1318 ( .A(n971), .Y(n972) );
  AND2X2 U1319 ( .A(\mem<15><0> ), .B(n77), .Y(n973) );
  INVX1 U1320 ( .A(n973), .Y(n974) );
  AND2X2 U1321 ( .A(\mem<39><0> ), .B(n617), .Y(n975) );
  INVX1 U1322 ( .A(n975), .Y(n976) );
  AND2X2 U1323 ( .A(\mem<19><0> ), .B(n186), .Y(n977) );
  INVX1 U1324 ( .A(n977), .Y(n978) );
  AND2X2 U1325 ( .A(\mem<23><0> ), .B(n77), .Y(n979) );
  INVX1 U1326 ( .A(n979), .Y(n980) );
  AND2X2 U1327 ( .A(n77), .B(\mem<55><0> ), .Y(n981) );
  INVX1 U1328 ( .A(n981), .Y(n982) );
  AND2X2 U1329 ( .A(\mem<4><0> ), .B(n161), .Y(n983) );
  INVX1 U1330 ( .A(n983), .Y(n984) );
  AND2X2 U1331 ( .A(\mem<35><1> ), .B(n185), .Y(n985) );
  INVX1 U1332 ( .A(n985), .Y(n986) );
  AND2X2 U1333 ( .A(n77), .B(\mem<39><1> ), .Y(n987) );
  INVX1 U1334 ( .A(n987), .Y(n988) );
  AND2X2 U1335 ( .A(\mem<23><1> ), .B(n205), .Y(n989) );
  INVX1 U1336 ( .A(n989), .Y(n990) );
  AND2X2 U1337 ( .A(\mem<55><1> ), .B(n79), .Y(n991) );
  INVX1 U1338 ( .A(n991), .Y(n992) );
  AND2X2 U1339 ( .A(\mem<47><1> ), .B(n3685), .Y(n993) );
  INVX1 U1340 ( .A(n993), .Y(n994) );
  AND2X2 U1341 ( .A(\mem<11><2> ), .B(n196), .Y(n995) );
  INVX1 U1342 ( .A(n995), .Y(n996) );
  AND2X2 U1343 ( .A(\mem<35><2> ), .B(n200), .Y(n997) );
  INVX1 U1344 ( .A(n997), .Y(n998) );
  AND2X2 U1345 ( .A(\mem<39><2> ), .B(n77), .Y(n999) );
  INVX1 U1346 ( .A(n999), .Y(n1000) );
  AND2X2 U1347 ( .A(\mem<19><2> ), .B(n193), .Y(n1001) );
  INVX1 U1348 ( .A(n1001), .Y(n1002) );
  AND2X2 U1349 ( .A(\mem<23><2> ), .B(n77), .Y(n1003) );
  INVX1 U1350 ( .A(n1003), .Y(n1004) );
  AND2X2 U1351 ( .A(\mem<55><2> ), .B(n77), .Y(n1005) );
  INVX1 U1352 ( .A(n1005), .Y(n1006) );
  AND2X2 U1353 ( .A(\mem<4><2> ), .B(n155), .Y(n1007) );
  INVX1 U1354 ( .A(n1007), .Y(n1008) );
  AND2X2 U1355 ( .A(\mem<47><2> ), .B(n225), .Y(n1009) );
  INVX1 U1356 ( .A(n1009), .Y(n1010) );
  AND2X2 U1357 ( .A(\mem<39><3> ), .B(n105), .Y(n1011) );
  INVX1 U1358 ( .A(n1011), .Y(n1012) );
  AND2X2 U1359 ( .A(\mem<23><3> ), .B(n205), .Y(n1013) );
  INVX1 U1360 ( .A(n1013), .Y(n1014) );
  AND2X2 U1361 ( .A(\mem<55><3> ), .B(n77), .Y(n1015) );
  INVX1 U1362 ( .A(n1015), .Y(n1016) );
  AND2X2 U1363 ( .A(\mem<47><3> ), .B(n3685), .Y(n1017) );
  INVX1 U1364 ( .A(n1017), .Y(n1018) );
  AND2X2 U1365 ( .A(\mem<11><4> ), .B(n184), .Y(n1019) );
  INVX1 U1366 ( .A(n1019), .Y(n1020) );
  AND2X2 U1367 ( .A(n205), .B(\mem<15><4> ), .Y(n1021) );
  INVX1 U1368 ( .A(n1021), .Y(n1022) );
  AND2X2 U1369 ( .A(n77), .B(\mem<39><4> ), .Y(n1023) );
  INVX1 U1370 ( .A(n1023), .Y(n1024) );
  AND2X2 U1371 ( .A(n183), .B(\mem<19><4> ), .Y(n1025) );
  INVX1 U1372 ( .A(n1025), .Y(n1026) );
  AND2X2 U1373 ( .A(n77), .B(\mem<23><4> ), .Y(n1027) );
  INVX1 U1374 ( .A(n1027), .Y(n1028) );
  AND2X2 U1375 ( .A(\mem<55><4> ), .B(n79), .Y(n1029) );
  INVX1 U1376 ( .A(n1029), .Y(n1030) );
  AND2X2 U1377 ( .A(\mem<7><4> ), .B(n224), .Y(n1031) );
  INVX1 U1378 ( .A(n1031), .Y(n1032) );
  AND2X2 U1379 ( .A(\mem<47><4> ), .B(n5728), .Y(n1033) );
  INVX1 U1380 ( .A(n1033), .Y(n1034) );
  AND2X2 U1381 ( .A(\mem<15><5> ), .B(n79), .Y(n1035) );
  INVX1 U1382 ( .A(n1035), .Y(n1036) );
  AND2X2 U1383 ( .A(n617), .B(\mem<39><5> ), .Y(n1037) );
  INVX1 U1384 ( .A(n1037), .Y(n1038) );
  AND2X2 U1385 ( .A(\mem<19><5> ), .B(n188), .Y(n1039) );
  INVX1 U1386 ( .A(n1039), .Y(n1040) );
  AND2X2 U1387 ( .A(\mem<23><5> ), .B(n79), .Y(n1041) );
  INVX1 U1388 ( .A(n1041), .Y(n1042) );
  AND2X2 U1389 ( .A(\mem<51><5> ), .B(n192), .Y(n1043) );
  INVX1 U1390 ( .A(n1043), .Y(n1044) );
  AND2X2 U1391 ( .A(\mem<55><5> ), .B(n77), .Y(n1045) );
  INVX1 U1392 ( .A(n1045), .Y(n1046) );
  AND2X2 U1393 ( .A(\mem<47><5> ), .B(n227), .Y(n1047) );
  INVX1 U1394 ( .A(n1047), .Y(n1048) );
  AND2X2 U1395 ( .A(\mem<11><6> ), .B(n202), .Y(n1049) );
  INVX1 U1396 ( .A(n1049), .Y(n1050) );
  AND2X2 U1397 ( .A(\mem<15><6> ), .B(n617), .Y(n1051) );
  INVX1 U1398 ( .A(n1051), .Y(n1052) );
  AND2X2 U1399 ( .A(\mem<35><6> ), .B(n198), .Y(n1053) );
  INVX1 U1400 ( .A(n1053), .Y(n1054) );
  AND2X2 U1401 ( .A(n77), .B(\mem<39><6> ), .Y(n1055) );
  INVX1 U1402 ( .A(n1055), .Y(n1056) );
  AND2X2 U1403 ( .A(\mem<19><6> ), .B(n169), .Y(n1057) );
  INVX1 U1404 ( .A(n1057), .Y(n1058) );
  AND2X2 U1405 ( .A(\mem<23><6> ), .B(n79), .Y(n1059) );
  INVX1 U1406 ( .A(n1059), .Y(n1060) );
  AND2X2 U1407 ( .A(\mem<55><6> ), .B(n77), .Y(n1061) );
  INVX1 U1408 ( .A(n1061), .Y(n1062) );
  AND2X2 U1409 ( .A(\mem<11><7> ), .B(n191), .Y(n1063) );
  INVX1 U1410 ( .A(n1063), .Y(n1064) );
  AND2X2 U1411 ( .A(n77), .B(\mem<15><7> ), .Y(n1065) );
  INVX1 U1412 ( .A(n1065), .Y(n1066) );
  AND2X2 U1413 ( .A(\mem<39><7> ), .B(n617), .Y(n1067) );
  INVX1 U1414 ( .A(n1067), .Y(n1068) );
  AND2X2 U1415 ( .A(\mem<19><7> ), .B(n190), .Y(n1069) );
  INVX1 U1416 ( .A(n1069), .Y(n1070) );
  AND2X2 U1417 ( .A(\mem<23><7> ), .B(n77), .Y(n1071) );
  INVX1 U1418 ( .A(n1071), .Y(n1072) );
  AND2X2 U1419 ( .A(\mem<55><7> ), .B(n77), .Y(n1073) );
  INVX1 U1420 ( .A(n1073), .Y(n1074) );
  AND2X2 U1421 ( .A(\mem<7><7> ), .B(n227), .Y(n1075) );
  INVX1 U1422 ( .A(n1075), .Y(n1076) );
  BUFX2 U1423 ( .A(n5913), .Y(n1077) );
  BUFX2 U1424 ( .A(n6067), .Y(n1078) );
  BUFX2 U1425 ( .A(n6216), .Y(n1079) );
  AND2X2 U1426 ( .A(n5604), .B(n3948), .Y(n1080) );
  INVX1 U1427 ( .A(n1080), .Y(n1081) );
  AND2X2 U1428 ( .A(n5185), .B(n5338), .Y(n1082) );
  INVX1 U1429 ( .A(n1082), .Y(n1083) );
  AND2X2 U1430 ( .A(n5311), .B(n3948), .Y(n1084) );
  INVX1 U1431 ( .A(n1084), .Y(n1085) );
  AND2X2 U1432 ( .A(n5302), .B(n5656), .Y(n1086) );
  INVX1 U1433 ( .A(n1086), .Y(n1087) );
  AND2X2 U1434 ( .A(n5395), .B(n5217), .Y(n1088) );
  INVX1 U1435 ( .A(n1088), .Y(n1089) );
  AND2X2 U1436 ( .A(n5656), .B(n5318), .Y(n1090) );
  INVX1 U1437 ( .A(n1090), .Y(n1091) );
  AND2X2 U1438 ( .A(n5646), .B(n5192), .Y(n1092) );
  INVX1 U1439 ( .A(n1092), .Y(n1093) );
  AND2X2 U1440 ( .A(n5657), .B(n5226), .Y(n1094) );
  INVX1 U1441 ( .A(n1094), .Y(n1095) );
  AND2X2 U1442 ( .A(n5185), .B(n5410), .Y(n1096) );
  INVX1 U1443 ( .A(n1096), .Y(n1097) );
  OR2X2 U1444 ( .A(n5930), .B(n5929), .Y(n1098) );
  INVX1 U1445 ( .A(n1098), .Y(n1099) );
  OR2X2 U1446 ( .A(n6086), .B(n6085), .Y(n1100) );
  INVX1 U1447 ( .A(n1100), .Y(n1101) );
  OR2X2 U1448 ( .A(n6237), .B(n6236), .Y(n1102) );
  INVX1 U1449 ( .A(n1102), .Y(n1103) );
  OR2X2 U1450 ( .A(n6317), .B(n6316), .Y(n1104) );
  INVX1 U1451 ( .A(n1104), .Y(n1105) );
  AND2X2 U1452 ( .A(\mem<57><7> ), .B(n5753), .Y(n1106) );
  INVX1 U1453 ( .A(n1106), .Y(n1107) );
  OR2X2 U1454 ( .A(n6396), .B(n6395), .Y(n1108) );
  INVX1 U1455 ( .A(n1108), .Y(n1109) );
  BUFX2 U1456 ( .A(n5914), .Y(n1110) );
  BUFX2 U1457 ( .A(n6068), .Y(n1111) );
  BUFX2 U1458 ( .A(n6217), .Y(n1112) );
  AND2X2 U1459 ( .A(n5388), .B(n5655), .Y(n1113) );
  INVX1 U1460 ( .A(n1113), .Y(n1114) );
  AND2X2 U1461 ( .A(n5700), .B(n92), .Y(n1115) );
  INVX1 U1462 ( .A(n1115), .Y(n1116) );
  AND2X2 U1463 ( .A(n3948), .B(n5287), .Y(n1117) );
  INVX1 U1464 ( .A(n1117), .Y(n1118) );
  AND2X2 U1465 ( .A(n653), .B(n652), .Y(n1119) );
  INVX1 U1466 ( .A(n1119), .Y(n1120) );
  OR2X2 U1467 ( .A(n5934), .B(n5933), .Y(n1121) );
  INVX1 U1468 ( .A(n1121), .Y(n1122) );
  OR2X2 U1469 ( .A(n6081), .B(n6080), .Y(n1123) );
  INVX1 U1470 ( .A(n1123), .Y(n1124) );
  OR2X2 U1471 ( .A(n6158), .B(n6157), .Y(n1125) );
  INVX1 U1472 ( .A(n1125), .Y(n1126) );
  OR2X2 U1473 ( .A(n6232), .B(n6231), .Y(n1127) );
  INVX1 U1474 ( .A(n1127), .Y(n1128) );
  OR2X2 U1475 ( .A(n6311), .B(n6310), .Y(n1129) );
  INVX1 U1476 ( .A(n1129), .Y(n1130) );
  OR2X2 U1477 ( .A(n6390), .B(n6389), .Y(n1131) );
  INVX1 U1478 ( .A(n1131), .Y(n1132) );
  AND2X2 U1479 ( .A(n5763), .B(n5762), .Y(n1133) );
  INVX1 U1480 ( .A(n1133), .Y(n1134) );
  BUFX2 U1481 ( .A(n6143), .Y(n1135) );
  AND2X2 U1482 ( .A(n65), .B(N181), .Y(n1136) );
  INVX1 U1483 ( .A(n1136), .Y(n1137) );
  AND2X2 U1484 ( .A(n905), .B(n942), .Y(n1138) );
  INVX1 U1485 ( .A(n1138), .Y(n1139) );
  BUFX2 U1486 ( .A(n5775), .Y(n1140) );
  AND2X2 U1487 ( .A(n5707), .B(n4173), .Y(n1141) );
  INVX1 U1488 ( .A(n1141), .Y(n1142) );
  INVX1 U1489 ( .A(n3763), .Y(n1143) );
  AND2X2 U1490 ( .A(n5770), .B(n5769), .Y(n1144) );
  INVX1 U1491 ( .A(n1144), .Y(n1145) );
  BUFX2 U1492 ( .A(n5829), .Y(n1146) );
  BUFX2 U1493 ( .A(n5993), .Y(n1147) );
  BUFX2 U1494 ( .A(n6293), .Y(n1148) );
  BUFX2 U1495 ( .A(n6373), .Y(n1149) );
  AND2X2 U1496 ( .A(n917), .B(n76), .Y(n1150) );
  INVX1 U1497 ( .A(n1150), .Y(n1151) );
  OR2X2 U1498 ( .A(\addr<10> ), .B(\addr<14> ), .Y(n1152) );
  AND2X2 U1499 ( .A(\data_in<0> ), .B(n1543), .Y(n1153) );
  INVX1 U1500 ( .A(n1153), .Y(n1154) );
  AND2X2 U1501 ( .A(\data_in<1> ), .B(n1543), .Y(n1155) );
  INVX1 U1502 ( .A(n1155), .Y(n1156) );
  AND2X2 U1503 ( .A(\data_in<2> ), .B(n1543), .Y(n1157) );
  INVX1 U1504 ( .A(n1157), .Y(n1158) );
  AND2X2 U1505 ( .A(\data_in<3> ), .B(n1543), .Y(n1159) );
  INVX1 U1506 ( .A(n1159), .Y(n1160) );
  AND2X2 U1507 ( .A(\data_in<4> ), .B(n1543), .Y(n1161) );
  INVX1 U1508 ( .A(n1161), .Y(n1162) );
  AND2X2 U1509 ( .A(\data_in<5> ), .B(n1543), .Y(n1163) );
  INVX1 U1510 ( .A(n1163), .Y(n1164) );
  AND2X2 U1511 ( .A(\data_in<6> ), .B(n1543), .Y(n1165) );
  INVX1 U1512 ( .A(n1165), .Y(n1166) );
  AND2X2 U1513 ( .A(\data_in<7> ), .B(n1543), .Y(n1167) );
  INVX1 U1514 ( .A(n1167), .Y(n1168) );
  AND2X2 U1515 ( .A(\data_in<8> ), .B(n43), .Y(n1169) );
  INVX1 U1516 ( .A(n1169), .Y(n1170) );
  AND2X2 U1517 ( .A(\data_in<9> ), .B(n1552), .Y(n1171) );
  INVX1 U1518 ( .A(n1171), .Y(n1172) );
  AND2X2 U1519 ( .A(\data_in<2> ), .B(n1551), .Y(n1173) );
  INVX1 U1520 ( .A(n1173), .Y(n1174) );
  AND2X2 U1521 ( .A(\data_in<11> ), .B(n1552), .Y(n1175) );
  INVX1 U1522 ( .A(n1175), .Y(n1176) );
  AND2X2 U1523 ( .A(\data_in<12> ), .B(n43), .Y(n1177) );
  INVX1 U1524 ( .A(n1177), .Y(n1178) );
  AND2X2 U1525 ( .A(\data_in<5> ), .B(n1551), .Y(n1179) );
  INVX1 U1526 ( .A(n1179), .Y(n1180) );
  AND2X2 U1527 ( .A(\data_in<14> ), .B(n43), .Y(n1181) );
  INVX1 U1528 ( .A(n1181), .Y(n1182) );
  AND2X2 U1529 ( .A(\data_in<15> ), .B(n1552), .Y(n1183) );
  INVX1 U1530 ( .A(n1183), .Y(n1184) );
  AND2X2 U1531 ( .A(\data_in<7> ), .B(n1553), .Y(n1185) );
  INVX1 U1532 ( .A(n1185), .Y(n1186) );
  AND2X2 U1533 ( .A(\data_in<0> ), .B(n1560), .Y(n1187) );
  INVX1 U1534 ( .A(n1187), .Y(n1188) );
  AND2X2 U1535 ( .A(\data_in<1> ), .B(n53), .Y(n1189) );
  INVX1 U1536 ( .A(n1189), .Y(n1190) );
  AND2X2 U1537 ( .A(\data_in<2> ), .B(n1560), .Y(n1191) );
  INVX1 U1538 ( .A(n1191), .Y(n1192) );
  AND2X2 U1539 ( .A(\data_in<3> ), .B(n53), .Y(n1193) );
  INVX1 U1540 ( .A(n1193), .Y(n1194) );
  AND2X2 U1541 ( .A(\data_in<4> ), .B(n1560), .Y(n1195) );
  INVX1 U1542 ( .A(n1195), .Y(n1196) );
  AND2X2 U1543 ( .A(\data_in<5> ), .B(n53), .Y(n1197) );
  INVX1 U1544 ( .A(n1197), .Y(n1198) );
  AND2X2 U1545 ( .A(\data_in<6> ), .B(n1560), .Y(n1199) );
  INVX1 U1546 ( .A(n1199), .Y(n1200) );
  AND2X2 U1547 ( .A(\data_in<7> ), .B(n53), .Y(n1201) );
  INVX1 U1548 ( .A(n1201), .Y(n1202) );
  AND2X2 U1549 ( .A(\data_in<0> ), .B(n1562), .Y(n1203) );
  INVX1 U1550 ( .A(n1203), .Y(n1204) );
  AND2X2 U1551 ( .A(\data_in<1> ), .B(n52), .Y(n1205) );
  INVX1 U1552 ( .A(n1205), .Y(n1206) );
  AND2X2 U1553 ( .A(\data_in<2> ), .B(n52), .Y(n1207) );
  INVX1 U1554 ( .A(n1207), .Y(n1208) );
  AND2X2 U1555 ( .A(\data_in<3> ), .B(n1562), .Y(n1209) );
  INVX1 U1556 ( .A(n1209), .Y(n1210) );
  AND2X2 U1557 ( .A(\data_in<4> ), .B(n52), .Y(n1211) );
  INVX1 U1558 ( .A(n1211), .Y(n1212) );
  AND2X2 U1559 ( .A(\data_in<5> ), .B(n1562), .Y(n1213) );
  INVX1 U1560 ( .A(n1213), .Y(n1214) );
  AND2X2 U1561 ( .A(\data_in<6> ), .B(n52), .Y(n1215) );
  INVX1 U1562 ( .A(n1215), .Y(n1216) );
  AND2X2 U1563 ( .A(\data_in<7> ), .B(n1562), .Y(n1217) );
  INVX1 U1564 ( .A(n1217), .Y(n1218) );
  AND2X2 U1565 ( .A(\data_in<0> ), .B(n1564), .Y(n1219) );
  INVX1 U1566 ( .A(n1219), .Y(n1220) );
  AND2X2 U1567 ( .A(\data_in<1> ), .B(n1564), .Y(n1221) );
  INVX1 U1568 ( .A(n1221), .Y(n1222) );
  AND2X2 U1569 ( .A(\data_in<2> ), .B(n1564), .Y(n1223) );
  INVX1 U1570 ( .A(n1223), .Y(n1224) );
  AND2X2 U1571 ( .A(\data_in<3> ), .B(n1564), .Y(n1225) );
  INVX1 U1572 ( .A(n1225), .Y(n1226) );
  AND2X2 U1573 ( .A(\data_in<4> ), .B(n1564), .Y(n1227) );
  INVX1 U1574 ( .A(n1227), .Y(n1228) );
  AND2X2 U1575 ( .A(\data_in<5> ), .B(n1564), .Y(n1229) );
  INVX1 U1576 ( .A(n1229), .Y(n1230) );
  AND2X2 U1577 ( .A(\data_in<6> ), .B(n1564), .Y(n1231) );
  INVX1 U1578 ( .A(n1231), .Y(n1232) );
  AND2X2 U1579 ( .A(\data_in<7> ), .B(n1564), .Y(n1233) );
  INVX1 U1580 ( .A(n1233), .Y(n1234) );
  AND2X2 U1581 ( .A(n51), .B(\data_in<0> ), .Y(n1235) );
  INVX1 U1582 ( .A(n1235), .Y(n1236) );
  AND2X2 U1583 ( .A(n51), .B(\data_in<1> ), .Y(n1237) );
  INVX1 U1584 ( .A(n1237), .Y(n1238) );
  AND2X2 U1585 ( .A(\data_in<2> ), .B(n1566), .Y(n1239) );
  INVX1 U1586 ( .A(n1239), .Y(n1240) );
  AND2X2 U1587 ( .A(n51), .B(\data_in<3> ), .Y(n1241) );
  INVX1 U1588 ( .A(n1241), .Y(n1242) );
  AND2X2 U1589 ( .A(\data_in<4> ), .B(n1566), .Y(n1243) );
  INVX1 U1590 ( .A(n1243), .Y(n1244) );
  AND2X2 U1591 ( .A(\data_in<5> ), .B(n1566), .Y(n1245) );
  INVX1 U1592 ( .A(n1245), .Y(n1246) );
  AND2X2 U1593 ( .A(\data_in<6> ), .B(n1566), .Y(n1247) );
  INVX1 U1594 ( .A(n1247), .Y(n1248) );
  AND2X2 U1595 ( .A(\data_in<7> ), .B(n51), .Y(n1249) );
  INVX1 U1596 ( .A(n1249), .Y(n1250) );
  AND2X2 U1597 ( .A(\data_in<0> ), .B(n1568), .Y(n1251) );
  INVX1 U1598 ( .A(n1251), .Y(n1252) );
  AND2X2 U1599 ( .A(\data_in<1> ), .B(n1568), .Y(n1253) );
  INVX1 U1600 ( .A(n1253), .Y(n1254) );
  AND2X2 U1601 ( .A(\data_in<2> ), .B(n1568), .Y(n1255) );
  INVX1 U1602 ( .A(n1255), .Y(n1256) );
  AND2X2 U1603 ( .A(\data_in<3> ), .B(n1568), .Y(n1257) );
  INVX1 U1604 ( .A(n1257), .Y(n1258) );
  AND2X2 U1605 ( .A(\data_in<4> ), .B(n1568), .Y(n1259) );
  INVX1 U1606 ( .A(n1259), .Y(n1260) );
  AND2X2 U1607 ( .A(\data_in<5> ), .B(n1568), .Y(n1261) );
  INVX1 U1608 ( .A(n1261), .Y(n1262) );
  AND2X2 U1609 ( .A(\data_in<6> ), .B(n1568), .Y(n1263) );
  INVX1 U1610 ( .A(n1263), .Y(n1264) );
  AND2X2 U1611 ( .A(\data_in<7> ), .B(n1568), .Y(n1265) );
  INVX1 U1612 ( .A(n1265), .Y(n1266) );
  AND2X2 U1613 ( .A(\data_in<0> ), .B(n1570), .Y(n1267) );
  INVX1 U1614 ( .A(n1267), .Y(n1268) );
  AND2X2 U1615 ( .A(\data_in<1> ), .B(n12), .Y(n1269) );
  INVX1 U1616 ( .A(n1269), .Y(n1270) );
  AND2X2 U1617 ( .A(\data_in<2> ), .B(n1570), .Y(n1271) );
  INVX1 U1618 ( .A(n1271), .Y(n1272) );
  AND2X2 U1619 ( .A(\data_in<3> ), .B(n12), .Y(n1273) );
  INVX1 U1620 ( .A(n1273), .Y(n1274) );
  AND2X2 U1621 ( .A(\data_in<4> ), .B(n12), .Y(n1275) );
  INVX1 U1622 ( .A(n1275), .Y(n1276) );
  AND2X2 U1623 ( .A(\data_in<5> ), .B(n1570), .Y(n1277) );
  INVX1 U1624 ( .A(n1277), .Y(n1278) );
  AND2X2 U1625 ( .A(\data_in<6> ), .B(n12), .Y(n1279) );
  INVX1 U1626 ( .A(n1279), .Y(n1280) );
  AND2X2 U1627 ( .A(\data_in<7> ), .B(n1570), .Y(n1281) );
  INVX1 U1628 ( .A(n1281), .Y(n1282) );
  AND2X2 U1629 ( .A(\data_in<0> ), .B(n1572), .Y(n1283) );
  INVX1 U1630 ( .A(n1283), .Y(n1284) );
  AND2X2 U1631 ( .A(\data_in<1> ), .B(n1572), .Y(n1285) );
  INVX1 U1632 ( .A(n1285), .Y(n1286) );
  AND2X2 U1633 ( .A(\data_in<2> ), .B(n1572), .Y(n1287) );
  INVX1 U1634 ( .A(n1287), .Y(n1288) );
  AND2X2 U1635 ( .A(\data_in<3> ), .B(n1572), .Y(n1289) );
  INVX1 U1636 ( .A(n1289), .Y(n1290) );
  AND2X2 U1637 ( .A(\data_in<4> ), .B(n1572), .Y(n1291) );
  INVX1 U1638 ( .A(n1291), .Y(n1292) );
  AND2X2 U1639 ( .A(\data_in<5> ), .B(n1572), .Y(n1293) );
  INVX1 U1640 ( .A(n1293), .Y(n1294) );
  AND2X2 U1641 ( .A(\data_in<6> ), .B(n1572), .Y(n1295) );
  INVX1 U1642 ( .A(n1295), .Y(n1296) );
  AND2X2 U1643 ( .A(\data_in<7> ), .B(n1572), .Y(n1297) );
  INVX1 U1644 ( .A(n1297), .Y(n1298) );
  AND2X2 U1645 ( .A(\data_in<2> ), .B(n49), .Y(n1299) );
  INVX1 U1646 ( .A(n1299), .Y(n1300) );
  AND2X2 U1647 ( .A(\data_in<5> ), .B(n49), .Y(n1301) );
  INVX1 U1648 ( .A(n1301), .Y(n1302) );
  AND2X2 U1649 ( .A(\data_in<0> ), .B(n1580), .Y(n1303) );
  INVX1 U1650 ( .A(n1303), .Y(n1304) );
  AND2X2 U1651 ( .A(\data_in<1> ), .B(n1580), .Y(n1305) );
  INVX1 U1652 ( .A(n1305), .Y(n1306) );
  AND2X2 U1653 ( .A(\data_in<3> ), .B(n1580), .Y(n1307) );
  INVX1 U1654 ( .A(n1307), .Y(n1308) );
  AND2X2 U1655 ( .A(\data_in<4> ), .B(n1580), .Y(n1309) );
  INVX1 U1656 ( .A(n1309), .Y(n1310) );
  AND2X2 U1657 ( .A(\data_in<6> ), .B(n1580), .Y(n1311) );
  INVX1 U1658 ( .A(n1311), .Y(n1312) );
  AND2X2 U1659 ( .A(\data_in<7> ), .B(n1580), .Y(n1313) );
  INVX1 U1660 ( .A(n1313), .Y(n1314) );
  AND2X2 U1661 ( .A(\data_in<0> ), .B(n1582), .Y(n1315) );
  INVX1 U1662 ( .A(n1315), .Y(n1316) );
  AND2X2 U1663 ( .A(\data_in<1> ), .B(n1582), .Y(n1317) );
  INVX1 U1664 ( .A(n1317), .Y(n1318) );
  AND2X2 U1665 ( .A(\data_in<2> ), .B(n1582), .Y(n1319) );
  INVX1 U1666 ( .A(n1319), .Y(n1320) );
  AND2X2 U1667 ( .A(\data_in<3> ), .B(n1582), .Y(n1321) );
  INVX1 U1668 ( .A(n1321), .Y(n1322) );
  AND2X2 U1669 ( .A(\data_in<4> ), .B(n1582), .Y(n1323) );
  INVX1 U1670 ( .A(n1323), .Y(n1324) );
  AND2X2 U1671 ( .A(\data_in<5> ), .B(n1582), .Y(n1325) );
  INVX1 U1672 ( .A(n1325), .Y(n1326) );
  AND2X2 U1673 ( .A(\data_in<6> ), .B(n1582), .Y(n1327) );
  INVX1 U1674 ( .A(n1327), .Y(n1328) );
  AND2X2 U1675 ( .A(\data_in<7> ), .B(n1582), .Y(n1329) );
  INVX1 U1676 ( .A(n1329), .Y(n1330) );
  AND2X2 U1677 ( .A(\data_in<0> ), .B(n48), .Y(n1331) );
  INVX1 U1678 ( .A(n1331), .Y(n1332) );
  AND2X2 U1679 ( .A(\data_in<1> ), .B(n1584), .Y(n1333) );
  INVX1 U1680 ( .A(n1333), .Y(n1334) );
  AND2X2 U1681 ( .A(\data_in<2> ), .B(n48), .Y(n1335) );
  INVX1 U1682 ( .A(n1335), .Y(n1336) );
  AND2X2 U1683 ( .A(\data_in<3> ), .B(n1584), .Y(n1337) );
  INVX1 U1684 ( .A(n1337), .Y(n1338) );
  AND2X2 U1685 ( .A(\data_in<4> ), .B(n48), .Y(n1339) );
  INVX1 U1686 ( .A(n1339), .Y(n1340) );
  AND2X2 U1687 ( .A(\data_in<5> ), .B(n1584), .Y(n1341) );
  INVX1 U1688 ( .A(n1341), .Y(n1342) );
  AND2X2 U1689 ( .A(\data_in<6> ), .B(n48), .Y(n1343) );
  INVX1 U1690 ( .A(n1343), .Y(n1344) );
  AND2X2 U1691 ( .A(\data_in<7> ), .B(n1584), .Y(n1345) );
  INVX1 U1692 ( .A(n1345), .Y(n1346) );
  AND2X2 U1693 ( .A(\data_in<7> ), .B(n1588), .Y(n1347) );
  INVX1 U1694 ( .A(n1347), .Y(n1348) );
  AND2X2 U1695 ( .A(\data_in<8> ), .B(n1605), .Y(n1349) );
  INVX1 U1696 ( .A(n1349), .Y(n1350) );
  AND2X2 U1697 ( .A(\data_in<9> ), .B(n1605), .Y(n1351) );
  INVX1 U1698 ( .A(n1351), .Y(n1352) );
  AND2X2 U1699 ( .A(\data_in<10> ), .B(n21), .Y(n1353) );
  INVX1 U1700 ( .A(n1353), .Y(n1354) );
  AND2X2 U1701 ( .A(\data_in<11> ), .B(n21), .Y(n1355) );
  INVX1 U1702 ( .A(n1355), .Y(n1356) );
  AND2X2 U1703 ( .A(\data_in<12> ), .B(n1605), .Y(n1357) );
  INVX1 U1704 ( .A(n1357), .Y(n1358) );
  AND2X2 U1705 ( .A(\data_in<13> ), .B(n1605), .Y(n1359) );
  INVX1 U1706 ( .A(n1359), .Y(n1360) );
  AND2X2 U1707 ( .A(\data_in<14> ), .B(n21), .Y(n1361) );
  INVX1 U1708 ( .A(n1361), .Y(n1362) );
  AND2X2 U1709 ( .A(\data_in<15> ), .B(n21), .Y(n1363) );
  INVX1 U1710 ( .A(n1363), .Y(n1364) );
  AND2X2 U1711 ( .A(\mem<16><2> ), .B(n5052), .Y(n1365) );
  INVX1 U1712 ( .A(n1365), .Y(n1366) );
  AND2X2 U1713 ( .A(\mem<16><5> ), .B(n5052), .Y(n1367) );
  INVX1 U1714 ( .A(n1367), .Y(n1368) );
  AND2X2 U1715 ( .A(\data_in<0> ), .B(n18), .Y(n1369) );
  INVX1 U1716 ( .A(n1369), .Y(n1370) );
  AND2X2 U1717 ( .A(\data_in<1> ), .B(n1621), .Y(n1371) );
  INVX1 U1718 ( .A(n1371), .Y(n1372) );
  AND2X2 U1719 ( .A(\data_in<2> ), .B(n1621), .Y(n1373) );
  INVX1 U1720 ( .A(n1373), .Y(n1374) );
  AND2X2 U1721 ( .A(\data_in<3> ), .B(n18), .Y(n1375) );
  INVX1 U1722 ( .A(n1375), .Y(n1376) );
  AND2X2 U1723 ( .A(\data_in<4> ), .B(n18), .Y(n1377) );
  INVX1 U1724 ( .A(n1377), .Y(n1378) );
  AND2X2 U1725 ( .A(\data_in<5> ), .B(n1621), .Y(n1379) );
  INVX1 U1726 ( .A(n1379), .Y(n1380) );
  AND2X2 U1727 ( .A(\data_in<6> ), .B(n1621), .Y(n1381) );
  INVX1 U1728 ( .A(n1381), .Y(n1382) );
  AND2X2 U1729 ( .A(\data_in<7> ), .B(n18), .Y(n1383) );
  INVX1 U1730 ( .A(n1383), .Y(n1384) );
  AND2X2 U1731 ( .A(\data_in<0> ), .B(n1630), .Y(n1385) );
  INVX1 U1732 ( .A(n1385), .Y(n1386) );
  AND2X2 U1733 ( .A(\data_in<1> ), .B(n1630), .Y(n1387) );
  INVX1 U1734 ( .A(n1387), .Y(n1388) );
  AND2X2 U1735 ( .A(\data_in<2> ), .B(n1630), .Y(n1389) );
  INVX1 U1736 ( .A(n1389), .Y(n1390) );
  AND2X2 U1737 ( .A(\data_in<3> ), .B(n1630), .Y(n1391) );
  INVX1 U1738 ( .A(n1391), .Y(n1392) );
  AND2X2 U1739 ( .A(\data_in<4> ), .B(n1630), .Y(n1393) );
  INVX1 U1740 ( .A(n1393), .Y(n1394) );
  AND2X2 U1741 ( .A(\data_in<5> ), .B(n1630), .Y(n1395) );
  INVX1 U1742 ( .A(n1395), .Y(n1396) );
  AND2X2 U1743 ( .A(\data_in<6> ), .B(n1630), .Y(n1397) );
  INVX1 U1744 ( .A(n1397), .Y(n1398) );
  AND2X2 U1745 ( .A(\data_in<7> ), .B(n1630), .Y(n1399) );
  INVX1 U1746 ( .A(n1399), .Y(n1400) );
  AND2X2 U1747 ( .A(\data_in<8> ), .B(n4209), .Y(n1401) );
  INVX1 U1748 ( .A(n1401), .Y(n1402) );
  AND2X2 U1749 ( .A(\data_in<9> ), .B(n4209), .Y(n1403) );
  INVX1 U1750 ( .A(n1403), .Y(n1404) );
  AND2X2 U1751 ( .A(\data_in<10> ), .B(n4209), .Y(n1405) );
  INVX1 U1752 ( .A(n1405), .Y(n1406) );
  AND2X2 U1753 ( .A(\data_in<11> ), .B(n4209), .Y(n1407) );
  INVX1 U1754 ( .A(n1407), .Y(n1408) );
  AND2X2 U1755 ( .A(\data_in<12> ), .B(n4209), .Y(n1409) );
  INVX1 U1756 ( .A(n1409), .Y(n1410) );
  AND2X2 U1757 ( .A(\data_in<13> ), .B(n4209), .Y(n1411) );
  INVX1 U1758 ( .A(n1411), .Y(n1412) );
  AND2X2 U1759 ( .A(\data_in<14> ), .B(n4209), .Y(n1413) );
  INVX1 U1760 ( .A(n1413), .Y(n1414) );
  AND2X2 U1761 ( .A(\data_in<15> ), .B(n4209), .Y(n1415) );
  INVX1 U1762 ( .A(n1415), .Y(n1416) );
  AND2X2 U1763 ( .A(\data_in<8> ), .B(n1636), .Y(n1417) );
  INVX1 U1764 ( .A(n1417), .Y(n1418) );
  AND2X2 U1765 ( .A(\data_in<9> ), .B(n1636), .Y(n1419) );
  INVX1 U1766 ( .A(n1419), .Y(n1420) );
  AND2X2 U1767 ( .A(\data_in<10> ), .B(n1636), .Y(n1421) );
  INVX1 U1768 ( .A(n1421), .Y(n1422) );
  AND2X2 U1769 ( .A(\data_in<11> ), .B(n1636), .Y(n1423) );
  INVX1 U1770 ( .A(n1423), .Y(n1424) );
  AND2X2 U1771 ( .A(\data_in<12> ), .B(n11), .Y(n1425) );
  INVX1 U1772 ( .A(n1425), .Y(n1426) );
  AND2X2 U1773 ( .A(\data_in<13> ), .B(n11), .Y(n1427) );
  INVX1 U1774 ( .A(n1427), .Y(n1428) );
  AND2X2 U1775 ( .A(\data_in<14> ), .B(n11), .Y(n1429) );
  INVX1 U1776 ( .A(n1429), .Y(n1430) );
  AND2X2 U1777 ( .A(\data_in<15> ), .B(n11), .Y(n1431) );
  INVX1 U1778 ( .A(n1431), .Y(n1432) );
  AND2X2 U1779 ( .A(\data_in<0> ), .B(n1637), .Y(n1433) );
  INVX1 U1780 ( .A(n1433), .Y(n1434) );
  AND2X2 U1781 ( .A(\data_in<1> ), .B(n1637), .Y(n1435) );
  INVX1 U1782 ( .A(n1435), .Y(n1436) );
  AND2X2 U1783 ( .A(\data_in<2> ), .B(n1637), .Y(n1437) );
  INVX1 U1784 ( .A(n1437), .Y(n1438) );
  AND2X2 U1785 ( .A(\data_in<3> ), .B(n1637), .Y(n1439) );
  INVX1 U1786 ( .A(n1439), .Y(n1440) );
  AND2X2 U1787 ( .A(\data_in<4> ), .B(n1637), .Y(n1441) );
  INVX1 U1788 ( .A(n1441), .Y(n1442) );
  AND2X2 U1789 ( .A(\data_in<5> ), .B(n1637), .Y(n1443) );
  INVX1 U1790 ( .A(n1443), .Y(n1444) );
  AND2X2 U1791 ( .A(\data_in<6> ), .B(n1637), .Y(n1445) );
  INVX1 U1792 ( .A(n1445), .Y(n1446) );
  AND2X2 U1793 ( .A(\data_in<7> ), .B(n1637), .Y(n1447) );
  INVX1 U1794 ( .A(n1447), .Y(n1448) );
  AND2X2 U1795 ( .A(\data_in<0> ), .B(n1639), .Y(n1449) );
  INVX1 U1796 ( .A(n1449), .Y(n1450) );
  AND2X2 U1797 ( .A(\data_in<1> ), .B(n1639), .Y(n1451) );
  INVX1 U1798 ( .A(n1451), .Y(n1452) );
  AND2X2 U1799 ( .A(\data_in<2> ), .B(n1639), .Y(n1453) );
  INVX1 U1800 ( .A(n1453), .Y(n1454) );
  AND2X2 U1801 ( .A(\data_in<3> ), .B(n1639), .Y(n1455) );
  INVX1 U1802 ( .A(n1455), .Y(n1456) );
  AND2X2 U1803 ( .A(\data_in<4> ), .B(n1639), .Y(n1457) );
  INVX1 U1804 ( .A(n1457), .Y(n1458) );
  AND2X2 U1805 ( .A(\data_in<5> ), .B(n1639), .Y(n1459) );
  INVX1 U1806 ( .A(n1459), .Y(n1460) );
  AND2X2 U1807 ( .A(\data_in<6> ), .B(n1639), .Y(n1461) );
  INVX1 U1808 ( .A(n1461), .Y(n1462) );
  AND2X2 U1809 ( .A(\data_in<7> ), .B(n1639), .Y(n1463) );
  INVX1 U1810 ( .A(n1463), .Y(n1464) );
  AND2X2 U1811 ( .A(\data_in<0> ), .B(n1641), .Y(n1465) );
  INVX1 U1812 ( .A(n1465), .Y(n1466) );
  AND2X2 U1813 ( .A(\data_in<1> ), .B(n1641), .Y(n1467) );
  INVX1 U1814 ( .A(n1467), .Y(n1468) );
  AND2X2 U1815 ( .A(\data_in<10> ), .B(n1642), .Y(n1469) );
  INVX1 U1816 ( .A(n1469), .Y(n1470) );
  AND2X2 U1817 ( .A(\data_in<3> ), .B(n1641), .Y(n1471) );
  INVX1 U1818 ( .A(n1471), .Y(n1472) );
  AND2X2 U1819 ( .A(\data_in<4> ), .B(n1641), .Y(n1473) );
  INVX1 U1820 ( .A(n1473), .Y(n1474) );
  AND2X2 U1821 ( .A(\data_in<13> ), .B(n1642), .Y(n1475) );
  INVX1 U1822 ( .A(n1475), .Y(n1476) );
  AND2X2 U1823 ( .A(\data_in<6> ), .B(n1641), .Y(n1477) );
  INVX1 U1824 ( .A(n1477), .Y(n1478) );
  AND2X2 U1825 ( .A(\data_in<7> ), .B(n1641), .Y(n1479) );
  INVX1 U1826 ( .A(n1479), .Y(n1480) );
  AND2X2 U1827 ( .A(\data_in<0> ), .B(n1643), .Y(n1481) );
  INVX1 U1828 ( .A(n1481), .Y(n1482) );
  AND2X2 U1829 ( .A(\data_in<1> ), .B(n1643), .Y(n1483) );
  INVX1 U1830 ( .A(n1483), .Y(n1484) );
  AND2X2 U1831 ( .A(\data_in<2> ), .B(n1643), .Y(n1485) );
  INVX1 U1832 ( .A(n1485), .Y(n1486) );
  AND2X2 U1833 ( .A(\data_in<3> ), .B(n1643), .Y(n1487) );
  INVX1 U1834 ( .A(n1487), .Y(n1488) );
  AND2X2 U1835 ( .A(\data_in<4> ), .B(n1643), .Y(n1489) );
  INVX1 U1836 ( .A(n1489), .Y(n1490) );
  AND2X2 U1837 ( .A(\data_in<5> ), .B(n1643), .Y(n1491) );
  INVX1 U1838 ( .A(n1491), .Y(n1492) );
  AND2X2 U1839 ( .A(\data_in<14> ), .B(n1644), .Y(n1493) );
  INVX1 U1840 ( .A(n1493), .Y(n1494) );
  AND2X2 U1841 ( .A(\data_in<15> ), .B(n1644), .Y(n1495) );
  INVX1 U1842 ( .A(n1495), .Y(n1496) );
  AND2X2 U1843 ( .A(\data_in<0> ), .B(n1645), .Y(n1497) );
  INVX1 U1844 ( .A(n1497), .Y(n1498) );
  AND2X2 U1845 ( .A(\data_in<1> ), .B(n1645), .Y(n1499) );
  INVX1 U1846 ( .A(n1499), .Y(n1500) );
  AND2X2 U1847 ( .A(\data_in<10> ), .B(n1646), .Y(n1501) );
  INVX1 U1848 ( .A(n1501), .Y(n1502) );
  AND2X2 U1849 ( .A(\data_in<3> ), .B(n1645), .Y(n1503) );
  INVX1 U1850 ( .A(n1503), .Y(n1504) );
  AND2X2 U1851 ( .A(\data_in<4> ), .B(n1645), .Y(n1505) );
  INVX1 U1852 ( .A(n1505), .Y(n1506) );
  AND2X2 U1853 ( .A(\data_in<13> ), .B(n1646), .Y(n1507) );
  INVX1 U1854 ( .A(n1507), .Y(n1508) );
  AND2X2 U1855 ( .A(\data_in<6> ), .B(n1645), .Y(n1509) );
  INVX1 U1856 ( .A(n1509), .Y(n1510) );
  AND2X2 U1857 ( .A(\data_in<7> ), .B(n1645), .Y(n1511) );
  INVX1 U1858 ( .A(n1511), .Y(n1512) );
  AND2X2 U1859 ( .A(\mem<1><0> ), .B(n6460), .Y(n1513) );
  INVX1 U1860 ( .A(n1513), .Y(n1514) );
  AND2X2 U1861 ( .A(\mem<1><1> ), .B(n6460), .Y(n1515) );
  INVX1 U1862 ( .A(n1515), .Y(n1516) );
  AND2X2 U1863 ( .A(\mem<1><2> ), .B(n6460), .Y(n1517) );
  INVX1 U1864 ( .A(n1517), .Y(n1518) );
  AND2X2 U1865 ( .A(\mem<1><3> ), .B(n6460), .Y(n1519) );
  INVX1 U1866 ( .A(n1519), .Y(n1520) );
  AND2X2 U1867 ( .A(\mem<1><4> ), .B(n6460), .Y(n1521) );
  INVX1 U1868 ( .A(n1521), .Y(n1522) );
  AND2X2 U1869 ( .A(\mem<1><5> ), .B(n6460), .Y(n1523) );
  INVX1 U1870 ( .A(n1523), .Y(n1524) );
  AND2X2 U1871 ( .A(\mem<1><6> ), .B(n6460), .Y(n1525) );
  INVX1 U1872 ( .A(n1525), .Y(n1526) );
  AND2X2 U1873 ( .A(\mem<1><7> ), .B(n6460), .Y(n1527) );
  INVX1 U1874 ( .A(n1527), .Y(n1528) );
  AND2X2 U1875 ( .A(n226), .B(n666), .Y(n1529) );
  AND2X2 U1876 ( .A(n220), .B(n666), .Y(n1530) );
  AND2X2 U1877 ( .A(n5732), .B(n667), .Y(n1531) );
  AND2X2 U1878 ( .A(n5735), .B(n667), .Y(n1532) );
  AND2X2 U1879 ( .A(n233), .B(n668), .Y(n1533) );
  AND2X2 U1880 ( .A(n5740), .B(n668), .Y(n1534) );
  AND2X2 U1881 ( .A(n154), .B(n669), .Y(n1535) );
  AND2X2 U1882 ( .A(n139), .B(n669), .Y(n1536) );
  AND2X2 U1883 ( .A(n201), .B(n670), .Y(n1537) );
  AND2X2 U1884 ( .A(n5747), .B(n670), .Y(n1538) );
  AND2X2 U1885 ( .A(n5141), .B(n671), .Y(n1539) );
  AND2X2 U1886 ( .A(n5118), .B(n671), .Y(n1540) );
  AND2X2 U1887 ( .A(n3928), .B(n6), .Y(n1542) );
  AND2X2 U1888 ( .A(n673), .B(n5726), .Y(n1543) );
  AND2X2 U1889 ( .A(n3667), .B(n673), .Y(n1544) );
  AND2X2 U1890 ( .A(n5729), .B(n675), .Y(n1545) );
  AND2X2 U1891 ( .A(n219), .B(n675), .Y(n1546) );
  AND2X2 U1892 ( .A(n5732), .B(n676), .Y(n1547) );
  AND2X2 U1893 ( .A(n5735), .B(n676), .Y(n1548) );
  AND2X2 U1894 ( .A(n5187), .B(n677), .Y(n1549) );
  AND2X2 U1895 ( .A(n5740), .B(n677), .Y(n1550) );
  AND2X2 U1896 ( .A(n678), .B(n155), .Y(n1551) );
  AND2X2 U1897 ( .A(n678), .B(n133), .Y(n1552) );
  AND2X2 U1898 ( .A(n196), .B(n691), .Y(n1553) );
  AND2X2 U1899 ( .A(n171), .B(n691), .Y(n1554) );
  AND2X2 U1900 ( .A(n5120), .B(n692), .Y(n1555) );
  AND2X2 U1901 ( .A(n5115), .B(n692), .Y(n1556) );
  AND2X2 U1902 ( .A(n92), .B(n693), .Y(n1557) );
  AND2X2 U1903 ( .A(n5751), .B(n693), .Y(n1558) );
  AND2X2 U1904 ( .A(n695), .B(n5099), .Y(n1559) );
  AND2X2 U1905 ( .A(n223), .B(n696), .Y(n1560) );
  AND2X2 U1906 ( .A(n222), .B(n696), .Y(n1561) );
  AND2X2 U1907 ( .A(n5732), .B(n713), .Y(n1562) );
  AND2X2 U1908 ( .A(n5735), .B(n713), .Y(n1563) );
  AND2X2 U1909 ( .A(n233), .B(n728), .Y(n1564) );
  AND2X2 U1910 ( .A(n5740), .B(n728), .Y(n1565) );
  AND2X2 U1911 ( .A(n162), .B(n740), .Y(n1566) );
  AND2X2 U1912 ( .A(n131), .B(n740), .Y(n1567) );
  AND2X2 U1913 ( .A(n197), .B(n752), .Y(n1568) );
  AND2X2 U1914 ( .A(n5747), .B(n752), .Y(n1569) );
  AND2X2 U1915 ( .A(n5140), .B(n765), .Y(n1570) );
  AND2X2 U1916 ( .A(n5121), .B(n765), .Y(n1571) );
  AND2X2 U1917 ( .A(n5753), .B(n777), .Y(n1572) );
  AND2X2 U1918 ( .A(n5751), .B(n777), .Y(n1573) );
  AND2X2 U1919 ( .A(n782), .B(n5726), .Y(n1574) );
  AND2X2 U1920 ( .A(n221), .B(n783), .Y(n1575) );
  AND2X2 U1921 ( .A(n5732), .B(n808), .Y(n1576) );
  AND2X2 U1922 ( .A(n5735), .B(n808), .Y(n1577) );
  AND2X2 U1923 ( .A(n233), .B(n809), .Y(n1578) );
  AND2X2 U1924 ( .A(n5740), .B(n809), .Y(n1579) );
  AND2X2 U1925 ( .A(n158), .B(n810), .Y(n1580) );
  AND2X2 U1926 ( .A(n128), .B(n810), .Y(n1581) );
  AND2X2 U1927 ( .A(n811), .B(n198), .Y(n1582) );
  AND2X2 U1928 ( .A(n811), .B(n177), .Y(n1583) );
  AND2X2 U1929 ( .A(n812), .B(n5120), .Y(n1584) );
  AND2X2 U1930 ( .A(n812), .B(n5119), .Y(n1585) );
  AND2X2 U1931 ( .A(n5753), .B(n824), .Y(n1586) );
  AND2X2 U1932 ( .A(n5751), .B(n824), .Y(n1587) );
  AND2X2 U1933 ( .A(n5726), .B(n5076), .Y(n1588) );
  AND2X2 U1934 ( .A(n3673), .B(n5076), .Y(n1589) );
  AND2X2 U1935 ( .A(n5729), .B(n825), .Y(n1590) );
  AND2X2 U1936 ( .A(n219), .B(n825), .Y(n1591) );
  AND2X2 U1937 ( .A(n5732), .B(n826), .Y(n1592) );
  AND2X2 U1938 ( .A(n5735), .B(n826), .Y(n1593) );
  AND2X2 U1939 ( .A(n5187), .B(n828), .Y(n1594) );
  AND2X2 U1940 ( .A(n5740), .B(n828), .Y(n1595) );
  AND2X2 U1941 ( .A(n157), .B(n829), .Y(n1596) );
  AND2X2 U1942 ( .A(n129), .B(n829), .Y(n1597) );
  AND2X2 U1943 ( .A(n200), .B(n830), .Y(n1598) );
  AND2X2 U1944 ( .A(n174), .B(n830), .Y(n1599) );
  AND2X2 U1945 ( .A(n5137), .B(n831), .Y(n1600) );
  AND2X2 U1946 ( .A(n5122), .B(n831), .Y(n1601) );
  AND2X2 U1947 ( .A(n92), .B(n832), .Y(n1602) );
  AND2X2 U1948 ( .A(n5750), .B(n832), .Y(n1603) );
  AND2X2 U1949 ( .A(n6428), .B(n19), .Y(n1604) );
  AND2X2 U1950 ( .A(n4940), .B(n833), .Y(n1605) );
  AND2X2 U1951 ( .A(n225), .B(n834), .Y(n1606) );
  AND2X2 U1952 ( .A(n217), .B(n834), .Y(n1607) );
  AND2X2 U1953 ( .A(n5732), .B(n835), .Y(n1608) );
  AND2X2 U1954 ( .A(n5735), .B(n835), .Y(n1609) );
  AND2X2 U1955 ( .A(n231), .B(n836), .Y(n1610) );
  AND2X2 U1956 ( .A(n5740), .B(n836), .Y(n1611) );
  AND2X2 U1957 ( .A(n161), .B(n837), .Y(n1612) );
  AND2X2 U1958 ( .A(n130), .B(n837), .Y(n1613) );
  AND2X2 U1959 ( .A(n199), .B(n869), .Y(n1614) );
  AND2X2 U1960 ( .A(n177), .B(n869), .Y(n1615) );
  AND2X2 U1961 ( .A(n5142), .B(n870), .Y(n1616) );
  AND2X2 U1962 ( .A(n5119), .B(n870), .Y(n1617) );
  AND2X2 U1963 ( .A(n5753), .B(n871), .Y(n1618) );
  AND2X2 U1964 ( .A(n5750), .B(n871), .Y(n1619) );
  AND2X2 U1965 ( .A(n5726), .B(n872), .Y(n1620) );
  AND2X2 U1966 ( .A(n224), .B(n873), .Y(n1621) );
  AND2X2 U1967 ( .A(n217), .B(n873), .Y(n1622) );
  AND2X2 U1968 ( .A(n5732), .B(n563), .Y(n1623) );
  AND2X2 U1969 ( .A(n5735), .B(n563), .Y(n1624) );
  AND2X2 U1970 ( .A(n233), .B(n874), .Y(n1625) );
  AND2X2 U1971 ( .A(n156), .B(n875), .Y(n1626) );
  AND2X2 U1972 ( .A(n137), .B(n875), .Y(n1627) );
  AND2X2 U1973 ( .A(n202), .B(n876), .Y(n1628) );
  AND2X2 U1974 ( .A(n176), .B(n876), .Y(n1629) );
  AND2X2 U1975 ( .A(n5143), .B(n877), .Y(n1630) );
  AND2X2 U1976 ( .A(n5121), .B(n877), .Y(n1631) );
  AND2X2 U1977 ( .A(n5753), .B(n878), .Y(n1632) );
  AND2X2 U1978 ( .A(n5751), .B(n878), .Y(n1633) );
  AND2X2 U1979 ( .A(n879), .B(n5726), .Y(n1634) );
  AND2X2 U1980 ( .A(n227), .B(n896), .Y(n1635) );
  AND2X2 U1981 ( .A(n220), .B(n896), .Y(n1636) );
  AND2X2 U1982 ( .A(n5732), .B(n897), .Y(n1637) );
  AND2X2 U1983 ( .A(n5735), .B(n897), .Y(n1638) );
  AND2X2 U1984 ( .A(n233), .B(n899), .Y(n1639) );
  AND2X2 U1985 ( .A(n5740), .B(n899), .Y(n1640) );
  AND2X2 U1986 ( .A(n160), .B(n900), .Y(n1641) );
  AND2X2 U1987 ( .A(n138), .B(n900), .Y(n1642) );
  AND2X2 U1988 ( .A(n195), .B(n901), .Y(n1643) );
  AND2X2 U1989 ( .A(n176), .B(n901), .Y(n1644) );
  AND2X2 U1990 ( .A(n5139), .B(n902), .Y(n1645) );
  AND2X2 U1991 ( .A(n5121), .B(n902), .Y(n1646) );
  AND2X2 U1992 ( .A(n3967), .B(n92), .Y(n1647) );
  AND2X2 U1993 ( .A(n3967), .B(n5750), .Y(n1648) );
  BUFX2 U1994 ( .A(n5857), .Y(n1649) );
  BUFX2 U1995 ( .A(n5935), .Y(n1650) );
  BUFX2 U1996 ( .A(n6016), .Y(n1651) );
  BUFX2 U1997 ( .A(n6087), .Y(n1652) );
  BUFX2 U1998 ( .A(n6238), .Y(n1653) );
  BUFX2 U1999 ( .A(n6318), .Y(n1654) );
  BUFX2 U2000 ( .A(n6397), .Y(n1655) );
  OR2X2 U2001 ( .A(n1139), .B(n1135), .Y(n1656) );
  INVX1 U2002 ( .A(n1656), .Y(n1657) );
  INVX1 U2003 ( .A(n5794), .Y(n1658) );
  INVX1 U2004 ( .A(n5795), .Y(n1659) );
  INVX1 U2005 ( .A(n5816), .Y(n1660) );
  INVX1 U2006 ( .A(n5817), .Y(n1661) );
  INVX1 U2007 ( .A(n5901), .Y(n1662) );
  INVX1 U2008 ( .A(n5902), .Y(n1663) );
  INVX1 U2009 ( .A(n5980), .Y(n1664) );
  INVX1 U2010 ( .A(n5981), .Y(n1665) );
  INVX1 U2011 ( .A(n6054), .Y(n1666) );
  INVX1 U2012 ( .A(n6055), .Y(n1667) );
  INVX1 U2013 ( .A(n6129), .Y(n1668) );
  INVX1 U2014 ( .A(n6204), .Y(n1669) );
  INVX1 U2015 ( .A(n6205), .Y(n1670) );
  INVX1 U2016 ( .A(n6280), .Y(n1671) );
  INVX1 U2017 ( .A(n6281), .Y(n1672) );
  INVX1 U2018 ( .A(n6360), .Y(n1673) );
  INVX1 U2019 ( .A(n6361), .Y(n1674) );
  INVX1 U2020 ( .A(n1675), .Y(n1676) );
  AND2X2 U2021 ( .A(n4108), .B(n962), .Y(n1677) );
  INVX1 U2022 ( .A(n1677), .Y(n1678) );
  AND2X2 U2023 ( .A(n925), .B(n952), .Y(n1679) );
  INVX1 U2024 ( .A(n1679), .Y(n1680) );
  AND2X2 U2025 ( .A(n929), .B(n956), .Y(n1681) );
  INVX1 U2026 ( .A(n1681), .Y(n1682) );
  AND2X2 U2027 ( .A(n3762), .B(n958), .Y(n1683) );
  INVX1 U2028 ( .A(n1683), .Y(n1684) );
  AND2X2 U2029 ( .A(n933), .B(n964), .Y(n1685) );
  INVX1 U2030 ( .A(n1685), .Y(n1686) );
  INVX1 U2031 ( .A(n1687), .Y(n1688) );
  AND2X2 U2032 ( .A(n939), .B(n968), .Y(n1689) );
  INVX1 U2033 ( .A(n1689), .Y(n1690) );
  AND2X2 U2034 ( .A(n941), .B(n970), .Y(n1691) );
  INVX1 U2035 ( .A(n1691), .Y(n1692) );
  INVX1 U2036 ( .A(n5880), .Y(n1693) );
  INVX1 U2037 ( .A(n5881), .Y(n1694) );
  INVX1 U2038 ( .A(n5960), .Y(n1695) );
  INVX1 U2039 ( .A(n5961), .Y(n1696) );
  INVX1 U2040 ( .A(n6036), .Y(n1697) );
  INVX1 U2041 ( .A(n6111), .Y(n1698) );
  INVX1 U2042 ( .A(n6112), .Y(n1699) );
  INVX1 U2043 ( .A(n6261), .Y(n1700) );
  INVX1 U2044 ( .A(n6262), .Y(n1701) );
  INVX1 U2045 ( .A(n6340), .Y(n1702) );
  INVX1 U2046 ( .A(n6341), .Y(n1703) );
  BUFX2 U2047 ( .A(n5994), .Y(n1704) );
  BUFX2 U2048 ( .A(n6294), .Y(n1705) );
  BUFX2 U2049 ( .A(n6374), .Y(n1706) );
  OR2X2 U2050 ( .A(n5812), .B(n5813), .Y(n1707) );
  OR2X2 U2051 ( .A(n5957), .B(n5956), .Y(n1708) );
  OR2X2 U2052 ( .A(n5977), .B(n5976), .Y(n1709) );
  OR2X2 U2053 ( .A(n6276), .B(n6277), .Y(n1710) );
  AND2X2 U2054 ( .A(\data_in<8> ), .B(n1530), .Y(n1711) );
  INVX1 U2055 ( .A(n1711), .Y(n1712) );
  AND2X2 U2056 ( .A(\data_in<9> ), .B(n1530), .Y(n1713) );
  INVX1 U2057 ( .A(n1713), .Y(n1714) );
  AND2X2 U2058 ( .A(\data_in<10> ), .B(n1530), .Y(n1715) );
  INVX1 U2059 ( .A(n1715), .Y(n1716) );
  AND2X2 U2060 ( .A(\data_in<11> ), .B(n1530), .Y(n1717) );
  INVX1 U2061 ( .A(n1717), .Y(n1718) );
  AND2X2 U2062 ( .A(\data_in<12> ), .B(n1530), .Y(n1719) );
  INVX1 U2063 ( .A(n1719), .Y(n1720) );
  AND2X2 U2064 ( .A(\data_in<13> ), .B(n1530), .Y(n1721) );
  INVX1 U2065 ( .A(n1721), .Y(n1722) );
  AND2X2 U2066 ( .A(\data_in<14> ), .B(n1530), .Y(n1723) );
  INVX1 U2067 ( .A(n1723), .Y(n1724) );
  AND2X2 U2068 ( .A(\data_in<15> ), .B(n1530), .Y(n1725) );
  INVX1 U2069 ( .A(n1725), .Y(n1726) );
  AND2X2 U2070 ( .A(\data_in<8> ), .B(n1532), .Y(n1727) );
  INVX1 U2071 ( .A(n1727), .Y(n1728) );
  AND2X2 U2072 ( .A(\data_in<9> ), .B(n1532), .Y(n1729) );
  INVX1 U2073 ( .A(n1729), .Y(n1730) );
  AND2X2 U2074 ( .A(\data_in<10> ), .B(n1532), .Y(n1731) );
  INVX1 U2075 ( .A(n1731), .Y(n1732) );
  AND2X2 U2076 ( .A(\data_in<11> ), .B(n1532), .Y(n1733) );
  INVX1 U2077 ( .A(n1733), .Y(n1734) );
  AND2X2 U2078 ( .A(\data_in<12> ), .B(n1532), .Y(n1735) );
  INVX1 U2079 ( .A(n1735), .Y(n1736) );
  AND2X2 U2080 ( .A(\data_in<13> ), .B(n1532), .Y(n1737) );
  INVX1 U2081 ( .A(n1737), .Y(n1738) );
  AND2X2 U2082 ( .A(\data_in<14> ), .B(n1532), .Y(n1739) );
  INVX1 U2083 ( .A(n1739), .Y(n1740) );
  AND2X2 U2084 ( .A(\data_in<15> ), .B(n1532), .Y(n1741) );
  INVX1 U2085 ( .A(n1741), .Y(n1742) );
  AND2X2 U2086 ( .A(\data_in<8> ), .B(n1534), .Y(n1743) );
  INVX1 U2087 ( .A(n1743), .Y(n1744) );
  AND2X2 U2088 ( .A(\data_in<9> ), .B(n1534), .Y(n1745) );
  INVX1 U2089 ( .A(n1745), .Y(n1746) );
  AND2X2 U2090 ( .A(\data_in<10> ), .B(n1534), .Y(n1747) );
  INVX1 U2091 ( .A(n1747), .Y(n1748) );
  AND2X2 U2092 ( .A(\data_in<11> ), .B(n1534), .Y(n1749) );
  INVX1 U2093 ( .A(n1749), .Y(n1750) );
  AND2X2 U2094 ( .A(\data_in<12> ), .B(n1534), .Y(n1751) );
  INVX1 U2095 ( .A(n1751), .Y(n1752) );
  AND2X2 U2096 ( .A(\data_in<13> ), .B(n1534), .Y(n1753) );
  INVX1 U2097 ( .A(n1753), .Y(n1754) );
  AND2X2 U2098 ( .A(\data_in<14> ), .B(n1534), .Y(n1755) );
  INVX1 U2099 ( .A(n1755), .Y(n1756) );
  AND2X2 U2100 ( .A(\data_in<15> ), .B(n1534), .Y(n1757) );
  INVX1 U2101 ( .A(n1757), .Y(n1758) );
  AND2X2 U2102 ( .A(\data_in<8> ), .B(n1536), .Y(n1759) );
  INVX1 U2103 ( .A(n1759), .Y(n1760) );
  AND2X2 U2104 ( .A(\data_in<9> ), .B(n1536), .Y(n1761) );
  INVX1 U2105 ( .A(n1761), .Y(n1762) );
  AND2X2 U2106 ( .A(\data_in<10> ), .B(n1536), .Y(n1763) );
  INVX1 U2107 ( .A(n1763), .Y(n1764) );
  AND2X2 U2108 ( .A(\data_in<11> ), .B(n1536), .Y(n1765) );
  INVX1 U2109 ( .A(n1765), .Y(n1766) );
  AND2X2 U2110 ( .A(\data_in<12> ), .B(n1536), .Y(n1767) );
  INVX1 U2111 ( .A(n1767), .Y(n1768) );
  AND2X2 U2112 ( .A(\data_in<13> ), .B(n1536), .Y(n1769) );
  INVX1 U2113 ( .A(n1769), .Y(n1770) );
  AND2X2 U2114 ( .A(\data_in<14> ), .B(n1536), .Y(n1771) );
  INVX1 U2115 ( .A(n1771), .Y(n1772) );
  AND2X2 U2116 ( .A(\data_in<15> ), .B(n1536), .Y(n1773) );
  INVX1 U2117 ( .A(n1773), .Y(n1774) );
  AND2X2 U2118 ( .A(\data_in<8> ), .B(n1538), .Y(n1775) );
  INVX1 U2119 ( .A(n1775), .Y(n1776) );
  AND2X2 U2120 ( .A(\data_in<9> ), .B(n1538), .Y(n1777) );
  INVX1 U2121 ( .A(n1777), .Y(n1778) );
  AND2X2 U2122 ( .A(\data_in<10> ), .B(n1538), .Y(n1779) );
  INVX1 U2123 ( .A(n1779), .Y(n1780) );
  AND2X2 U2124 ( .A(\data_in<11> ), .B(n1538), .Y(n1781) );
  INVX1 U2125 ( .A(n1781), .Y(n1782) );
  AND2X2 U2126 ( .A(\data_in<12> ), .B(n1538), .Y(n1783) );
  INVX1 U2127 ( .A(n1783), .Y(n1784) );
  AND2X2 U2128 ( .A(\data_in<13> ), .B(n1538), .Y(n1785) );
  INVX1 U2129 ( .A(n1785), .Y(n1786) );
  AND2X2 U2130 ( .A(\data_in<14> ), .B(n1538), .Y(n1787) );
  INVX1 U2131 ( .A(n1787), .Y(n1788) );
  AND2X2 U2132 ( .A(\data_in<15> ), .B(n1538), .Y(n1789) );
  INVX1 U2133 ( .A(n1789), .Y(n1790) );
  AND2X2 U2134 ( .A(\data_in<8> ), .B(n1540), .Y(n1791) );
  INVX1 U2135 ( .A(n1791), .Y(n1792) );
  AND2X2 U2136 ( .A(\data_in<9> ), .B(n1540), .Y(n1793) );
  INVX1 U2137 ( .A(n1793), .Y(n1794) );
  AND2X2 U2138 ( .A(\data_in<10> ), .B(n1540), .Y(n1795) );
  INVX1 U2139 ( .A(n1795), .Y(n1796) );
  AND2X2 U2140 ( .A(\data_in<11> ), .B(n1540), .Y(n1797) );
  INVX1 U2141 ( .A(n1797), .Y(n1798) );
  AND2X2 U2142 ( .A(\data_in<12> ), .B(n1540), .Y(n1799) );
  INVX1 U2143 ( .A(n1799), .Y(n1800) );
  AND2X2 U2144 ( .A(\data_in<13> ), .B(n1540), .Y(n1801) );
  INVX1 U2145 ( .A(n1801), .Y(n1802) );
  AND2X2 U2146 ( .A(\data_in<14> ), .B(n1540), .Y(n1803) );
  INVX1 U2147 ( .A(n1803), .Y(n1804) );
  AND2X2 U2148 ( .A(\data_in<15> ), .B(n1540), .Y(n1805) );
  INVX1 U2149 ( .A(n1805), .Y(n1806) );
  AND2X2 U2150 ( .A(\data_in<8> ), .B(n1542), .Y(n1807) );
  INVX1 U2151 ( .A(n1807), .Y(n1808) );
  AND2X2 U2152 ( .A(\data_in<9> ), .B(n1542), .Y(n1809) );
  INVX1 U2153 ( .A(n1809), .Y(n1810) );
  AND2X2 U2154 ( .A(\data_in<10> ), .B(n1542), .Y(n1811) );
  INVX1 U2155 ( .A(n1811), .Y(n1812) );
  AND2X2 U2156 ( .A(\data_in<11> ), .B(n1542), .Y(n1813) );
  INVX1 U2157 ( .A(n1813), .Y(n1814) );
  AND2X2 U2158 ( .A(\data_in<12> ), .B(n1542), .Y(n1815) );
  INVX1 U2159 ( .A(n1815), .Y(n2328) );
  AND2X2 U2160 ( .A(\data_in<13> ), .B(n1542), .Y(n2329) );
  INVX1 U2161 ( .A(n2329), .Y(n2330) );
  AND2X2 U2162 ( .A(\data_in<14> ), .B(n1542), .Y(n2331) );
  INVX1 U2163 ( .A(n2331), .Y(n2332) );
  AND2X2 U2164 ( .A(\data_in<15> ), .B(n1542), .Y(n2333) );
  INVX1 U2165 ( .A(n2333), .Y(n2334) );
  AND2X2 U2166 ( .A(\data_in<8> ), .B(n1544), .Y(n2335) );
  INVX1 U2167 ( .A(n2335), .Y(n2336) );
  AND2X2 U2168 ( .A(\data_in<9> ), .B(n1544), .Y(n2337) );
  INVX1 U2169 ( .A(n2337), .Y(n2338) );
  AND2X2 U2170 ( .A(\data_in<10> ), .B(n1544), .Y(n2339) );
  INVX1 U2171 ( .A(n2339), .Y(n2340) );
  AND2X2 U2172 ( .A(\data_in<11> ), .B(n1544), .Y(n2341) );
  INVX1 U2173 ( .A(n2341), .Y(n2342) );
  AND2X2 U2174 ( .A(\data_in<12> ), .B(n1544), .Y(n2343) );
  INVX1 U2175 ( .A(n2343), .Y(n2344) );
  AND2X2 U2176 ( .A(\data_in<13> ), .B(n1544), .Y(n2345) );
  INVX1 U2177 ( .A(n2345), .Y(n2346) );
  AND2X2 U2178 ( .A(\data_in<14> ), .B(n1544), .Y(n2347) );
  INVX1 U2179 ( .A(n2347), .Y(n2348) );
  AND2X2 U2180 ( .A(\data_in<15> ), .B(n1544), .Y(n2349) );
  INVX1 U2181 ( .A(n2349), .Y(n2350) );
  AND2X2 U2182 ( .A(\data_in<8> ), .B(n1546), .Y(n2351) );
  INVX1 U2183 ( .A(n2351), .Y(n2352) );
  AND2X2 U2184 ( .A(\data_in<9> ), .B(n1546), .Y(n2353) );
  INVX1 U2185 ( .A(n2353), .Y(n2354) );
  AND2X2 U2186 ( .A(\data_in<10> ), .B(n1546), .Y(n2355) );
  INVX1 U2187 ( .A(n2355), .Y(n2356) );
  AND2X2 U2188 ( .A(\data_in<11> ), .B(n1546), .Y(n2357) );
  INVX1 U2189 ( .A(n2357), .Y(n2358) );
  AND2X2 U2190 ( .A(\data_in<12> ), .B(n1546), .Y(n2359) );
  INVX1 U2191 ( .A(n2359), .Y(n2360) );
  AND2X2 U2192 ( .A(\data_in<13> ), .B(n1546), .Y(n2361) );
  INVX1 U2193 ( .A(n2361), .Y(n2362) );
  AND2X2 U2194 ( .A(\data_in<14> ), .B(n1546), .Y(n2363) );
  INVX1 U2195 ( .A(n2363), .Y(n2364) );
  AND2X2 U2196 ( .A(\data_in<15> ), .B(n1546), .Y(n2365) );
  INVX1 U2197 ( .A(n2365), .Y(n2366) );
  AND2X2 U2198 ( .A(\data_in<8> ), .B(n1548), .Y(n2367) );
  INVX1 U2199 ( .A(n2367), .Y(n2368) );
  AND2X2 U2200 ( .A(\data_in<9> ), .B(n1548), .Y(n2369) );
  INVX1 U2201 ( .A(n2369), .Y(n2370) );
  AND2X2 U2202 ( .A(\data_in<10> ), .B(n1548), .Y(n2371) );
  INVX1 U2203 ( .A(n2371), .Y(n2372) );
  AND2X2 U2204 ( .A(\data_in<11> ), .B(n1548), .Y(n2373) );
  INVX1 U2205 ( .A(n2373), .Y(n2374) );
  AND2X2 U2206 ( .A(\data_in<12> ), .B(n1548), .Y(n2375) );
  INVX1 U2207 ( .A(n2375), .Y(n2376) );
  AND2X2 U2208 ( .A(\data_in<13> ), .B(n1548), .Y(n2377) );
  INVX1 U2209 ( .A(n2377), .Y(n2378) );
  AND2X2 U2210 ( .A(\data_in<14> ), .B(n1548), .Y(n2379) );
  INVX1 U2211 ( .A(n2379), .Y(n2380) );
  AND2X2 U2212 ( .A(\data_in<15> ), .B(n1548), .Y(n2381) );
  INVX1 U2213 ( .A(n2381), .Y(n2382) );
  AND2X2 U2214 ( .A(\data_in<8> ), .B(n1550), .Y(n2383) );
  INVX1 U2215 ( .A(n2383), .Y(n2384) );
  AND2X2 U2216 ( .A(\data_in<9> ), .B(n1550), .Y(n2385) );
  INVX1 U2217 ( .A(n2385), .Y(n2386) );
  AND2X2 U2218 ( .A(\data_in<10> ), .B(n1550), .Y(n2387) );
  INVX1 U2219 ( .A(n2387), .Y(n2388) );
  AND2X2 U2220 ( .A(\data_in<11> ), .B(n1550), .Y(n2389) );
  INVX1 U2221 ( .A(n2389), .Y(n2390) );
  AND2X2 U2222 ( .A(\data_in<12> ), .B(n1550), .Y(n2391) );
  INVX1 U2223 ( .A(n2391), .Y(n2392) );
  AND2X2 U2224 ( .A(\data_in<13> ), .B(n1550), .Y(n2393) );
  INVX1 U2225 ( .A(n2393), .Y(n2394) );
  AND2X2 U2226 ( .A(\data_in<14> ), .B(n1550), .Y(n2395) );
  INVX1 U2227 ( .A(n2395), .Y(n2396) );
  AND2X2 U2228 ( .A(\data_in<15> ), .B(n1550), .Y(n2397) );
  INVX1 U2229 ( .A(n2397), .Y(n2398) );
  AND2X2 U2230 ( .A(\data_in<10> ), .B(n1552), .Y(n2399) );
  INVX1 U2231 ( .A(n2399), .Y(n2400) );
  AND2X2 U2232 ( .A(\data_in<13> ), .B(n43), .Y(n2401) );
  INVX1 U2233 ( .A(n2401), .Y(n2402) );
  AND2X2 U2234 ( .A(\data_in<8> ), .B(n1554), .Y(n2403) );
  INVX1 U2235 ( .A(n2403), .Y(n2404) );
  AND2X2 U2236 ( .A(\data_in<9> ), .B(n1554), .Y(n2405) );
  INVX1 U2237 ( .A(n2405), .Y(n2406) );
  AND2X2 U2238 ( .A(\data_in<10> ), .B(n1554), .Y(n2407) );
  INVX1 U2239 ( .A(n2407), .Y(n2408) );
  AND2X2 U2240 ( .A(\data_in<11> ), .B(n1554), .Y(n2409) );
  INVX1 U2241 ( .A(n2409), .Y(n2410) );
  AND2X2 U2242 ( .A(\data_in<12> ), .B(n1554), .Y(n2411) );
  INVX1 U2243 ( .A(n2411), .Y(n2412) );
  AND2X2 U2244 ( .A(\data_in<13> ), .B(n1554), .Y(n2413) );
  INVX1 U2245 ( .A(n2413), .Y(n2414) );
  AND2X2 U2246 ( .A(\data_in<14> ), .B(n1554), .Y(n2415) );
  INVX1 U2247 ( .A(n2415), .Y(n2416) );
  AND2X2 U2248 ( .A(\data_in<15> ), .B(n1554), .Y(n2417) );
  INVX1 U2249 ( .A(n2417), .Y(n2418) );
  AND2X2 U2250 ( .A(\data_in<8> ), .B(n1556), .Y(n2419) );
  INVX1 U2251 ( .A(n2419), .Y(n2420) );
  AND2X2 U2252 ( .A(\data_in<9> ), .B(n1556), .Y(n2421) );
  INVX1 U2253 ( .A(n2421), .Y(n2422) );
  AND2X2 U2254 ( .A(\data_in<10> ), .B(n1556), .Y(n2423) );
  INVX1 U2255 ( .A(n2423), .Y(n2424) );
  AND2X2 U2256 ( .A(\data_in<11> ), .B(n1556), .Y(n2425) );
  INVX1 U2257 ( .A(n2425), .Y(n2426) );
  AND2X2 U2258 ( .A(\data_in<12> ), .B(n1556), .Y(n2427) );
  INVX1 U2259 ( .A(n2427), .Y(n2428) );
  AND2X2 U2260 ( .A(\data_in<13> ), .B(n1556), .Y(n2429) );
  INVX1 U2261 ( .A(n2429), .Y(n2430) );
  AND2X2 U2262 ( .A(\data_in<14> ), .B(n1556), .Y(n2431) );
  INVX1 U2263 ( .A(n2431), .Y(n2432) );
  AND2X2 U2264 ( .A(\data_in<15> ), .B(n1556), .Y(n2433) );
  INVX1 U2265 ( .A(n2433), .Y(n2434) );
  AND2X2 U2266 ( .A(\data_in<8> ), .B(n1558), .Y(n2435) );
  INVX1 U2267 ( .A(n2435), .Y(n2436) );
  AND2X2 U2268 ( .A(\data_in<9> ), .B(n1558), .Y(n2437) );
  INVX1 U2269 ( .A(n2437), .Y(n2438) );
  AND2X2 U2270 ( .A(\data_in<10> ), .B(n1558), .Y(n2439) );
  INVX1 U2271 ( .A(n2439), .Y(n2440) );
  AND2X2 U2272 ( .A(\data_in<11> ), .B(n1558), .Y(n2441) );
  INVX1 U2273 ( .A(n2441), .Y(n2442) );
  AND2X2 U2274 ( .A(\data_in<12> ), .B(n1558), .Y(n2443) );
  INVX1 U2275 ( .A(n2443), .Y(n2444) );
  AND2X2 U2276 ( .A(\data_in<13> ), .B(n1558), .Y(n2445) );
  INVX1 U2277 ( .A(n2445), .Y(n2446) );
  AND2X2 U2278 ( .A(\data_in<14> ), .B(n1558), .Y(n2447) );
  INVX1 U2279 ( .A(n2447), .Y(n2448) );
  AND2X2 U2280 ( .A(\data_in<15> ), .B(n1558), .Y(n2449) );
  INVX1 U2281 ( .A(n2449), .Y(n2450) );
  AND2X2 U2282 ( .A(\data_in<8> ), .B(n1559), .Y(n2451) );
  INVX1 U2283 ( .A(n2451), .Y(n2452) );
  AND2X2 U2284 ( .A(\data_in<9> ), .B(n1559), .Y(n2453) );
  INVX1 U2285 ( .A(n2453), .Y(n2454) );
  AND2X2 U2286 ( .A(\data_in<10> ), .B(n1559), .Y(n2455) );
  INVX1 U2287 ( .A(n2455), .Y(n2456) );
  AND2X2 U2288 ( .A(\data_in<11> ), .B(n1559), .Y(n2457) );
  INVX1 U2289 ( .A(n2457), .Y(n2458) );
  AND2X2 U2290 ( .A(\data_in<12> ), .B(n1559), .Y(n2459) );
  INVX1 U2291 ( .A(n2459), .Y(n2460) );
  AND2X2 U2292 ( .A(\data_in<13> ), .B(n1559), .Y(n2461) );
  INVX1 U2293 ( .A(n2461), .Y(n2462) );
  AND2X2 U2294 ( .A(\data_in<14> ), .B(n1559), .Y(n2463) );
  INVX1 U2295 ( .A(n2463), .Y(n2464) );
  AND2X2 U2296 ( .A(\data_in<15> ), .B(n1559), .Y(n2465) );
  INVX1 U2297 ( .A(n2465), .Y(n2466) );
  AND2X2 U2298 ( .A(\data_in<10> ), .B(n1565), .Y(n2467) );
  INVX1 U2299 ( .A(n2467), .Y(n2468) );
  AND2X2 U2300 ( .A(\data_in<13> ), .B(n1565), .Y(n2469) );
  INVX1 U2301 ( .A(n2469), .Y(n2470) );
  AND2X2 U2302 ( .A(\data_in<10> ), .B(n13), .Y(n2471) );
  INVX1 U2303 ( .A(n2471), .Y(n2472) );
  AND2X2 U2304 ( .A(n1567), .B(\data_in<13> ), .Y(n2473) );
  INVX1 U2305 ( .A(n2473), .Y(n2474) );
  AND2X2 U2306 ( .A(\data_in<10> ), .B(n1569), .Y(n2475) );
  INVX1 U2307 ( .A(n2475), .Y(n2476) );
  AND2X2 U2308 ( .A(\data_in<13> ), .B(n1569), .Y(n2477) );
  INVX1 U2309 ( .A(n2477), .Y(n2478) );
  AND2X2 U2310 ( .A(\data_in<10> ), .B(n64), .Y(n2479) );
  INVX1 U2311 ( .A(n2479), .Y(n2480) );
  AND2X2 U2312 ( .A(\data_in<13> ), .B(n64), .Y(n2481) );
  INVX1 U2313 ( .A(n2481), .Y(n2482) );
  AND2X2 U2314 ( .A(\data_in<8> ), .B(n3843), .Y(n2483) );
  INVX1 U2315 ( .A(n2483), .Y(n2484) );
  AND2X2 U2316 ( .A(\data_in<9> ), .B(n3843), .Y(n2485) );
  INVX1 U2317 ( .A(n2485), .Y(n2486) );
  AND2X2 U2318 ( .A(\data_in<10> ), .B(n3843), .Y(n2487) );
  INVX1 U2319 ( .A(n2487), .Y(n2488) );
  AND2X2 U2320 ( .A(\data_in<11> ), .B(n3843), .Y(n2489) );
  INVX1 U2321 ( .A(n2489), .Y(n2490) );
  AND2X2 U2322 ( .A(\data_in<12> ), .B(n3843), .Y(n2491) );
  INVX1 U2323 ( .A(n2491), .Y(n2492) );
  AND2X2 U2324 ( .A(\data_in<13> ), .B(n3843), .Y(n2493) );
  INVX1 U2325 ( .A(n2493), .Y(n2494) );
  AND2X2 U2326 ( .A(\data_in<14> ), .B(n3843), .Y(n2495) );
  INVX1 U2327 ( .A(n2495), .Y(n2496) );
  AND2X2 U2328 ( .A(\data_in<15> ), .B(n3843), .Y(n2497) );
  INVX1 U2329 ( .A(n2497), .Y(n2498) );
  AND2X2 U2330 ( .A(\data_in<10> ), .B(n1575), .Y(n2499) );
  INVX1 U2331 ( .A(n2499), .Y(n2500) );
  AND2X2 U2332 ( .A(\data_in<13> ), .B(n1575), .Y(n2501) );
  INVX1 U2333 ( .A(n2501), .Y(n2502) );
  AND2X2 U2334 ( .A(\data_in<8> ), .B(n1577), .Y(n2503) );
  INVX1 U2335 ( .A(n2503), .Y(n2504) );
  AND2X2 U2336 ( .A(\data_in<9> ), .B(n1577), .Y(n2505) );
  INVX1 U2337 ( .A(n2505), .Y(n2506) );
  AND2X2 U2338 ( .A(\data_in<10> ), .B(n1577), .Y(n2507) );
  INVX1 U2339 ( .A(n2507), .Y(n2508) );
  AND2X2 U2340 ( .A(\data_in<11> ), .B(n1577), .Y(n2509) );
  INVX1 U2341 ( .A(n2509), .Y(n2510) );
  AND2X2 U2342 ( .A(\data_in<12> ), .B(n1577), .Y(n2511) );
  INVX1 U2343 ( .A(n2511), .Y(n2512) );
  AND2X2 U2344 ( .A(\data_in<13> ), .B(n1577), .Y(n2513) );
  INVX1 U2345 ( .A(n2513), .Y(n2514) );
  AND2X2 U2346 ( .A(\data_in<14> ), .B(n1577), .Y(n2515) );
  INVX1 U2347 ( .A(n2515), .Y(n2516) );
  AND2X2 U2348 ( .A(\data_in<15> ), .B(n1577), .Y(n2517) );
  INVX1 U2349 ( .A(n2517), .Y(n2518) );
  AND2X2 U2350 ( .A(\data_in<8> ), .B(n1579), .Y(n2519) );
  INVX1 U2351 ( .A(n2519), .Y(n2520) );
  AND2X2 U2352 ( .A(\data_in<9> ), .B(n1579), .Y(n2521) );
  INVX1 U2353 ( .A(n2521), .Y(n2522) );
  AND2X2 U2354 ( .A(\data_in<10> ), .B(n1579), .Y(n2523) );
  INVX1 U2355 ( .A(n2523), .Y(n2524) );
  AND2X2 U2356 ( .A(\data_in<11> ), .B(n1579), .Y(n2525) );
  INVX1 U2357 ( .A(n2525), .Y(n2526) );
  AND2X2 U2358 ( .A(\data_in<12> ), .B(n1579), .Y(n2527) );
  INVX1 U2359 ( .A(n2527), .Y(n2528) );
  AND2X2 U2360 ( .A(\data_in<13> ), .B(n1579), .Y(n2529) );
  INVX1 U2361 ( .A(n2529), .Y(n2530) );
  AND2X2 U2362 ( .A(\data_in<14> ), .B(n1579), .Y(n2531) );
  INVX1 U2363 ( .A(n2531), .Y(n2532) );
  AND2X2 U2364 ( .A(\data_in<15> ), .B(n1579), .Y(n2533) );
  INVX1 U2365 ( .A(n2533), .Y(n2534) );
  AND2X2 U2366 ( .A(\data_in<8> ), .B(n1581), .Y(n2535) );
  INVX1 U2367 ( .A(n2535), .Y(n2536) );
  AND2X2 U2368 ( .A(\data_in<9> ), .B(n1581), .Y(n2537) );
  INVX1 U2369 ( .A(n2537), .Y(n2538) );
  AND2X2 U2370 ( .A(\data_in<10> ), .B(n1581), .Y(n2539) );
  INVX1 U2371 ( .A(n2539), .Y(n2540) );
  AND2X2 U2372 ( .A(\data_in<11> ), .B(n1581), .Y(n2541) );
  INVX1 U2373 ( .A(n2541), .Y(n2542) );
  AND2X2 U2374 ( .A(\data_in<12> ), .B(n1581), .Y(n2543) );
  INVX1 U2375 ( .A(n2543), .Y(n2544) );
  AND2X2 U2376 ( .A(\data_in<13> ), .B(n1581), .Y(n2545) );
  INVX1 U2377 ( .A(n2545), .Y(n2546) );
  AND2X2 U2378 ( .A(\data_in<14> ), .B(n1581), .Y(n2547) );
  INVX1 U2379 ( .A(n2547), .Y(n2548) );
  AND2X2 U2380 ( .A(\data_in<15> ), .B(n1581), .Y(n2549) );
  INVX1 U2381 ( .A(n2549), .Y(n2550) );
  AND2X2 U2382 ( .A(\data_in<8> ), .B(n1583), .Y(n2551) );
  INVX1 U2383 ( .A(n2551), .Y(n2552) );
  AND2X2 U2384 ( .A(\data_in<9> ), .B(n1583), .Y(n2553) );
  INVX1 U2385 ( .A(n2553), .Y(n2554) );
  AND2X2 U2386 ( .A(\data_in<10> ), .B(n1583), .Y(n2555) );
  INVX1 U2387 ( .A(n2555), .Y(n2556) );
  AND2X2 U2388 ( .A(\data_in<11> ), .B(n1583), .Y(n2557) );
  INVX1 U2389 ( .A(n2557), .Y(n2558) );
  AND2X2 U2390 ( .A(\data_in<12> ), .B(n1583), .Y(n2559) );
  INVX1 U2391 ( .A(n2559), .Y(n2560) );
  AND2X2 U2392 ( .A(\data_in<13> ), .B(n1583), .Y(n2561) );
  INVX1 U2393 ( .A(n2561), .Y(n2562) );
  AND2X2 U2394 ( .A(\data_in<14> ), .B(n1583), .Y(n2563) );
  INVX1 U2395 ( .A(n2563), .Y(n2564) );
  AND2X2 U2396 ( .A(\data_in<15> ), .B(n1583), .Y(n2565) );
  INVX1 U2397 ( .A(n2565), .Y(n2566) );
  AND2X2 U2398 ( .A(\data_in<10> ), .B(n1585), .Y(n2567) );
  INVX1 U2399 ( .A(n2567), .Y(n2568) );
  AND2X2 U2400 ( .A(\data_in<13> ), .B(n9), .Y(n2569) );
  INVX1 U2401 ( .A(n2569), .Y(n2570) );
  AND2X2 U2402 ( .A(\data_in<8> ), .B(n1587), .Y(n2571) );
  INVX1 U2403 ( .A(n2571), .Y(n2572) );
  AND2X2 U2404 ( .A(\data_in<9> ), .B(n1587), .Y(n2573) );
  INVX1 U2405 ( .A(n2573), .Y(n2574) );
  AND2X2 U2406 ( .A(\data_in<10> ), .B(n1587), .Y(n2575) );
  INVX1 U2407 ( .A(n2575), .Y(n2576) );
  AND2X2 U2408 ( .A(\data_in<11> ), .B(n1587), .Y(n2577) );
  INVX1 U2409 ( .A(n2577), .Y(n2578) );
  AND2X2 U2410 ( .A(\data_in<12> ), .B(n1587), .Y(n2579) );
  INVX1 U2411 ( .A(n2579), .Y(n2580) );
  AND2X2 U2412 ( .A(\data_in<13> ), .B(n1587), .Y(n2581) );
  INVX1 U2413 ( .A(n2581), .Y(n2582) );
  AND2X2 U2414 ( .A(\data_in<14> ), .B(n1587), .Y(n2583) );
  INVX1 U2415 ( .A(n2583), .Y(n2584) );
  AND2X2 U2416 ( .A(\data_in<15> ), .B(n1587), .Y(n2585) );
  INVX1 U2417 ( .A(n2585), .Y(n2586) );
  AND2X2 U2418 ( .A(\data_in<8> ), .B(n1589), .Y(n2587) );
  INVX1 U2419 ( .A(n2587), .Y(n2588) );
  AND2X2 U2420 ( .A(\data_in<9> ), .B(n1589), .Y(n2589) );
  INVX1 U2421 ( .A(n2589), .Y(n2590) );
  AND2X2 U2422 ( .A(\data_in<10> ), .B(n1589), .Y(n2591) );
  INVX1 U2423 ( .A(n2591), .Y(n2592) );
  AND2X2 U2424 ( .A(\data_in<11> ), .B(n1589), .Y(n2593) );
  INVX1 U2425 ( .A(n2593), .Y(n2594) );
  AND2X2 U2426 ( .A(\data_in<12> ), .B(n1589), .Y(n2595) );
  INVX1 U2427 ( .A(n2595), .Y(n2596) );
  AND2X2 U2428 ( .A(\data_in<13> ), .B(n1589), .Y(n2597) );
  INVX1 U2429 ( .A(n2597), .Y(n2598) );
  AND2X2 U2430 ( .A(\data_in<14> ), .B(n1589), .Y(n2599) );
  INVX1 U2431 ( .A(n2599), .Y(n2600) );
  AND2X2 U2432 ( .A(\data_in<15> ), .B(n1589), .Y(n2601) );
  INVX1 U2433 ( .A(n2601), .Y(n2602) );
  AND2X2 U2434 ( .A(\data_in<8> ), .B(n1591), .Y(n2603) );
  INVX1 U2435 ( .A(n2603), .Y(n2604) );
  AND2X2 U2436 ( .A(\data_in<9> ), .B(n1591), .Y(n2605) );
  INVX1 U2437 ( .A(n2605), .Y(n2606) );
  AND2X2 U2438 ( .A(\data_in<10> ), .B(n1591), .Y(n2607) );
  INVX1 U2439 ( .A(n2607), .Y(n2608) );
  AND2X2 U2440 ( .A(\data_in<11> ), .B(n1591), .Y(n2609) );
  INVX1 U2441 ( .A(n2609), .Y(n2610) );
  AND2X2 U2442 ( .A(\data_in<12> ), .B(n1591), .Y(n2611) );
  INVX1 U2443 ( .A(n2611), .Y(n2612) );
  AND2X2 U2444 ( .A(\data_in<13> ), .B(n1591), .Y(n2613) );
  INVX1 U2445 ( .A(n2613), .Y(n2614) );
  AND2X2 U2446 ( .A(\data_in<14> ), .B(n1591), .Y(n2615) );
  INVX1 U2447 ( .A(n2615), .Y(n2616) );
  AND2X2 U2448 ( .A(\data_in<15> ), .B(n1591), .Y(n2617) );
  INVX1 U2449 ( .A(n2617), .Y(n2618) );
  AND2X2 U2450 ( .A(\data_in<8> ), .B(n1593), .Y(n2619) );
  INVX1 U2451 ( .A(n2619), .Y(n2620) );
  AND2X2 U2452 ( .A(\data_in<9> ), .B(n1593), .Y(n2621) );
  INVX1 U2453 ( .A(n2621), .Y(n2622) );
  AND2X2 U2454 ( .A(\data_in<10> ), .B(n1593), .Y(n2623) );
  INVX1 U2455 ( .A(n2623), .Y(n2624) );
  AND2X2 U2456 ( .A(\data_in<11> ), .B(n1593), .Y(n2625) );
  INVX1 U2457 ( .A(n2625), .Y(n2626) );
  AND2X2 U2458 ( .A(\data_in<12> ), .B(n1593), .Y(n2627) );
  INVX1 U2459 ( .A(n2627), .Y(n2628) );
  AND2X2 U2460 ( .A(\data_in<13> ), .B(n1593), .Y(n2629) );
  INVX1 U2461 ( .A(n2629), .Y(n2630) );
  AND2X2 U2462 ( .A(\data_in<14> ), .B(n1593), .Y(n2631) );
  INVX1 U2463 ( .A(n2631), .Y(n2632) );
  AND2X2 U2464 ( .A(\data_in<15> ), .B(n1593), .Y(n2633) );
  INVX1 U2465 ( .A(n2633), .Y(n2634) );
  AND2X2 U2466 ( .A(\data_in<8> ), .B(n1595), .Y(n2635) );
  INVX1 U2467 ( .A(n2635), .Y(n2636) );
  AND2X2 U2468 ( .A(\data_in<9> ), .B(n1595), .Y(n2637) );
  INVX1 U2469 ( .A(n2637), .Y(n2638) );
  AND2X2 U2470 ( .A(\data_in<10> ), .B(n1595), .Y(n2639) );
  INVX1 U2471 ( .A(n2639), .Y(n2640) );
  AND2X2 U2472 ( .A(\data_in<11> ), .B(n1595), .Y(n2641) );
  INVX1 U2473 ( .A(n2641), .Y(n2642) );
  AND2X2 U2474 ( .A(\data_in<12> ), .B(n1595), .Y(n2643) );
  INVX1 U2475 ( .A(n2643), .Y(n2644) );
  AND2X2 U2476 ( .A(\data_in<13> ), .B(n1595), .Y(n2645) );
  INVX1 U2477 ( .A(n2645), .Y(n2646) );
  AND2X2 U2478 ( .A(\data_in<14> ), .B(n1595), .Y(n2647) );
  INVX1 U2479 ( .A(n2647), .Y(n2648) );
  AND2X2 U2480 ( .A(\data_in<15> ), .B(n1595), .Y(n2649) );
  INVX1 U2481 ( .A(n2649), .Y(n2650) );
  AND2X2 U2482 ( .A(\data_in<8> ), .B(n1597), .Y(n2651) );
  INVX1 U2483 ( .A(n2651), .Y(n2652) );
  AND2X2 U2484 ( .A(\data_in<9> ), .B(n1597), .Y(n2653) );
  INVX1 U2485 ( .A(n2653), .Y(n2654) );
  AND2X2 U2486 ( .A(\data_in<10> ), .B(n1597), .Y(n2655) );
  INVX1 U2487 ( .A(n2655), .Y(n2656) );
  AND2X2 U2488 ( .A(\data_in<11> ), .B(n1597), .Y(n2657) );
  INVX1 U2489 ( .A(n2657), .Y(n2658) );
  AND2X2 U2490 ( .A(\data_in<12> ), .B(n1597), .Y(n2659) );
  INVX1 U2491 ( .A(n2659), .Y(n2660) );
  AND2X2 U2492 ( .A(\data_in<13> ), .B(n1597), .Y(n2661) );
  INVX1 U2493 ( .A(n2661), .Y(n2662) );
  AND2X2 U2494 ( .A(\data_in<14> ), .B(n1597), .Y(n2663) );
  INVX1 U2495 ( .A(n2663), .Y(n2664) );
  AND2X2 U2496 ( .A(\data_in<15> ), .B(n1597), .Y(n2665) );
  INVX1 U2497 ( .A(n2665), .Y(n2666) );
  AND2X2 U2498 ( .A(\data_in<8> ), .B(n1599), .Y(n2667) );
  INVX1 U2499 ( .A(n2667), .Y(n2668) );
  AND2X2 U2500 ( .A(\data_in<9> ), .B(n1599), .Y(n2669) );
  INVX1 U2501 ( .A(n2669), .Y(n2670) );
  AND2X2 U2502 ( .A(\data_in<10> ), .B(n1599), .Y(n2671) );
  INVX1 U2503 ( .A(n2671), .Y(n2672) );
  AND2X2 U2504 ( .A(\data_in<11> ), .B(n1599), .Y(n2673) );
  INVX1 U2505 ( .A(n2673), .Y(n2674) );
  AND2X2 U2506 ( .A(\data_in<12> ), .B(n1599), .Y(n2675) );
  INVX1 U2507 ( .A(n2675), .Y(n2676) );
  AND2X2 U2508 ( .A(\data_in<13> ), .B(n1599), .Y(n2677) );
  INVX1 U2509 ( .A(n2677), .Y(n2678) );
  AND2X2 U2510 ( .A(\data_in<14> ), .B(n1599), .Y(n2679) );
  INVX1 U2511 ( .A(n2679), .Y(n2680) );
  AND2X2 U2512 ( .A(\data_in<15> ), .B(n1599), .Y(n2681) );
  INVX1 U2513 ( .A(n2681), .Y(n2682) );
  AND2X2 U2514 ( .A(\data_in<8> ), .B(n1601), .Y(n2683) );
  INVX1 U2515 ( .A(n2683), .Y(n2684) );
  AND2X2 U2516 ( .A(\data_in<9> ), .B(n1601), .Y(n2685) );
  INVX1 U2517 ( .A(n2685), .Y(n2686) );
  AND2X2 U2518 ( .A(\data_in<10> ), .B(n1601), .Y(n2687) );
  INVX1 U2519 ( .A(n2687), .Y(n2688) );
  AND2X2 U2520 ( .A(\data_in<11> ), .B(n1601), .Y(n2689) );
  INVX1 U2521 ( .A(n2689), .Y(n2690) );
  AND2X2 U2522 ( .A(\data_in<12> ), .B(n1601), .Y(n2691) );
  INVX1 U2523 ( .A(n2691), .Y(n2692) );
  AND2X2 U2524 ( .A(\data_in<13> ), .B(n1601), .Y(n2693) );
  INVX1 U2525 ( .A(n2693), .Y(n2694) );
  AND2X2 U2526 ( .A(\data_in<14> ), .B(n1601), .Y(n2695) );
  INVX1 U2527 ( .A(n2695), .Y(n2696) );
  AND2X2 U2528 ( .A(\data_in<15> ), .B(n1601), .Y(n2697) );
  INVX1 U2529 ( .A(n2697), .Y(n2698) );
  AND2X2 U2530 ( .A(\data_in<8> ), .B(n1603), .Y(n2699) );
  INVX1 U2531 ( .A(n2699), .Y(n2700) );
  AND2X2 U2532 ( .A(\data_in<9> ), .B(n1603), .Y(n2701) );
  INVX1 U2533 ( .A(n2701), .Y(n2702) );
  AND2X2 U2534 ( .A(\data_in<10> ), .B(n1603), .Y(n2703) );
  INVX1 U2535 ( .A(n2703), .Y(n2704) );
  AND2X2 U2536 ( .A(\data_in<11> ), .B(n1603), .Y(n2705) );
  INVX1 U2537 ( .A(n2705), .Y(n2706) );
  AND2X2 U2538 ( .A(\data_in<12> ), .B(n1603), .Y(n2707) );
  INVX1 U2539 ( .A(n2707), .Y(n2708) );
  AND2X2 U2540 ( .A(\data_in<13> ), .B(n1603), .Y(n2709) );
  INVX1 U2541 ( .A(n2709), .Y(n2710) );
  AND2X2 U2542 ( .A(\data_in<14> ), .B(n1603), .Y(n2711) );
  INVX1 U2543 ( .A(n2711), .Y(n2712) );
  AND2X2 U2544 ( .A(\data_in<15> ), .B(n1603), .Y(n2713) );
  INVX1 U2545 ( .A(n2713), .Y(n2714) );
  AND2X2 U2546 ( .A(\data_in<8> ), .B(n1607), .Y(n2715) );
  INVX1 U2547 ( .A(n2715), .Y(n2716) );
  AND2X2 U2548 ( .A(\data_in<9> ), .B(n1607), .Y(n2717) );
  INVX1 U2549 ( .A(n2717), .Y(n2718) );
  AND2X2 U2550 ( .A(\data_in<10> ), .B(n1607), .Y(n2719) );
  INVX1 U2551 ( .A(n2719), .Y(n2720) );
  AND2X2 U2552 ( .A(\data_in<11> ), .B(n1607), .Y(n2721) );
  INVX1 U2553 ( .A(n2721), .Y(n2722) );
  AND2X2 U2554 ( .A(\data_in<12> ), .B(n1607), .Y(n2723) );
  INVX1 U2555 ( .A(n2723), .Y(n2724) );
  AND2X2 U2556 ( .A(\data_in<13> ), .B(n1607), .Y(n2725) );
  INVX1 U2557 ( .A(n2725), .Y(n2726) );
  AND2X2 U2558 ( .A(\data_in<14> ), .B(n1607), .Y(n2727) );
  INVX1 U2559 ( .A(n2727), .Y(n2728) );
  AND2X2 U2560 ( .A(\data_in<15> ), .B(n1607), .Y(n2729) );
  INVX1 U2561 ( .A(n2729), .Y(n2730) );
  AND2X2 U2562 ( .A(\data_in<8> ), .B(n1609), .Y(n2731) );
  INVX1 U2563 ( .A(n2731), .Y(n2732) );
  AND2X2 U2564 ( .A(\data_in<9> ), .B(n1609), .Y(n2733) );
  INVX1 U2565 ( .A(n2733), .Y(n2734) );
  AND2X2 U2566 ( .A(\data_in<10> ), .B(n1609), .Y(n2735) );
  INVX1 U2567 ( .A(n2735), .Y(n2736) );
  AND2X2 U2568 ( .A(\data_in<11> ), .B(n1609), .Y(n2737) );
  INVX1 U2569 ( .A(n2737), .Y(n2738) );
  AND2X2 U2570 ( .A(\data_in<12> ), .B(n1609), .Y(n2739) );
  INVX1 U2571 ( .A(n2739), .Y(n2740) );
  AND2X2 U2572 ( .A(\data_in<13> ), .B(n1609), .Y(n2741) );
  INVX1 U2573 ( .A(n2741), .Y(n2742) );
  AND2X2 U2574 ( .A(\data_in<14> ), .B(n1609), .Y(n2743) );
  INVX1 U2575 ( .A(n2743), .Y(n2744) );
  AND2X2 U2576 ( .A(\data_in<15> ), .B(n1609), .Y(n2745) );
  INVX1 U2577 ( .A(n2745), .Y(n2746) );
  AND2X2 U2578 ( .A(\data_in<8> ), .B(n1611), .Y(n2747) );
  INVX1 U2579 ( .A(n2747), .Y(n2748) );
  AND2X2 U2580 ( .A(\data_in<9> ), .B(n1611), .Y(n2749) );
  INVX1 U2581 ( .A(n2749), .Y(n2750) );
  AND2X2 U2582 ( .A(\data_in<10> ), .B(n1611), .Y(n2751) );
  INVX1 U2583 ( .A(n2751), .Y(n2752) );
  AND2X2 U2584 ( .A(\data_in<11> ), .B(n1611), .Y(n2753) );
  INVX1 U2585 ( .A(n2753), .Y(n2754) );
  AND2X2 U2586 ( .A(\data_in<12> ), .B(n1611), .Y(n2755) );
  INVX1 U2587 ( .A(n2755), .Y(n2756) );
  AND2X2 U2588 ( .A(\data_in<13> ), .B(n1611), .Y(n2757) );
  INVX1 U2589 ( .A(n2757), .Y(n2758) );
  AND2X2 U2590 ( .A(\data_in<14> ), .B(n1611), .Y(n2759) );
  INVX1 U2591 ( .A(n2759), .Y(n2760) );
  AND2X2 U2592 ( .A(\data_in<15> ), .B(n1611), .Y(n2761) );
  INVX1 U2593 ( .A(n2761), .Y(n2762) );
  AND2X2 U2594 ( .A(\data_in<8> ), .B(n1615), .Y(n2763) );
  INVX1 U2595 ( .A(n2763), .Y(n2764) );
  AND2X2 U2596 ( .A(\data_in<9> ), .B(n1615), .Y(n2765) );
  INVX1 U2597 ( .A(n2765), .Y(n2766) );
  AND2X2 U2598 ( .A(\data_in<10> ), .B(n1615), .Y(n2767) );
  INVX1 U2599 ( .A(n2767), .Y(n2768) );
  AND2X2 U2600 ( .A(\data_in<11> ), .B(n1615), .Y(n2769) );
  INVX1 U2601 ( .A(n2769), .Y(n2770) );
  AND2X2 U2602 ( .A(\data_in<12> ), .B(n1615), .Y(n2771) );
  INVX1 U2603 ( .A(n2771), .Y(n2772) );
  AND2X2 U2604 ( .A(\data_in<13> ), .B(n1615), .Y(n2773) );
  INVX1 U2605 ( .A(n2773), .Y(n2774) );
  AND2X2 U2606 ( .A(\data_in<14> ), .B(n1615), .Y(n2775) );
  INVX1 U2607 ( .A(n2775), .Y(n2776) );
  AND2X2 U2608 ( .A(\data_in<15> ), .B(n1615), .Y(n2777) );
  INVX1 U2609 ( .A(n2777), .Y(n2778) );
  AND2X2 U2610 ( .A(\data_in<8> ), .B(n1617), .Y(n2779) );
  INVX1 U2611 ( .A(n2779), .Y(n2780) );
  AND2X2 U2612 ( .A(\data_in<9> ), .B(n1617), .Y(n2781) );
  INVX1 U2613 ( .A(n2781), .Y(n2782) );
  AND2X2 U2614 ( .A(\data_in<10> ), .B(n1617), .Y(n2783) );
  INVX1 U2615 ( .A(n2783), .Y(n2784) );
  AND2X2 U2616 ( .A(\data_in<11> ), .B(n1617), .Y(n2785) );
  INVX1 U2617 ( .A(n2785), .Y(n2786) );
  AND2X2 U2618 ( .A(\data_in<12> ), .B(n1617), .Y(n2787) );
  INVX1 U2619 ( .A(n2787), .Y(n2788) );
  AND2X2 U2620 ( .A(\data_in<13> ), .B(n1617), .Y(n2789) );
  INVX1 U2621 ( .A(n2789), .Y(n2790) );
  AND2X2 U2622 ( .A(\data_in<14> ), .B(n1617), .Y(n2791) );
  INVX1 U2623 ( .A(n2791), .Y(n2792) );
  AND2X2 U2624 ( .A(\data_in<15> ), .B(n1617), .Y(n2793) );
  INVX1 U2625 ( .A(n2793), .Y(n2794) );
  AND2X2 U2626 ( .A(\data_in<8> ), .B(n1619), .Y(n2795) );
  INVX1 U2627 ( .A(n2795), .Y(n2796) );
  AND2X2 U2628 ( .A(\data_in<9> ), .B(n1619), .Y(n2797) );
  INVX1 U2629 ( .A(n2797), .Y(n2798) );
  AND2X2 U2630 ( .A(\data_in<10> ), .B(n1619), .Y(n2799) );
  INVX1 U2631 ( .A(n2799), .Y(n2800) );
  AND2X2 U2632 ( .A(\data_in<11> ), .B(n1619), .Y(n2801) );
  INVX1 U2633 ( .A(n2801), .Y(n2802) );
  AND2X2 U2634 ( .A(\data_in<12> ), .B(n1619), .Y(n2803) );
  INVX1 U2635 ( .A(n2803), .Y(n2804) );
  AND2X2 U2636 ( .A(\data_in<13> ), .B(n1619), .Y(n2805) );
  INVX1 U2637 ( .A(n2805), .Y(n2806) );
  AND2X2 U2638 ( .A(\data_in<14> ), .B(n1619), .Y(n2807) );
  INVX1 U2639 ( .A(n2807), .Y(n2808) );
  AND2X2 U2640 ( .A(\data_in<15> ), .B(n1619), .Y(n2809) );
  INVX1 U2641 ( .A(n2809), .Y(n2810) );
  AND2X2 U2642 ( .A(\data_in<8> ), .B(n3844), .Y(n2811) );
  INVX1 U2643 ( .A(n2811), .Y(n2812) );
  AND2X2 U2644 ( .A(\data_in<9> ), .B(n3844), .Y(n2813) );
  INVX1 U2645 ( .A(n2813), .Y(n2814) );
  AND2X2 U2646 ( .A(\data_in<10> ), .B(n3844), .Y(n2815) );
  INVX1 U2647 ( .A(n2815), .Y(n2816) );
  AND2X2 U2648 ( .A(\data_in<11> ), .B(n3844), .Y(n2817) );
  INVX1 U2649 ( .A(n2817), .Y(n2818) );
  AND2X2 U2650 ( .A(\data_in<12> ), .B(n3844), .Y(n2819) );
  INVX1 U2651 ( .A(n2819), .Y(n2820) );
  AND2X2 U2652 ( .A(\data_in<13> ), .B(n3844), .Y(n2821) );
  INVX1 U2653 ( .A(n2821), .Y(n2822) );
  AND2X2 U2654 ( .A(\data_in<14> ), .B(n3844), .Y(n2823) );
  INVX1 U2655 ( .A(n2823), .Y(n2824) );
  AND2X2 U2656 ( .A(\data_in<15> ), .B(n3844), .Y(n2825) );
  INVX1 U2657 ( .A(n2825), .Y(n2826) );
  AND2X2 U2658 ( .A(\data_in<8> ), .B(n1622), .Y(n2827) );
  INVX1 U2659 ( .A(n2827), .Y(n2828) );
  AND2X2 U2660 ( .A(\data_in<9> ), .B(n17), .Y(n2829) );
  INVX1 U2661 ( .A(n2829), .Y(n2830) );
  AND2X2 U2662 ( .A(\data_in<10> ), .B(n17), .Y(n2831) );
  INVX1 U2663 ( .A(n2831), .Y(n2832) );
  AND2X2 U2664 ( .A(\data_in<11> ), .B(n1622), .Y(n2833) );
  INVX1 U2665 ( .A(n2833), .Y(n2834) );
  AND2X2 U2666 ( .A(\data_in<12> ), .B(n1622), .Y(n2835) );
  INVX1 U2667 ( .A(n2835), .Y(n2836) );
  AND2X2 U2668 ( .A(\data_in<13> ), .B(n17), .Y(n2837) );
  INVX1 U2669 ( .A(n2837), .Y(n2838) );
  AND2X2 U2670 ( .A(\data_in<14> ), .B(n17), .Y(n2839) );
  INVX1 U2671 ( .A(n2839), .Y(n2840) );
  AND2X2 U2672 ( .A(\data_in<15> ), .B(n1622), .Y(n2841) );
  INVX1 U2673 ( .A(n2841), .Y(n2842) );
  AND2X2 U2674 ( .A(\data_in<8> ), .B(n1624), .Y(n2843) );
  INVX1 U2675 ( .A(n2843), .Y(n2844) );
  AND2X2 U2676 ( .A(\data_in<9> ), .B(n1624), .Y(n2845) );
  INVX1 U2677 ( .A(n2845), .Y(n2846) );
  AND2X2 U2678 ( .A(\data_in<10> ), .B(n1624), .Y(n2847) );
  INVX1 U2679 ( .A(n2847), .Y(n2848) );
  AND2X2 U2680 ( .A(\data_in<11> ), .B(n1624), .Y(n2849) );
  INVX1 U2681 ( .A(n2849), .Y(n2850) );
  AND2X2 U2682 ( .A(\data_in<12> ), .B(n1624), .Y(n2851) );
  INVX1 U2683 ( .A(n2851), .Y(n2852) );
  AND2X2 U2684 ( .A(\data_in<13> ), .B(n1624), .Y(n2853) );
  INVX1 U2685 ( .A(n2853), .Y(n2854) );
  AND2X2 U2686 ( .A(\data_in<14> ), .B(n1624), .Y(n2855) );
  INVX1 U2687 ( .A(n2855), .Y(n2856) );
  AND2X2 U2688 ( .A(\data_in<15> ), .B(n1624), .Y(n2857) );
  INVX1 U2689 ( .A(n2857), .Y(n2858) );
  AND2X2 U2690 ( .A(\data_in<8> ), .B(n6437), .Y(n2859) );
  INVX1 U2691 ( .A(n2859), .Y(n2860) );
  AND2X2 U2692 ( .A(\data_in<9> ), .B(n6437), .Y(n2861) );
  INVX1 U2693 ( .A(n2861), .Y(n2862) );
  AND2X2 U2694 ( .A(\data_in<10> ), .B(n6437), .Y(n2863) );
  INVX1 U2695 ( .A(n2863), .Y(n2864) );
  AND2X2 U2696 ( .A(\data_in<11> ), .B(n6437), .Y(n2865) );
  INVX1 U2697 ( .A(n2865), .Y(n2866) );
  AND2X2 U2698 ( .A(\data_in<12> ), .B(n6437), .Y(n2867) );
  INVX1 U2699 ( .A(n2867), .Y(n2868) );
  AND2X2 U2700 ( .A(\data_in<13> ), .B(n6437), .Y(n2869) );
  INVX1 U2701 ( .A(n2869), .Y(n2870) );
  AND2X2 U2702 ( .A(\data_in<14> ), .B(n6437), .Y(n2871) );
  INVX1 U2703 ( .A(n2871), .Y(n2872) );
  AND2X2 U2704 ( .A(\data_in<15> ), .B(n6437), .Y(n2873) );
  INVX1 U2705 ( .A(n2873), .Y(n2874) );
  AND2X2 U2706 ( .A(\data_in<8> ), .B(n1627), .Y(n2875) );
  INVX1 U2707 ( .A(n2875), .Y(n2876) );
  AND2X2 U2708 ( .A(\data_in<9> ), .B(n1627), .Y(n2877) );
  INVX1 U2709 ( .A(n2877), .Y(n2878) );
  AND2X2 U2710 ( .A(\data_in<10> ), .B(n1627), .Y(n2879) );
  INVX1 U2711 ( .A(n2879), .Y(n2880) );
  AND2X2 U2712 ( .A(\data_in<11> ), .B(n1627), .Y(n2881) );
  INVX1 U2713 ( .A(n2881), .Y(n2882) );
  AND2X2 U2714 ( .A(\data_in<12> ), .B(n1627), .Y(n2883) );
  INVX1 U2715 ( .A(n2883), .Y(n2884) );
  AND2X2 U2716 ( .A(\data_in<13> ), .B(n1627), .Y(n2885) );
  INVX1 U2717 ( .A(n2885), .Y(n2886) );
  AND2X2 U2718 ( .A(\data_in<14> ), .B(n1627), .Y(n2887) );
  INVX1 U2719 ( .A(n2887), .Y(n2888) );
  AND2X2 U2720 ( .A(\data_in<15> ), .B(n1627), .Y(n2889) );
  INVX1 U2721 ( .A(n2889), .Y(n2890) );
  AND2X2 U2722 ( .A(\data_in<8> ), .B(n1629), .Y(n2891) );
  INVX1 U2723 ( .A(n2891), .Y(n2892) );
  AND2X2 U2724 ( .A(\data_in<9> ), .B(n1629), .Y(n2893) );
  INVX1 U2725 ( .A(n2893), .Y(n2894) );
  AND2X2 U2726 ( .A(\data_in<10> ), .B(n1629), .Y(n2895) );
  INVX1 U2727 ( .A(n2895), .Y(n2896) );
  AND2X2 U2728 ( .A(\data_in<11> ), .B(n1629), .Y(n2897) );
  INVX1 U2729 ( .A(n2897), .Y(n2898) );
  AND2X2 U2730 ( .A(\data_in<12> ), .B(n1629), .Y(n2899) );
  INVX1 U2731 ( .A(n2899), .Y(n2900) );
  AND2X2 U2732 ( .A(\data_in<13> ), .B(n1629), .Y(n2901) );
  INVX1 U2733 ( .A(n2901), .Y(n2902) );
  AND2X2 U2734 ( .A(\data_in<14> ), .B(n1629), .Y(n2903) );
  INVX1 U2735 ( .A(n2903), .Y(n2904) );
  AND2X2 U2736 ( .A(\data_in<15> ), .B(n1629), .Y(n2905) );
  INVX1 U2737 ( .A(n2905), .Y(n2906) );
  AND2X2 U2738 ( .A(\data_in<8> ), .B(n1631), .Y(n2907) );
  INVX1 U2739 ( .A(n2907), .Y(n2908) );
  AND2X2 U2740 ( .A(\data_in<9> ), .B(n1631), .Y(n2909) );
  INVX1 U2741 ( .A(n2909), .Y(n2910) );
  AND2X2 U2742 ( .A(\data_in<10> ), .B(n1631), .Y(n2911) );
  INVX1 U2743 ( .A(n2911), .Y(n2912) );
  AND2X2 U2744 ( .A(\data_in<11> ), .B(n1631), .Y(n2913) );
  INVX1 U2745 ( .A(n2913), .Y(n2914) );
  AND2X2 U2746 ( .A(\data_in<12> ), .B(n1631), .Y(n2915) );
  INVX1 U2747 ( .A(n2915), .Y(n2916) );
  AND2X2 U2748 ( .A(\data_in<13> ), .B(n1631), .Y(n2917) );
  INVX1 U2749 ( .A(n2917), .Y(n2918) );
  AND2X2 U2750 ( .A(\data_in<14> ), .B(n1631), .Y(n2919) );
  INVX1 U2751 ( .A(n2919), .Y(n2920) );
  AND2X2 U2752 ( .A(\data_in<15> ), .B(n1631), .Y(n2921) );
  INVX1 U2753 ( .A(n2921), .Y(n2922) );
  AND2X2 U2754 ( .A(\data_in<8> ), .B(n1633), .Y(n2923) );
  INVX1 U2755 ( .A(n2923), .Y(n2924) );
  AND2X2 U2756 ( .A(\data_in<9> ), .B(n1633), .Y(n2925) );
  INVX1 U2757 ( .A(n2925), .Y(n2926) );
  AND2X2 U2758 ( .A(\data_in<10> ), .B(n1633), .Y(n2927) );
  INVX1 U2759 ( .A(n2927), .Y(n2928) );
  AND2X2 U2760 ( .A(\data_in<11> ), .B(n1633), .Y(n2929) );
  INVX1 U2761 ( .A(n2929), .Y(n2930) );
  AND2X2 U2762 ( .A(\data_in<12> ), .B(n1633), .Y(n2931) );
  INVX1 U2763 ( .A(n2931), .Y(n2932) );
  AND2X2 U2764 ( .A(\data_in<13> ), .B(n1633), .Y(n2933) );
  INVX1 U2765 ( .A(n2933), .Y(n2934) );
  AND2X2 U2766 ( .A(\data_in<14> ), .B(n1633), .Y(n2935) );
  INVX1 U2767 ( .A(n2935), .Y(n2936) );
  AND2X2 U2768 ( .A(\data_in<15> ), .B(n1633), .Y(n2937) );
  INVX1 U2769 ( .A(n2937), .Y(n2938) );
  AND2X2 U2770 ( .A(\data_in<8> ), .B(n1638), .Y(n2939) );
  INVX1 U2771 ( .A(n2939), .Y(n2940) );
  AND2X2 U2772 ( .A(\data_in<9> ), .B(n1638), .Y(n2941) );
  INVX1 U2773 ( .A(n2941), .Y(n2942) );
  AND2X2 U2774 ( .A(\data_in<10> ), .B(n1638), .Y(n2943) );
  INVX1 U2775 ( .A(n2943), .Y(n2944) );
  AND2X2 U2776 ( .A(\data_in<11> ), .B(n1638), .Y(n2945) );
  INVX1 U2777 ( .A(n2945), .Y(n2946) );
  AND2X2 U2778 ( .A(\data_in<12> ), .B(n1638), .Y(n2947) );
  INVX1 U2779 ( .A(n2947), .Y(n2948) );
  AND2X2 U2780 ( .A(\data_in<13> ), .B(n1638), .Y(n2949) );
  INVX1 U2781 ( .A(n2949), .Y(n2950) );
  AND2X2 U2782 ( .A(\data_in<14> ), .B(n1638), .Y(n2951) );
  INVX1 U2783 ( .A(n2951), .Y(n2952) );
  AND2X2 U2784 ( .A(\data_in<15> ), .B(n1638), .Y(n2953) );
  INVX1 U2785 ( .A(n2953), .Y(n2954) );
  AND2X2 U2786 ( .A(\data_in<8> ), .B(n1640), .Y(n2955) );
  INVX1 U2787 ( .A(n2955), .Y(n2956) );
  AND2X2 U2788 ( .A(\data_in<9> ), .B(n1640), .Y(n2957) );
  INVX1 U2789 ( .A(n2957), .Y(n2958) );
  AND2X2 U2790 ( .A(\data_in<10> ), .B(n1640), .Y(n2959) );
  INVX1 U2791 ( .A(n2959), .Y(n2960) );
  AND2X2 U2792 ( .A(\data_in<11> ), .B(n1640), .Y(n2961) );
  INVX1 U2793 ( .A(n2961), .Y(n2962) );
  AND2X2 U2794 ( .A(\data_in<12> ), .B(n1640), .Y(n2963) );
  INVX1 U2795 ( .A(n2963), .Y(n2964) );
  AND2X2 U2796 ( .A(\data_in<13> ), .B(n1640), .Y(n2965) );
  INVX1 U2797 ( .A(n2965), .Y(n2966) );
  AND2X2 U2798 ( .A(\data_in<14> ), .B(n1640), .Y(n2967) );
  INVX1 U2799 ( .A(n2967), .Y(n2968) );
  AND2X2 U2800 ( .A(\data_in<15> ), .B(n1640), .Y(n2969) );
  INVX1 U2801 ( .A(n2969), .Y(n2970) );
  AND2X2 U2802 ( .A(\data_in<8> ), .B(n1642), .Y(n2971) );
  INVX1 U2803 ( .A(n2971), .Y(n2972) );
  AND2X2 U2804 ( .A(\data_in<9> ), .B(n1642), .Y(n2973) );
  INVX1 U2805 ( .A(n2973), .Y(n2974) );
  AND2X2 U2806 ( .A(\data_in<11> ), .B(n1642), .Y(n2975) );
  INVX1 U2807 ( .A(n2975), .Y(n2976) );
  AND2X2 U2808 ( .A(\data_in<12> ), .B(n1642), .Y(n2977) );
  INVX1 U2809 ( .A(n2977), .Y(n2978) );
  AND2X2 U2810 ( .A(\data_in<14> ), .B(n1642), .Y(n2979) );
  INVX1 U2811 ( .A(n2979), .Y(n2980) );
  AND2X2 U2812 ( .A(\data_in<15> ), .B(n1642), .Y(n2981) );
  INVX1 U2813 ( .A(n2981), .Y(n2982) );
  AND2X2 U2814 ( .A(\data_in<8> ), .B(n1644), .Y(n2983) );
  INVX1 U2815 ( .A(n2983), .Y(n2984) );
  AND2X2 U2816 ( .A(\data_in<9> ), .B(n1644), .Y(n2985) );
  INVX1 U2817 ( .A(n2985), .Y(n2986) );
  AND2X2 U2818 ( .A(\data_in<10> ), .B(n1644), .Y(n2987) );
  INVX1 U2819 ( .A(n2987), .Y(n2988) );
  AND2X2 U2820 ( .A(\data_in<11> ), .B(n1644), .Y(n2989) );
  INVX1 U2821 ( .A(n2989), .Y(n2990) );
  AND2X2 U2822 ( .A(\data_in<12> ), .B(n1644), .Y(n2991) );
  INVX1 U2823 ( .A(n2991), .Y(n2992) );
  AND2X2 U2824 ( .A(\data_in<13> ), .B(n1644), .Y(n2993) );
  INVX1 U2825 ( .A(n2993), .Y(n2994) );
  AND2X2 U2826 ( .A(\data_in<8> ), .B(n1646), .Y(n2995) );
  INVX1 U2827 ( .A(n2995), .Y(n2996) );
  AND2X2 U2828 ( .A(\data_in<9> ), .B(n1646), .Y(n2997) );
  INVX1 U2829 ( .A(n2997), .Y(n2998) );
  AND2X2 U2830 ( .A(\data_in<11> ), .B(n1646), .Y(n2999) );
  INVX1 U2831 ( .A(n2999), .Y(n3000) );
  AND2X2 U2832 ( .A(\data_in<12> ), .B(n1646), .Y(n3001) );
  INVX1 U2833 ( .A(n3001), .Y(n3002) );
  AND2X2 U2834 ( .A(\data_in<14> ), .B(n1646), .Y(n3003) );
  INVX1 U2835 ( .A(n3003), .Y(n3004) );
  AND2X2 U2836 ( .A(\data_in<15> ), .B(n1646), .Y(n3005) );
  INVX1 U2837 ( .A(n3005), .Y(n3006) );
  INVX1 U2838 ( .A(n6018), .Y(n3007) );
  INVX1 U2839 ( .A(n6164), .Y(n3008) );
  AND2X2 U2840 ( .A(n5859), .B(n537), .Y(n3009) );
  INVX1 U2841 ( .A(n3009), .Y(n3010) );
  AND2X2 U2842 ( .A(n5938), .B(n542), .Y(n3011) );
  INVX1 U2843 ( .A(n3011), .Y(n3012) );
  AND2X2 U2844 ( .A(n6090), .B(n543), .Y(n3013) );
  INVX1 U2845 ( .A(n3013), .Y(n3014) );
  INVX1 U2846 ( .A(n5805), .Y(n3015) );
  INVX1 U2847 ( .A(n5806), .Y(n3016) );
  INVX1 U2848 ( .A(n5991), .Y(n3017) );
  INVX1 U2849 ( .A(n5992), .Y(n3018) );
  INVX1 U2850 ( .A(n6065), .Y(n3019) );
  INVX1 U2851 ( .A(n6066), .Y(n3020) );
  INVX1 U2852 ( .A(n6291), .Y(n3021) );
  INVX1 U2853 ( .A(n6292), .Y(n3022) );
  AND2X2 U2854 ( .A(n592), .B(n4106), .Y(n3023) );
  INVX1 U2855 ( .A(n3023), .Y(n3024) );
  AND2X2 U2856 ( .A(n921), .B(n5784), .Y(n3025) );
  INVX1 U2857 ( .A(n3025), .Y(n3026) );
  AND2X2 U2858 ( .A(n927), .B(n954), .Y(n3027) );
  INVX1 U2859 ( .A(n3027), .Y(n3028) );
  AND2X2 U2860 ( .A(n931), .B(n960), .Y(n3029) );
  INVX1 U2861 ( .A(n3029), .Y(n3030) );
  OR2X2 U2862 ( .A(n5897), .B(n5898), .Y(n3031) );
  AND2X2 U2863 ( .A(n915), .B(n76), .Y(n3032) );
  INVX1 U2864 ( .A(n3032), .Y(n3033) );
  OR2X2 U2865 ( .A(\addr<12> ), .B(\addr<9> ), .Y(n3034) );
  OR2X2 U2866 ( .A(n6033), .B(n6034), .Y(n3035) );
  OR2X2 U2867 ( .A(n6050), .B(n6051), .Y(n3036) );
  AND2X2 U2868 ( .A(\data_in<0> ), .B(n1529), .Y(n3037) );
  INVX1 U2869 ( .A(n3037), .Y(n3038) );
  AND2X2 U2870 ( .A(\data_in<1> ), .B(n1529), .Y(n3039) );
  INVX1 U2871 ( .A(n3039), .Y(n3040) );
  AND2X2 U2872 ( .A(\data_in<2> ), .B(n1529), .Y(n3041) );
  INVX1 U2873 ( .A(n3041), .Y(n3042) );
  AND2X2 U2874 ( .A(\data_in<3> ), .B(n1529), .Y(n3043) );
  INVX1 U2875 ( .A(n3043), .Y(n3044) );
  AND2X2 U2876 ( .A(\data_in<4> ), .B(n1529), .Y(n3045) );
  INVX1 U2877 ( .A(n3045), .Y(n3046) );
  AND2X2 U2878 ( .A(\data_in<5> ), .B(n1529), .Y(n3047) );
  INVX1 U2879 ( .A(n3047), .Y(n3048) );
  AND2X2 U2880 ( .A(\data_in<6> ), .B(n1529), .Y(n3049) );
  INVX1 U2881 ( .A(n3049), .Y(n3050) );
  AND2X2 U2882 ( .A(\data_in<7> ), .B(n1529), .Y(n3051) );
  INVX1 U2883 ( .A(n3051), .Y(n3052) );
  AND2X2 U2884 ( .A(\data_in<0> ), .B(n1531), .Y(n3053) );
  INVX1 U2885 ( .A(n3053), .Y(n3054) );
  AND2X2 U2886 ( .A(\data_in<1> ), .B(n1531), .Y(n3055) );
  INVX1 U2887 ( .A(n3055), .Y(n3056) );
  AND2X2 U2888 ( .A(\data_in<2> ), .B(n1531), .Y(n3057) );
  INVX1 U2889 ( .A(n3057), .Y(n3058) );
  AND2X2 U2890 ( .A(\data_in<3> ), .B(n1531), .Y(n3059) );
  INVX1 U2891 ( .A(n3059), .Y(n3060) );
  AND2X2 U2892 ( .A(\data_in<4> ), .B(n1531), .Y(n3061) );
  INVX1 U2893 ( .A(n3061), .Y(n3062) );
  AND2X2 U2894 ( .A(\data_in<5> ), .B(n1531), .Y(n3063) );
  INVX1 U2895 ( .A(n3063), .Y(n3064) );
  AND2X2 U2896 ( .A(\data_in<6> ), .B(n1531), .Y(n3065) );
  INVX1 U2897 ( .A(n3065), .Y(n3066) );
  AND2X2 U2898 ( .A(\data_in<7> ), .B(n1531), .Y(n3067) );
  INVX1 U2899 ( .A(n3067), .Y(n3068) );
  AND2X2 U2900 ( .A(\data_in<0> ), .B(n1533), .Y(n3069) );
  INVX1 U2901 ( .A(n3069), .Y(n3070) );
  AND2X2 U2902 ( .A(\data_in<1> ), .B(n1533), .Y(n3071) );
  INVX1 U2903 ( .A(n3071), .Y(n3072) );
  AND2X2 U2904 ( .A(\data_in<2> ), .B(n1533), .Y(n3073) );
  INVX1 U2905 ( .A(n3073), .Y(n3074) );
  AND2X2 U2906 ( .A(\data_in<3> ), .B(n1533), .Y(n3075) );
  INVX1 U2907 ( .A(n3075), .Y(n3076) );
  AND2X2 U2908 ( .A(\data_in<4> ), .B(n1533), .Y(n3077) );
  INVX1 U2909 ( .A(n3077), .Y(n3078) );
  AND2X2 U2910 ( .A(\data_in<5> ), .B(n1533), .Y(n3079) );
  INVX1 U2911 ( .A(n3079), .Y(n3080) );
  AND2X2 U2912 ( .A(\data_in<6> ), .B(n1533), .Y(n3081) );
  INVX1 U2913 ( .A(n3081), .Y(n3082) );
  AND2X2 U2914 ( .A(\data_in<7> ), .B(n1533), .Y(n3083) );
  INVX1 U2915 ( .A(n3083), .Y(n3084) );
  AND2X2 U2916 ( .A(\data_in<0> ), .B(n1535), .Y(n3085) );
  INVX1 U2917 ( .A(n3085), .Y(n3086) );
  AND2X2 U2918 ( .A(\data_in<1> ), .B(n1535), .Y(n3087) );
  INVX1 U2919 ( .A(n3087), .Y(n3088) );
  AND2X2 U2920 ( .A(\data_in<2> ), .B(n1535), .Y(n3089) );
  INVX1 U2921 ( .A(n3089), .Y(n3090) );
  AND2X2 U2922 ( .A(\data_in<3> ), .B(n1535), .Y(n3091) );
  INVX1 U2923 ( .A(n3091), .Y(n3092) );
  AND2X2 U2924 ( .A(\data_in<4> ), .B(n1535), .Y(n3093) );
  INVX1 U2925 ( .A(n3093), .Y(n3094) );
  AND2X2 U2926 ( .A(\data_in<5> ), .B(n1535), .Y(n3095) );
  INVX1 U2927 ( .A(n3095), .Y(n3096) );
  AND2X2 U2928 ( .A(\data_in<6> ), .B(n1535), .Y(n3097) );
  INVX1 U2929 ( .A(n3097), .Y(n3098) );
  AND2X2 U2930 ( .A(\data_in<7> ), .B(n1535), .Y(n3099) );
  INVX1 U2931 ( .A(n3099), .Y(n3100) );
  AND2X2 U2932 ( .A(\data_in<0> ), .B(n1537), .Y(n3101) );
  INVX1 U2933 ( .A(n3101), .Y(n3102) );
  AND2X2 U2934 ( .A(\data_in<1> ), .B(n1537), .Y(n3103) );
  INVX1 U2935 ( .A(n3103), .Y(n3104) );
  AND2X2 U2936 ( .A(\data_in<2> ), .B(n1537), .Y(n3105) );
  INVX1 U2937 ( .A(n3105), .Y(n3106) );
  AND2X2 U2938 ( .A(\data_in<3> ), .B(n1537), .Y(n3107) );
  INVX1 U2939 ( .A(n3107), .Y(n3108) );
  AND2X2 U2940 ( .A(\data_in<4> ), .B(n1537), .Y(n3109) );
  INVX1 U2941 ( .A(n3109), .Y(n3110) );
  AND2X2 U2942 ( .A(\data_in<5> ), .B(n1537), .Y(n3111) );
  INVX1 U2943 ( .A(n3111), .Y(n3112) );
  AND2X2 U2944 ( .A(\data_in<6> ), .B(n1537), .Y(n3113) );
  INVX1 U2945 ( .A(n3113), .Y(n3114) );
  AND2X2 U2946 ( .A(\data_in<7> ), .B(n1537), .Y(n3115) );
  INVX1 U2947 ( .A(n3115), .Y(n3116) );
  AND2X2 U2948 ( .A(\data_in<0> ), .B(n1539), .Y(n3117) );
  INVX1 U2949 ( .A(n3117), .Y(n3118) );
  AND2X2 U2950 ( .A(\data_in<1> ), .B(n1539), .Y(n3119) );
  INVX1 U2951 ( .A(n3119), .Y(n3120) );
  AND2X2 U2952 ( .A(\data_in<2> ), .B(n1539), .Y(n3121) );
  INVX1 U2953 ( .A(n3121), .Y(n3122) );
  AND2X2 U2954 ( .A(\data_in<3> ), .B(n1539), .Y(n3123) );
  INVX1 U2955 ( .A(n3123), .Y(n3124) );
  AND2X2 U2956 ( .A(\data_in<4> ), .B(n1539), .Y(n3125) );
  INVX1 U2957 ( .A(n3125), .Y(n3126) );
  AND2X2 U2958 ( .A(\data_in<5> ), .B(n1539), .Y(n3127) );
  INVX1 U2959 ( .A(n3127), .Y(n3128) );
  AND2X2 U2960 ( .A(\data_in<6> ), .B(n1539), .Y(n3129) );
  INVX1 U2961 ( .A(n3129), .Y(n3130) );
  AND2X2 U2962 ( .A(\data_in<7> ), .B(n1539), .Y(n3131) );
  INVX1 U2963 ( .A(n3131), .Y(n3132) );
  AND2X2 U2964 ( .A(\data_in<0> ), .B(n5), .Y(n3133) );
  INVX1 U2965 ( .A(n3133), .Y(n3134) );
  AND2X2 U2966 ( .A(n672), .B(n4), .Y(n3135) );
  INVX1 U2967 ( .A(n3135), .Y(n3136) );
  AND2X2 U2968 ( .A(\data_in<2> ), .B(n1541), .Y(n3137) );
  INVX1 U2969 ( .A(n3137), .Y(n3138) );
  AND2X2 U2970 ( .A(\data_in<3> ), .B(n1541), .Y(n3139) );
  INVX1 U2971 ( .A(n3139), .Y(n3140) );
  AND2X2 U2972 ( .A(\data_in<4> ), .B(n5), .Y(n3141) );
  INVX1 U2973 ( .A(n3141), .Y(n3142) );
  AND2X2 U2974 ( .A(\data_in<5> ), .B(n5), .Y(n3143) );
  INVX1 U2975 ( .A(n3143), .Y(n3144) );
  AND2X2 U2976 ( .A(\data_in<6> ), .B(n1541), .Y(n3145) );
  INVX1 U2977 ( .A(n3145), .Y(n3146) );
  AND2X2 U2978 ( .A(\data_in<7> ), .B(n1541), .Y(n3147) );
  INVX1 U2979 ( .A(n3147), .Y(n3148) );
  AND2X2 U2980 ( .A(\mem<56><2> ), .B(n4984), .Y(n3149) );
  INVX1 U2981 ( .A(n3149), .Y(n3150) );
  AND2X2 U2982 ( .A(\mem<56><5> ), .B(n4985), .Y(n3151) );
  INVX1 U2983 ( .A(n3151), .Y(n3152) );
  AND2X2 U2984 ( .A(\data_in<0> ), .B(n1545), .Y(n3153) );
  INVX1 U2985 ( .A(n3153), .Y(n3154) );
  AND2X2 U2986 ( .A(\data_in<1> ), .B(n1545), .Y(n3155) );
  INVX1 U2987 ( .A(n3155), .Y(n3156) );
  AND2X2 U2988 ( .A(\data_in<2> ), .B(n1545), .Y(n3157) );
  INVX1 U2989 ( .A(n3157), .Y(n3158) );
  AND2X2 U2990 ( .A(\data_in<3> ), .B(n1545), .Y(n3159) );
  INVX1 U2991 ( .A(n3159), .Y(n3160) );
  AND2X2 U2992 ( .A(\data_in<4> ), .B(n1545), .Y(n3161) );
  INVX1 U2993 ( .A(n3161), .Y(n3162) );
  AND2X2 U2994 ( .A(\data_in<5> ), .B(n1545), .Y(n3163) );
  INVX1 U2995 ( .A(n3163), .Y(n3164) );
  AND2X2 U2996 ( .A(\data_in<6> ), .B(n1545), .Y(n3165) );
  INVX1 U2997 ( .A(n3165), .Y(n3166) );
  AND2X2 U2998 ( .A(\data_in<7> ), .B(n1545), .Y(n3167) );
  INVX1 U2999 ( .A(n3167), .Y(n3168) );
  AND2X2 U3000 ( .A(\data_in<0> ), .B(n1547), .Y(n3169) );
  INVX1 U3001 ( .A(n3169), .Y(n3170) );
  AND2X2 U3002 ( .A(\data_in<1> ), .B(n1547), .Y(n3171) );
  INVX1 U3003 ( .A(n3171), .Y(n3172) );
  AND2X2 U3004 ( .A(\data_in<2> ), .B(n1547), .Y(n3173) );
  INVX1 U3005 ( .A(n3173), .Y(n3174) );
  AND2X2 U3006 ( .A(\data_in<3> ), .B(n1547), .Y(n3175) );
  INVX1 U3007 ( .A(n3175), .Y(n3176) );
  AND2X2 U3008 ( .A(\data_in<4> ), .B(n1547), .Y(n3177) );
  INVX1 U3009 ( .A(n3177), .Y(n3178) );
  AND2X2 U3010 ( .A(\data_in<5> ), .B(n1547), .Y(n3179) );
  INVX1 U3011 ( .A(n3179), .Y(n3180) );
  AND2X2 U3012 ( .A(\data_in<6> ), .B(n1547), .Y(n3181) );
  INVX1 U3013 ( .A(n3181), .Y(n3182) );
  AND2X2 U3014 ( .A(\data_in<7> ), .B(n1547), .Y(n3183) );
  INVX1 U3015 ( .A(n3183), .Y(n3184) );
  AND2X2 U3016 ( .A(\data_in<0> ), .B(n1549), .Y(n3185) );
  INVX1 U3017 ( .A(n3185), .Y(n3186) );
  AND2X2 U3018 ( .A(\data_in<1> ), .B(n1549), .Y(n3187) );
  INVX1 U3019 ( .A(n3187), .Y(n3188) );
  AND2X2 U3020 ( .A(\data_in<2> ), .B(n1549), .Y(n3189) );
  INVX1 U3021 ( .A(n3189), .Y(n3190) );
  AND2X2 U3022 ( .A(\data_in<3> ), .B(n1549), .Y(n3191) );
  INVX1 U3023 ( .A(n3191), .Y(n3192) );
  AND2X2 U3024 ( .A(\data_in<4> ), .B(n1549), .Y(n3193) );
  INVX1 U3025 ( .A(n3193), .Y(n3194) );
  AND2X2 U3026 ( .A(\data_in<5> ), .B(n1549), .Y(n3195) );
  INVX1 U3027 ( .A(n3195), .Y(n3196) );
  AND2X2 U3028 ( .A(\data_in<6> ), .B(n1549), .Y(n3197) );
  INVX1 U3029 ( .A(n3197), .Y(n3198) );
  AND2X2 U3030 ( .A(\data_in<7> ), .B(n1549), .Y(n3199) );
  INVX1 U3031 ( .A(n3199), .Y(n3200) );
  AND2X2 U3032 ( .A(\data_in<0> ), .B(n1553), .Y(n3201) );
  INVX1 U3033 ( .A(n3201), .Y(n3202) );
  AND2X2 U3034 ( .A(\data_in<1> ), .B(n1553), .Y(n3203) );
  INVX1 U3035 ( .A(n3203), .Y(n3204) );
  AND2X2 U3036 ( .A(\data_in<2> ), .B(n1553), .Y(n3205) );
  INVX1 U3037 ( .A(n3205), .Y(n3206) );
  AND2X2 U3038 ( .A(\data_in<3> ), .B(n1553), .Y(n3207) );
  INVX1 U3039 ( .A(n3207), .Y(n3208) );
  AND2X2 U3040 ( .A(\data_in<4> ), .B(n1553), .Y(n3209) );
  INVX1 U3041 ( .A(n3209), .Y(n3210) );
  AND2X2 U3042 ( .A(\data_in<5> ), .B(n1553), .Y(n3211) );
  INVX1 U3043 ( .A(n3211), .Y(n3212) );
  AND2X2 U3044 ( .A(\data_in<6> ), .B(n1553), .Y(n3213) );
  INVX1 U3045 ( .A(n3213), .Y(n3214) );
  AND2X2 U3046 ( .A(\data_in<0> ), .B(n1555), .Y(n3215) );
  INVX1 U3047 ( .A(n3215), .Y(n3216) );
  AND2X2 U3048 ( .A(\data_in<1> ), .B(n1555), .Y(n3217) );
  INVX1 U3049 ( .A(n3217), .Y(n3218) );
  AND2X2 U3050 ( .A(\data_in<2> ), .B(n1555), .Y(n3219) );
  INVX1 U3051 ( .A(n3219), .Y(n3220) );
  AND2X2 U3052 ( .A(\data_in<3> ), .B(n1555), .Y(n3221) );
  INVX1 U3053 ( .A(n3221), .Y(n3222) );
  AND2X2 U3054 ( .A(\data_in<4> ), .B(n1555), .Y(n3223) );
  INVX1 U3055 ( .A(n3223), .Y(n3224) );
  AND2X2 U3056 ( .A(\data_in<5> ), .B(n1555), .Y(n3225) );
  INVX1 U3057 ( .A(n3225), .Y(n3226) );
  AND2X2 U3058 ( .A(\data_in<6> ), .B(n1555), .Y(n3227) );
  INVX1 U3059 ( .A(n3227), .Y(n3228) );
  AND2X2 U3060 ( .A(\data_in<7> ), .B(n1555), .Y(n3229) );
  INVX1 U3061 ( .A(n3229), .Y(n3230) );
  AND2X2 U3062 ( .A(\data_in<0> ), .B(n1557), .Y(n3231) );
  INVX1 U3063 ( .A(n3231), .Y(n3232) );
  AND2X2 U3064 ( .A(\data_in<1> ), .B(n1557), .Y(n3233) );
  INVX1 U3065 ( .A(n3233), .Y(n3234) );
  AND2X2 U3066 ( .A(\data_in<2> ), .B(n1557), .Y(n3235) );
  INVX1 U3067 ( .A(n3235), .Y(n3236) );
  AND2X2 U3068 ( .A(\data_in<3> ), .B(n1557), .Y(n3237) );
  INVX1 U3069 ( .A(n3237), .Y(n3238) );
  AND2X2 U3070 ( .A(\data_in<4> ), .B(n1557), .Y(n3239) );
  INVX1 U3071 ( .A(n3239), .Y(n3240) );
  AND2X2 U3072 ( .A(\data_in<5> ), .B(n1557), .Y(n3241) );
  INVX1 U3073 ( .A(n3241), .Y(n3242) );
  AND2X2 U3074 ( .A(\data_in<6> ), .B(n1557), .Y(n3243) );
  INVX1 U3075 ( .A(n3243), .Y(n3244) );
  AND2X2 U3076 ( .A(\data_in<7> ), .B(n1557), .Y(n3245) );
  INVX1 U3077 ( .A(n3245), .Y(n3246) );
  AND2X2 U3078 ( .A(\mem<45><2> ), .B(n5002), .Y(n3247) );
  INVX1 U3079 ( .A(n3247), .Y(n3248) );
  AND2X2 U3080 ( .A(\mem<45><5> ), .B(n5003), .Y(n3249) );
  INVX1 U3081 ( .A(n3249), .Y(n3250) );
  AND2X2 U3082 ( .A(\mem<44><2> ), .B(n5004), .Y(n3251) );
  INVX1 U3083 ( .A(n3251), .Y(n3252) );
  AND2X2 U3084 ( .A(\mem<44><5> ), .B(n5005), .Y(n3253) );
  INVX1 U3085 ( .A(n3253), .Y(n3254) );
  AND2X2 U3086 ( .A(\mem<43><2> ), .B(n5006), .Y(n3255) );
  INVX1 U3087 ( .A(n3255), .Y(n3256) );
  AND2X2 U3088 ( .A(\mem<43><5> ), .B(n5006), .Y(n3257) );
  INVX1 U3089 ( .A(n3257), .Y(n3258) );
  AND2X2 U3090 ( .A(\mem<42><2> ), .B(n5008), .Y(n3259) );
  INVX1 U3091 ( .A(n3259), .Y(n3260) );
  AND2X2 U3092 ( .A(\mem<42><5> ), .B(n5008), .Y(n3261) );
  INVX1 U3093 ( .A(n3261), .Y(n3262) );
  AND2X2 U3094 ( .A(\data_in<0> ), .B(n1576), .Y(n3263) );
  INVX1 U3095 ( .A(n3263), .Y(n3264) );
  AND2X2 U3096 ( .A(\data_in<1> ), .B(n1576), .Y(n3265) );
  INVX1 U3097 ( .A(n3265), .Y(n3266) );
  AND2X2 U3098 ( .A(\data_in<2> ), .B(n1576), .Y(n3267) );
  INVX1 U3099 ( .A(n3267), .Y(n3268) );
  AND2X2 U3100 ( .A(\data_in<3> ), .B(n1576), .Y(n3269) );
  INVX1 U3101 ( .A(n3269), .Y(n3270) );
  AND2X2 U3102 ( .A(\data_in<4> ), .B(n1576), .Y(n3271) );
  INVX1 U3103 ( .A(n3271), .Y(n3272) );
  AND2X2 U3104 ( .A(\data_in<5> ), .B(n1576), .Y(n3273) );
  INVX1 U3105 ( .A(n3273), .Y(n3274) );
  AND2X2 U3106 ( .A(\data_in<6> ), .B(n1576), .Y(n3275) );
  INVX1 U3107 ( .A(n3275), .Y(n3276) );
  AND2X2 U3108 ( .A(\data_in<7> ), .B(n1576), .Y(n3277) );
  INVX1 U3109 ( .A(n3277), .Y(n3278) );
  AND2X2 U3110 ( .A(\data_in<0> ), .B(n1578), .Y(n3279) );
  INVX1 U3111 ( .A(n3279), .Y(n3280) );
  AND2X2 U3112 ( .A(\data_in<1> ), .B(n1578), .Y(n3281) );
  INVX1 U3113 ( .A(n3281), .Y(n3282) );
  AND2X2 U3114 ( .A(\data_in<2> ), .B(n1578), .Y(n3283) );
  INVX1 U3115 ( .A(n3283), .Y(n3284) );
  AND2X2 U3116 ( .A(\data_in<3> ), .B(n1578), .Y(n3285) );
  INVX1 U3117 ( .A(n3285), .Y(n3286) );
  AND2X2 U3118 ( .A(\data_in<4> ), .B(n1578), .Y(n3287) );
  INVX1 U3119 ( .A(n3287), .Y(n3288) );
  AND2X2 U3120 ( .A(\data_in<5> ), .B(n1578), .Y(n3289) );
  INVX1 U3121 ( .A(n3289), .Y(n3290) );
  AND2X2 U3122 ( .A(\data_in<6> ), .B(n1578), .Y(n3291) );
  INVX1 U3123 ( .A(n3291), .Y(n3292) );
  AND2X2 U3124 ( .A(\data_in<7> ), .B(n1578), .Y(n3293) );
  INVX1 U3125 ( .A(n3293), .Y(n3294) );
  AND2X2 U3126 ( .A(\data_in<2> ), .B(n1580), .Y(n3295) );
  INVX1 U3127 ( .A(n3295), .Y(n3296) );
  AND2X2 U3128 ( .A(\data_in<5> ), .B(n1580), .Y(n3297) );
  INVX1 U3129 ( .A(n3297), .Y(n3298) );
  AND2X2 U3130 ( .A(\data_in<0> ), .B(n1586), .Y(n3299) );
  INVX1 U3131 ( .A(n3299), .Y(n3300) );
  AND2X2 U3132 ( .A(\data_in<1> ), .B(n1586), .Y(n3301) );
  INVX1 U3133 ( .A(n3301), .Y(n3302) );
  AND2X2 U3134 ( .A(\data_in<2> ), .B(n1586), .Y(n3303) );
  INVX1 U3135 ( .A(n3303), .Y(n3304) );
  AND2X2 U3136 ( .A(\data_in<3> ), .B(n1586), .Y(n3305) );
  INVX1 U3137 ( .A(n3305), .Y(n3306) );
  AND2X2 U3138 ( .A(\data_in<4> ), .B(n1586), .Y(n3307) );
  INVX1 U3139 ( .A(n3307), .Y(n3308) );
  AND2X2 U3140 ( .A(\data_in<5> ), .B(n1586), .Y(n3309) );
  INVX1 U3141 ( .A(n3309), .Y(n3310) );
  AND2X2 U3142 ( .A(\data_in<6> ), .B(n1586), .Y(n3311) );
  INVX1 U3143 ( .A(n3311), .Y(n3312) );
  AND2X2 U3144 ( .A(\data_in<7> ), .B(n1586), .Y(n3313) );
  INVX1 U3145 ( .A(n3313), .Y(n3314) );
  AND2X2 U3146 ( .A(\data_in<0> ), .B(n1588), .Y(n3315) );
  INVX1 U3147 ( .A(n3315), .Y(n3316) );
  AND2X2 U3148 ( .A(\data_in<1> ), .B(n1588), .Y(n3317) );
  INVX1 U3149 ( .A(n3317), .Y(n3318) );
  AND2X2 U3150 ( .A(\data_in<2> ), .B(n1588), .Y(n3319) );
  INVX1 U3151 ( .A(n3319), .Y(n3320) );
  AND2X2 U3152 ( .A(\data_in<3> ), .B(n1588), .Y(n3321) );
  INVX1 U3153 ( .A(n3321), .Y(n3322) );
  AND2X2 U3154 ( .A(\data_in<4> ), .B(n1588), .Y(n3323) );
  INVX1 U3155 ( .A(n3323), .Y(n3324) );
  AND2X2 U3156 ( .A(\data_in<5> ), .B(n1588), .Y(n3325) );
  INVX1 U3157 ( .A(n3325), .Y(n3326) );
  AND2X2 U3158 ( .A(\data_in<6> ), .B(n1588), .Y(n3327) );
  INVX1 U3159 ( .A(n3327), .Y(n3328) );
  AND2X2 U3160 ( .A(\data_in<0> ), .B(n1590), .Y(n3329) );
  INVX1 U3161 ( .A(n3329), .Y(n3330) );
  AND2X2 U3162 ( .A(\data_in<1> ), .B(n1590), .Y(n3331) );
  INVX1 U3163 ( .A(n3331), .Y(n3332) );
  AND2X2 U3164 ( .A(\data_in<2> ), .B(n1590), .Y(n3333) );
  INVX1 U3165 ( .A(n3333), .Y(n3334) );
  AND2X2 U3166 ( .A(\data_in<3> ), .B(n1590), .Y(n3335) );
  INVX1 U3167 ( .A(n3335), .Y(n3336) );
  AND2X2 U3168 ( .A(\data_in<4> ), .B(n1590), .Y(n3337) );
  INVX1 U3169 ( .A(n3337), .Y(n3338) );
  AND2X2 U3170 ( .A(\data_in<5> ), .B(n1590), .Y(n3339) );
  INVX1 U3171 ( .A(n3339), .Y(n3340) );
  AND2X2 U3172 ( .A(\data_in<6> ), .B(n1590), .Y(n3341) );
  INVX1 U3173 ( .A(n3341), .Y(n3342) );
  AND2X2 U3174 ( .A(\data_in<7> ), .B(n1590), .Y(n3343) );
  INVX1 U3175 ( .A(n3343), .Y(n3344) );
  AND2X2 U3176 ( .A(\data_in<0> ), .B(n1592), .Y(n3345) );
  INVX1 U3177 ( .A(n3345), .Y(n3346) );
  AND2X2 U3178 ( .A(\data_in<1> ), .B(n1592), .Y(n3347) );
  INVX1 U3179 ( .A(n3347), .Y(n3348) );
  AND2X2 U3180 ( .A(\data_in<2> ), .B(n1592), .Y(n3349) );
  INVX1 U3181 ( .A(n3349), .Y(n3350) );
  AND2X2 U3182 ( .A(\data_in<3> ), .B(n1592), .Y(n3351) );
  INVX1 U3183 ( .A(n3351), .Y(n3352) );
  AND2X2 U3184 ( .A(\data_in<4> ), .B(n1592), .Y(n3353) );
  INVX1 U3185 ( .A(n3353), .Y(n3354) );
  AND2X2 U3186 ( .A(\data_in<5> ), .B(n1592), .Y(n3355) );
  INVX1 U3187 ( .A(n3355), .Y(n3356) );
  AND2X2 U3188 ( .A(\data_in<6> ), .B(n1592), .Y(n3357) );
  INVX1 U3189 ( .A(n3357), .Y(n3358) );
  AND2X2 U3190 ( .A(\data_in<7> ), .B(n1592), .Y(n3359) );
  INVX1 U3191 ( .A(n3359), .Y(n3360) );
  AND2X2 U3192 ( .A(\data_in<0> ), .B(n1594), .Y(n3361) );
  INVX1 U3193 ( .A(n3361), .Y(n3362) );
  AND2X2 U3194 ( .A(\data_in<1> ), .B(n1594), .Y(n3363) );
  INVX1 U3195 ( .A(n3363), .Y(n3364) );
  AND2X2 U3196 ( .A(\data_in<2> ), .B(n1594), .Y(n3365) );
  INVX1 U3197 ( .A(n3365), .Y(n3366) );
  AND2X2 U3198 ( .A(\data_in<3> ), .B(n1594), .Y(n3367) );
  INVX1 U3199 ( .A(n3367), .Y(n3368) );
  AND2X2 U3200 ( .A(\data_in<4> ), .B(n1594), .Y(n3369) );
  INVX1 U3201 ( .A(n3369), .Y(n3370) );
  AND2X2 U3202 ( .A(\data_in<5> ), .B(n1594), .Y(n3371) );
  INVX1 U3203 ( .A(n3371), .Y(n3372) );
  AND2X2 U3204 ( .A(\data_in<6> ), .B(n1594), .Y(n3373) );
  INVX1 U3205 ( .A(n3373), .Y(n3374) );
  AND2X2 U3206 ( .A(\data_in<7> ), .B(n1594), .Y(n3375) );
  INVX1 U3207 ( .A(n3375), .Y(n3376) );
  AND2X2 U3208 ( .A(\data_in<0> ), .B(n1596), .Y(n3377) );
  INVX1 U3209 ( .A(n3377), .Y(n3378) );
  AND2X2 U3210 ( .A(\data_in<1> ), .B(n1596), .Y(n3379) );
  INVX1 U3211 ( .A(n3379), .Y(n3380) );
  AND2X2 U3212 ( .A(\data_in<2> ), .B(n1596), .Y(n3381) );
  INVX1 U3213 ( .A(n3381), .Y(n3382) );
  AND2X2 U3214 ( .A(\data_in<3> ), .B(n1596), .Y(n3383) );
  INVX1 U3215 ( .A(n3383), .Y(n3384) );
  AND2X2 U3216 ( .A(\data_in<4> ), .B(n1596), .Y(n3385) );
  INVX1 U3217 ( .A(n3385), .Y(n3386) );
  AND2X2 U3218 ( .A(\data_in<5> ), .B(n1596), .Y(n3387) );
  INVX1 U3219 ( .A(n3387), .Y(n3388) );
  AND2X2 U3220 ( .A(\data_in<6> ), .B(n1596), .Y(n3389) );
  INVX1 U3221 ( .A(n3389), .Y(n3390) );
  AND2X2 U3222 ( .A(\data_in<7> ), .B(n1596), .Y(n3391) );
  INVX1 U3223 ( .A(n3391), .Y(n3392) );
  AND2X2 U3224 ( .A(\data_in<0> ), .B(n1598), .Y(n3393) );
  INVX1 U3225 ( .A(n3393), .Y(n3394) );
  AND2X2 U3226 ( .A(\data_in<1> ), .B(n1598), .Y(n3395) );
  INVX1 U3227 ( .A(n3395), .Y(n3396) );
  AND2X2 U3228 ( .A(\data_in<2> ), .B(n1598), .Y(n3397) );
  INVX1 U3229 ( .A(n3397), .Y(n3398) );
  AND2X2 U3230 ( .A(\data_in<3> ), .B(n1598), .Y(n3399) );
  INVX1 U3231 ( .A(n3399), .Y(n3400) );
  AND2X2 U3232 ( .A(\data_in<4> ), .B(n1598), .Y(n3401) );
  INVX1 U3233 ( .A(n3401), .Y(n3402) );
  AND2X2 U3234 ( .A(\data_in<5> ), .B(n1598), .Y(n3403) );
  INVX1 U3235 ( .A(n3403), .Y(n3404) );
  AND2X2 U3236 ( .A(\data_in<6> ), .B(n1598), .Y(n3405) );
  INVX1 U3237 ( .A(n3405), .Y(n3406) );
  AND2X2 U3238 ( .A(\data_in<7> ), .B(n1598), .Y(n3407) );
  INVX1 U3239 ( .A(n3407), .Y(n3408) );
  AND2X2 U3240 ( .A(\data_in<0> ), .B(n1600), .Y(n3409) );
  INVX1 U3241 ( .A(n3409), .Y(n3410) );
  AND2X2 U3242 ( .A(\data_in<1> ), .B(n1600), .Y(n3411) );
  INVX1 U3243 ( .A(n3411), .Y(n3412) );
  AND2X2 U3244 ( .A(\data_in<2> ), .B(n1600), .Y(n3413) );
  INVX1 U3245 ( .A(n3413), .Y(n3414) );
  AND2X2 U3246 ( .A(\data_in<3> ), .B(n1600), .Y(n3415) );
  INVX1 U3247 ( .A(n3415), .Y(n3416) );
  AND2X2 U3248 ( .A(\data_in<4> ), .B(n1600), .Y(n3417) );
  INVX1 U3249 ( .A(n3417), .Y(n3418) );
  AND2X2 U3250 ( .A(\data_in<5> ), .B(n1600), .Y(n3419) );
  INVX1 U3251 ( .A(n3419), .Y(n3420) );
  AND2X2 U3252 ( .A(\data_in<6> ), .B(n1600), .Y(n3421) );
  INVX1 U3253 ( .A(n3421), .Y(n3422) );
  AND2X2 U3254 ( .A(\data_in<7> ), .B(n1600), .Y(n3423) );
  INVX1 U3255 ( .A(n3423), .Y(n3424) );
  AND2X2 U3256 ( .A(\data_in<0> ), .B(n1602), .Y(n3425) );
  INVX1 U3257 ( .A(n3425), .Y(n3426) );
  AND2X2 U3258 ( .A(\data_in<1> ), .B(n1602), .Y(n3427) );
  INVX1 U3259 ( .A(n3427), .Y(n3428) );
  AND2X2 U3260 ( .A(\data_in<2> ), .B(n1602), .Y(n3429) );
  INVX1 U3261 ( .A(n3429), .Y(n3430) );
  AND2X2 U3262 ( .A(\data_in<3> ), .B(n1602), .Y(n3431) );
  INVX1 U3263 ( .A(n3431), .Y(n3432) );
  AND2X2 U3264 ( .A(\data_in<4> ), .B(n1602), .Y(n3433) );
  INVX1 U3265 ( .A(n3433), .Y(n3434) );
  AND2X2 U3266 ( .A(\data_in<5> ), .B(n1602), .Y(n3435) );
  INVX1 U3267 ( .A(n3435), .Y(n3436) );
  AND2X2 U3268 ( .A(\data_in<6> ), .B(n1602), .Y(n3437) );
  INVX1 U3269 ( .A(n3437), .Y(n3438) );
  AND2X2 U3270 ( .A(\data_in<7> ), .B(n1602), .Y(n3439) );
  INVX1 U3271 ( .A(n3439), .Y(n3440) );
  AND2X2 U3272 ( .A(\data_in<0> ), .B(n1604), .Y(n3441) );
  INVX1 U3273 ( .A(n3441), .Y(n3442) );
  AND2X2 U3274 ( .A(\data_in<1> ), .B(n1604), .Y(n3443) );
  INVX1 U3275 ( .A(n3443), .Y(n3444) );
  AND2X2 U3276 ( .A(\data_in<2> ), .B(n1604), .Y(n3445) );
  INVX1 U3277 ( .A(n3445), .Y(n3446) );
  AND2X2 U3278 ( .A(\data_in<3> ), .B(n1604), .Y(n3447) );
  INVX1 U3279 ( .A(n3447), .Y(n3448) );
  AND2X2 U3280 ( .A(\data_in<4> ), .B(n1604), .Y(n3449) );
  INVX1 U3281 ( .A(n3449), .Y(n3450) );
  AND2X2 U3282 ( .A(\data_in<5> ), .B(n1604), .Y(n3451) );
  INVX1 U3283 ( .A(n3451), .Y(n3452) );
  AND2X2 U3284 ( .A(\data_in<6> ), .B(n1604), .Y(n3453) );
  INVX1 U3285 ( .A(n3453), .Y(n3454) );
  AND2X2 U3286 ( .A(\data_in<7> ), .B(n1604), .Y(n3455) );
  INVX1 U3287 ( .A(n3455), .Y(n3456) );
  AND2X2 U3288 ( .A(\data_in<0> ), .B(n1606), .Y(n3457) );
  INVX1 U3289 ( .A(n3457), .Y(n3458) );
  AND2X2 U3290 ( .A(\data_in<1> ), .B(n1606), .Y(n3459) );
  INVX1 U3291 ( .A(n3459), .Y(n3460) );
  AND2X2 U3292 ( .A(\data_in<2> ), .B(n1606), .Y(n3461) );
  INVX1 U3293 ( .A(n3461), .Y(n3462) );
  AND2X2 U3294 ( .A(\data_in<3> ), .B(n1606), .Y(n3463) );
  INVX1 U3295 ( .A(n3463), .Y(n3464) );
  AND2X2 U3296 ( .A(\data_in<4> ), .B(n1606), .Y(n3465) );
  INVX1 U3297 ( .A(n3465), .Y(n3466) );
  AND2X2 U3298 ( .A(\data_in<5> ), .B(n1606), .Y(n3467) );
  INVX1 U3299 ( .A(n3467), .Y(n3468) );
  AND2X2 U3300 ( .A(\data_in<6> ), .B(n1606), .Y(n3469) );
  INVX1 U3301 ( .A(n3469), .Y(n3470) );
  AND2X2 U3302 ( .A(\data_in<7> ), .B(n1606), .Y(n3471) );
  INVX1 U3303 ( .A(n3471), .Y(n3472) );
  AND2X2 U3304 ( .A(\data_in<0> ), .B(n1608), .Y(n3473) );
  INVX1 U3305 ( .A(n3473), .Y(n3474) );
  AND2X2 U3306 ( .A(\data_in<1> ), .B(n1608), .Y(n3475) );
  INVX1 U3307 ( .A(n3475), .Y(n3476) );
  AND2X2 U3308 ( .A(\data_in<2> ), .B(n1608), .Y(n3477) );
  INVX1 U3309 ( .A(n3477), .Y(n3478) );
  AND2X2 U3310 ( .A(\data_in<3> ), .B(n1608), .Y(n3479) );
  INVX1 U3311 ( .A(n3479), .Y(n3480) );
  AND2X2 U3312 ( .A(\data_in<4> ), .B(n1608), .Y(n3481) );
  INVX1 U3313 ( .A(n3481), .Y(n3482) );
  AND2X2 U3314 ( .A(\data_in<5> ), .B(n1608), .Y(n3483) );
  INVX1 U3315 ( .A(n3483), .Y(n3484) );
  AND2X2 U3316 ( .A(\data_in<6> ), .B(n1608), .Y(n3485) );
  INVX1 U3317 ( .A(n3485), .Y(n3486) );
  AND2X2 U3318 ( .A(\data_in<7> ), .B(n1608), .Y(n3487) );
  INVX1 U3319 ( .A(n3487), .Y(n3488) );
  AND2X2 U3320 ( .A(\data_in<0> ), .B(n1610), .Y(n3489) );
  INVX1 U3321 ( .A(n3489), .Y(n3490) );
  AND2X2 U3322 ( .A(\data_in<1> ), .B(n1610), .Y(n3491) );
  INVX1 U3323 ( .A(n3491), .Y(n3492) );
  AND2X2 U3324 ( .A(\data_in<2> ), .B(n1610), .Y(n3493) );
  INVX1 U3325 ( .A(n3493), .Y(n3494) );
  AND2X2 U3326 ( .A(\data_in<3> ), .B(n1610), .Y(n3495) );
  INVX1 U3327 ( .A(n3495), .Y(n3496) );
  AND2X2 U3328 ( .A(\data_in<4> ), .B(n1610), .Y(n3497) );
  INVX1 U3329 ( .A(n3497), .Y(n3498) );
  AND2X2 U3330 ( .A(\data_in<5> ), .B(n1610), .Y(n3499) );
  INVX1 U3331 ( .A(n3499), .Y(n3500) );
  AND2X2 U3332 ( .A(\data_in<6> ), .B(n1610), .Y(n3501) );
  INVX1 U3333 ( .A(n3501), .Y(n3502) );
  AND2X2 U3334 ( .A(\data_in<7> ), .B(n1610), .Y(n3503) );
  INVX1 U3335 ( .A(n3503), .Y(n3504) );
  AND2X2 U3336 ( .A(\data_in<0> ), .B(n1614), .Y(n3505) );
  INVX1 U3337 ( .A(n3505), .Y(n3506) );
  AND2X2 U3338 ( .A(\data_in<1> ), .B(n1614), .Y(n3507) );
  INVX1 U3339 ( .A(n3507), .Y(n3508) );
  AND2X2 U3340 ( .A(\data_in<2> ), .B(n1614), .Y(n3509) );
  INVX1 U3341 ( .A(n3509), .Y(n3510) );
  AND2X2 U3342 ( .A(\data_in<3> ), .B(n1614), .Y(n3511) );
  INVX1 U3343 ( .A(n3511), .Y(n3512) );
  AND2X2 U3344 ( .A(\data_in<4> ), .B(n1614), .Y(n3513) );
  INVX1 U3345 ( .A(n3513), .Y(n3514) );
  AND2X2 U3346 ( .A(\data_in<5> ), .B(n1614), .Y(n3515) );
  INVX1 U3347 ( .A(n3515), .Y(n3516) );
  AND2X2 U3348 ( .A(\data_in<6> ), .B(n1614), .Y(n3517) );
  INVX1 U3349 ( .A(n3517), .Y(n3518) );
  AND2X2 U3350 ( .A(\data_in<7> ), .B(n1614), .Y(n3519) );
  INVX1 U3351 ( .A(n3519), .Y(n3520) );
  AND2X2 U3352 ( .A(\data_in<0> ), .B(n1616), .Y(n3521) );
  INVX1 U3353 ( .A(n3521), .Y(n3522) );
  AND2X2 U3354 ( .A(\data_in<1> ), .B(n1616), .Y(n3523) );
  INVX1 U3355 ( .A(n3523), .Y(n3524) );
  AND2X2 U3356 ( .A(\data_in<2> ), .B(n1616), .Y(n3525) );
  INVX1 U3357 ( .A(n3525), .Y(n3526) );
  AND2X2 U3358 ( .A(\data_in<3> ), .B(n1616), .Y(n3527) );
  INVX1 U3359 ( .A(n3527), .Y(n3528) );
  AND2X2 U3360 ( .A(\data_in<4> ), .B(n1616), .Y(n3529) );
  INVX1 U3361 ( .A(n3529), .Y(n3530) );
  AND2X2 U3362 ( .A(\data_in<5> ), .B(n1616), .Y(n3531) );
  INVX1 U3363 ( .A(n3531), .Y(n3532) );
  AND2X2 U3364 ( .A(\data_in<6> ), .B(n1616), .Y(n3533) );
  INVX1 U3365 ( .A(n3533), .Y(n3534) );
  AND2X2 U3366 ( .A(\data_in<7> ), .B(n1616), .Y(n3535) );
  INVX1 U3367 ( .A(n3535), .Y(n3536) );
  AND2X2 U3368 ( .A(\data_in<0> ), .B(n1618), .Y(n3537) );
  INVX1 U3369 ( .A(n3537), .Y(n3538) );
  AND2X2 U3370 ( .A(\data_in<1> ), .B(n1618), .Y(n3539) );
  INVX1 U3371 ( .A(n3539), .Y(n3540) );
  AND2X2 U3372 ( .A(\data_in<2> ), .B(n1618), .Y(n3541) );
  INVX1 U3373 ( .A(n3541), .Y(n3542) );
  AND2X2 U3374 ( .A(\data_in<3> ), .B(n1618), .Y(n3543) );
  INVX1 U3375 ( .A(n3543), .Y(n3544) );
  AND2X2 U3376 ( .A(\data_in<4> ), .B(n1618), .Y(n3545) );
  INVX1 U3377 ( .A(n3545), .Y(n3546) );
  AND2X2 U3378 ( .A(\data_in<5> ), .B(n1618), .Y(n3547) );
  INVX1 U3379 ( .A(n3547), .Y(n3548) );
  AND2X2 U3380 ( .A(\data_in<6> ), .B(n1618), .Y(n3549) );
  INVX1 U3381 ( .A(n3549), .Y(n3550) );
  AND2X2 U3382 ( .A(\data_in<7> ), .B(n1618), .Y(n3551) );
  INVX1 U3383 ( .A(n3551), .Y(n3552) );
  AND2X2 U3384 ( .A(\data_in<0> ), .B(n1623), .Y(n3553) );
  INVX1 U3385 ( .A(n3553), .Y(n3554) );
  AND2X2 U3386 ( .A(\data_in<1> ), .B(n1623), .Y(n3555) );
  INVX1 U3387 ( .A(n3555), .Y(n3556) );
  AND2X2 U3388 ( .A(\data_in<2> ), .B(n1623), .Y(n3557) );
  INVX1 U3389 ( .A(n3557), .Y(n3558) );
  AND2X2 U3390 ( .A(\data_in<3> ), .B(n1623), .Y(n3559) );
  INVX1 U3391 ( .A(n3559), .Y(n3560) );
  AND2X2 U3392 ( .A(\data_in<4> ), .B(n1623), .Y(n3561) );
  INVX1 U3393 ( .A(n3561), .Y(n3562) );
  AND2X2 U3394 ( .A(\data_in<5> ), .B(n1623), .Y(n3563) );
  INVX1 U3395 ( .A(n3563), .Y(n3564) );
  AND2X2 U3396 ( .A(\data_in<6> ), .B(n1623), .Y(n3565) );
  INVX1 U3397 ( .A(n3565), .Y(n3566) );
  AND2X2 U3398 ( .A(\data_in<7> ), .B(n1623), .Y(n3567) );
  INVX1 U3399 ( .A(n3567), .Y(n3568) );
  AND2X2 U3400 ( .A(\data_in<0> ), .B(n1625), .Y(n3569) );
  INVX1 U3401 ( .A(n3569), .Y(n3570) );
  AND2X2 U3402 ( .A(\data_in<1> ), .B(n1625), .Y(n3571) );
  INVX1 U3403 ( .A(n3571), .Y(n3572) );
  AND2X2 U3404 ( .A(\data_in<2> ), .B(n1625), .Y(n3573) );
  INVX1 U3405 ( .A(n3573), .Y(n3574) );
  AND2X2 U3406 ( .A(\data_in<3> ), .B(n1625), .Y(n3575) );
  INVX1 U3407 ( .A(n3575), .Y(n3576) );
  AND2X2 U3408 ( .A(\data_in<4> ), .B(n1625), .Y(n3577) );
  INVX1 U3409 ( .A(n3577), .Y(n3578) );
  AND2X2 U3410 ( .A(\data_in<5> ), .B(n1625), .Y(n3579) );
  INVX1 U3411 ( .A(n3579), .Y(n3580) );
  AND2X2 U3412 ( .A(\data_in<6> ), .B(n1625), .Y(n3581) );
  INVX1 U3413 ( .A(n3581), .Y(n3582) );
  AND2X2 U3414 ( .A(\data_in<7> ), .B(n1625), .Y(n3583) );
  INVX1 U3415 ( .A(n3583), .Y(n3584) );
  AND2X2 U3416 ( .A(\data_in<0> ), .B(n1626), .Y(n3585) );
  INVX1 U3417 ( .A(n3585), .Y(n3586) );
  AND2X2 U3418 ( .A(\data_in<1> ), .B(n1626), .Y(n3587) );
  INVX1 U3419 ( .A(n3587), .Y(n3588) );
  AND2X2 U3420 ( .A(\data_in<2> ), .B(n1626), .Y(n3589) );
  INVX1 U3421 ( .A(n3589), .Y(n3590) );
  AND2X2 U3422 ( .A(\data_in<3> ), .B(n1626), .Y(n3591) );
  INVX1 U3423 ( .A(n3591), .Y(n3592) );
  AND2X2 U3424 ( .A(\data_in<4> ), .B(n1626), .Y(n3593) );
  INVX1 U3425 ( .A(n3593), .Y(n3594) );
  AND2X2 U3426 ( .A(\data_in<5> ), .B(n1626), .Y(n3595) );
  INVX1 U3427 ( .A(n3595), .Y(n3596) );
  AND2X2 U3428 ( .A(\data_in<6> ), .B(n1626), .Y(n3597) );
  INVX1 U3429 ( .A(n3597), .Y(n3598) );
  AND2X2 U3430 ( .A(\data_in<7> ), .B(n1626), .Y(n3599) );
  INVX1 U3431 ( .A(n3599), .Y(n3600) );
  AND2X2 U3432 ( .A(\data_in<0> ), .B(n1628), .Y(n3601) );
  INVX1 U3433 ( .A(n3601), .Y(n3602) );
  AND2X2 U3434 ( .A(\data_in<1> ), .B(n1628), .Y(n3603) );
  INVX1 U3435 ( .A(n3603), .Y(n3604) );
  AND2X2 U3436 ( .A(\data_in<2> ), .B(n1628), .Y(n3605) );
  INVX1 U3437 ( .A(n3605), .Y(n3606) );
  AND2X2 U3438 ( .A(\data_in<3> ), .B(n1628), .Y(n3607) );
  INVX1 U3439 ( .A(n3607), .Y(n3608) );
  AND2X2 U3440 ( .A(\data_in<4> ), .B(n1628), .Y(n3609) );
  INVX1 U3441 ( .A(n3609), .Y(n3610) );
  AND2X2 U3442 ( .A(\data_in<5> ), .B(n1628), .Y(n3611) );
  INVX1 U3443 ( .A(n3611), .Y(n3612) );
  AND2X2 U3444 ( .A(\data_in<6> ), .B(n1628), .Y(n3613) );
  INVX1 U3445 ( .A(n3613), .Y(n3614) );
  AND2X2 U3446 ( .A(\data_in<7> ), .B(n1628), .Y(n3615) );
  INVX1 U3447 ( .A(n3615), .Y(n3616) );
  AND2X2 U3448 ( .A(\mem<10><3> ), .B(n5060), .Y(n3617) );
  INVX1 U3449 ( .A(n3617), .Y(n3618) );
  AND2X2 U3450 ( .A(\mem<10><7> ), .B(n5060), .Y(n3619) );
  INVX1 U3451 ( .A(n3619), .Y(n3620) );
  AND2X2 U3452 ( .A(\data_in<0> ), .B(n1632), .Y(n3621) );
  INVX1 U3453 ( .A(n3621), .Y(n3622) );
  AND2X2 U3454 ( .A(\data_in<1> ), .B(n1632), .Y(n3623) );
  INVX1 U3455 ( .A(n3623), .Y(n3624) );
  AND2X2 U3456 ( .A(\data_in<2> ), .B(n1632), .Y(n3625) );
  INVX1 U3457 ( .A(n3625), .Y(n3626) );
  AND2X2 U3458 ( .A(\data_in<3> ), .B(n1632), .Y(n3627) );
  INVX1 U3459 ( .A(n3627), .Y(n3628) );
  AND2X2 U3460 ( .A(\data_in<4> ), .B(n1632), .Y(n3629) );
  INVX1 U3461 ( .A(n3629), .Y(n3630) );
  AND2X2 U3462 ( .A(\data_in<5> ), .B(n1632), .Y(n3631) );
  INVX1 U3463 ( .A(n3631), .Y(n3632) );
  AND2X2 U3464 ( .A(\data_in<6> ), .B(n1632), .Y(n3633) );
  INVX1 U3465 ( .A(n3633), .Y(n3634) );
  AND2X2 U3466 ( .A(\data_in<7> ), .B(n1632), .Y(n3635) );
  INVX1 U3467 ( .A(n3635), .Y(n3636) );
  AND2X2 U3468 ( .A(\mem<5><2> ), .B(n5065), .Y(n3637) );
  INVX1 U3469 ( .A(n3637), .Y(n3638) );
  AND2X2 U3470 ( .A(\mem<5><5> ), .B(n5066), .Y(n3639) );
  INVX1 U3471 ( .A(n3639), .Y(n3640) );
  AND2X2 U3472 ( .A(\data_in<2> ), .B(n1641), .Y(n3641) );
  INVX1 U3473 ( .A(n3641), .Y(n3642) );
  AND2X2 U3474 ( .A(\data_in<5> ), .B(n1641), .Y(n3643) );
  INVX1 U3475 ( .A(n3643), .Y(n3644) );
  AND2X2 U3476 ( .A(\data_in<6> ), .B(n1643), .Y(n3645) );
  INVX1 U3477 ( .A(n3645), .Y(n3646) );
  AND2X2 U3478 ( .A(\data_in<7> ), .B(n1643), .Y(n3647) );
  INVX1 U3479 ( .A(n3647), .Y(n3648) );
  AND2X2 U3480 ( .A(\data_in<2> ), .B(n1645), .Y(n3649) );
  INVX1 U3481 ( .A(n3649), .Y(n3650) );
  AND2X2 U3482 ( .A(\data_in<5> ), .B(n1645), .Y(n3651) );
  INVX1 U3483 ( .A(n3651), .Y(n3652) );
  OR2X2 U3484 ( .A(n5153), .B(n5766), .Y(n3653) );
  INVX1 U3485 ( .A(n3653), .Y(n3654) );
  INVX1 U3486 ( .A(n3653), .Y(n3655) );
  OR2X2 U3487 ( .A(n5080), .B(n634), .Y(n3656) );
  OR2X2 U3488 ( .A(n5113), .B(n5761), .Y(n3658) );
  OR2X2 U3489 ( .A(n4171), .B(\addr<15> ), .Y(n3661) );
  INVX1 U3490 ( .A(n3661), .Y(n3662) );
  OR2X2 U3491 ( .A(n5184), .B(n4172), .Y(n3663) );
  INVX1 U3492 ( .A(n3663), .Y(n3664) );
  AND2X2 U3493 ( .A(n5726), .B(n5700), .Y(n3665) );
  INVX1 U3494 ( .A(n3665), .Y(n3666) );
  INVX1 U3495 ( .A(n3665), .Y(n3667) );
  AND2X2 U3496 ( .A(n212), .B(n5726), .Y(n3668) );
  INVX1 U3497 ( .A(n3668), .Y(n3669) );
  INVX1 U3498 ( .A(n3668), .Y(n3670) );
  AND2X2 U3499 ( .A(n5726), .B(n5708), .Y(n3671) );
  INVX1 U3500 ( .A(n3671), .Y(n3672) );
  INVX1 U3501 ( .A(n3671), .Y(n3673) );
  OR2X2 U3502 ( .A(n3926), .B(n4943), .Y(n3674) );
  INVX1 U3503 ( .A(n3674), .Y(n3675) );
  AND2X2 U3504 ( .A(n5726), .B(n409), .Y(n3676) );
  INVX1 U3505 ( .A(n3676), .Y(n3677) );
  INVX1 U3506 ( .A(n3676), .Y(n3678) );
  AND2X2 U3507 ( .A(n5725), .B(n5181), .Y(n3679) );
  INVX1 U3508 ( .A(n3679), .Y(n3680) );
  INVX1 U3509 ( .A(n3679), .Y(n3681) );
  BUFX2 U3510 ( .A(n6458), .Y(n5716) );
  OR2X2 U3511 ( .A(\addr<15> ), .B(n1137), .Y(n3682) );
  INVX1 U3512 ( .A(n3682), .Y(n3683) );
  OR2X2 U3513 ( .A(n3764), .B(n3964), .Y(n3684) );
  INVX1 U3514 ( .A(n3684), .Y(n3685) );
  AND2X2 U3515 ( .A(enable), .B(n5856), .Y(n3686) );
  AND2X2 U3516 ( .A(n5516), .B(n5654), .Y(n3687) );
  INVX1 U3517 ( .A(n3687), .Y(n3688) );
  AND2X2 U3518 ( .A(n5366), .B(n5185), .Y(n3689) );
  INVX1 U3519 ( .A(n3689), .Y(n3690) );
  AND2X2 U3520 ( .A(n5374), .B(n5656), .Y(n3691) );
  INVX1 U3521 ( .A(n3691), .Y(n3692) );
  AND2X2 U3522 ( .A(n5278), .B(n3919), .Y(n3693) );
  INVX1 U3523 ( .A(n3693), .Y(n3694) );
  AND2X2 U3524 ( .A(n5467), .B(n3948), .Y(n3695) );
  INVX1 U3525 ( .A(n3695), .Y(n3696) );
  AND2X2 U3526 ( .A(n5474), .B(n5654), .Y(n3697) );
  INVX1 U3527 ( .A(n3697), .Y(n3698) );
  AND2X2 U3528 ( .A(n5326), .B(n5656), .Y(n3699) );
  INVX1 U3529 ( .A(n3699), .Y(n3700) );
  AND2X2 U3530 ( .A(n5469), .B(n5654), .Y(n3701) );
  INVX1 U3531 ( .A(n3701), .Y(n3702) );
  AND2X2 U3532 ( .A(n5461), .B(n5654), .Y(n3703) );
  INVX1 U3533 ( .A(n3703), .Y(n3704) );
  AND2X2 U3534 ( .A(n5453), .B(n5084), .Y(n3705) );
  INVX1 U3535 ( .A(n3705), .Y(n3706) );
  AND2X2 U3536 ( .A(n5384), .B(n5655), .Y(n3707) );
  INVX1 U3537 ( .A(n3707), .Y(n3708) );
  AND2X2 U3538 ( .A(n5390), .B(n5217), .Y(n3709) );
  INVX1 U3539 ( .A(n3709), .Y(n3710) );
  AND2X2 U3540 ( .A(n5243), .B(n5191), .Y(n3711) );
  INVX1 U3541 ( .A(n3711), .Y(n3712) );
  AND2X2 U3542 ( .A(n5343), .B(n5204), .Y(n3713) );
  INVX1 U3543 ( .A(n3713), .Y(n3714) );
  AND2X2 U3544 ( .A(n5383), .B(n5217), .Y(n3715) );
  INVX1 U3545 ( .A(n3715), .Y(n3716) );
  AND2X2 U3546 ( .A(n5553), .B(n5653), .Y(n3717) );
  INVX1 U3547 ( .A(n3717), .Y(n3718) );
  OR2X2 U3548 ( .A(n6162), .B(n6161), .Y(n3719) );
  INVX1 U3549 ( .A(n3719), .Y(n3720) );
  AND2X2 U3550 ( .A(n5519), .B(n3956), .Y(n3721) );
  INVX1 U3551 ( .A(n3721), .Y(n3722) );
  INVX1 U3552 ( .A(n3723), .Y(n3724) );
  AND2X2 U3553 ( .A(n5376), .B(n5206), .Y(n3725) );
  INVX1 U3554 ( .A(n3725), .Y(n3726) );
  AND2X2 U3555 ( .A(n5275), .B(n3918), .Y(n3727) );
  INVX1 U3556 ( .A(n3727), .Y(n3728) );
  AND2X2 U3557 ( .A(n5479), .B(n5084), .Y(n3729) );
  INVX1 U3558 ( .A(n3729), .Y(n3730) );
  AND2X2 U3559 ( .A(n5476), .B(n3949), .Y(n3731) );
  INVX1 U3560 ( .A(n3731), .Y(n3732) );
  AND2X2 U3561 ( .A(n5329), .B(n3996), .Y(n3733) );
  INVX1 U3562 ( .A(n3733), .Y(n3734) );
  AND2X2 U3563 ( .A(n5472), .B(n5209), .Y(n3735) );
  INVX1 U3564 ( .A(n3735), .Y(n3736) );
  AND2X2 U3565 ( .A(n5464), .B(n5173), .Y(n3737) );
  INVX1 U3566 ( .A(n3737), .Y(n3738) );
  INVX1 U3567 ( .A(n3739), .Y(n3740) );
  AND2X2 U3568 ( .A(n5618), .B(n3955), .Y(n3741) );
  INVX1 U3569 ( .A(n3741), .Y(n3742) );
  AND2X2 U3570 ( .A(n5386), .B(n5208), .Y(n3743) );
  INVX1 U3571 ( .A(n3743), .Y(n3744) );
  AND2X2 U3572 ( .A(n5240), .B(n3973), .Y(n3745) );
  INVX1 U3573 ( .A(n3745), .Y(n3746) );
  AND2X2 U3574 ( .A(n5352), .B(n3984), .Y(n3747) );
  INVX1 U3575 ( .A(n3747), .Y(n3748) );
  AND2X2 U3576 ( .A(n5340), .B(n3985), .Y(n3749) );
  INVX1 U3577 ( .A(n3749), .Y(n3750) );
  AND2X2 U3578 ( .A(n5324), .B(n5086), .Y(n3751) );
  INVX1 U3579 ( .A(n3751), .Y(n3752) );
  AND2X2 U3580 ( .A(n5304), .B(n5209), .Y(n3753) );
  INVX1 U3581 ( .A(n3753), .Y(n3754) );
  AND2X2 U3582 ( .A(n5381), .B(n5655), .Y(n3755) );
  INVX1 U3583 ( .A(n3755), .Y(n3756) );
  AND2X2 U3584 ( .A(n5556), .B(n3996), .Y(n3757) );
  INVX1 U3585 ( .A(n3757), .Y(n3758) );
  AND2X2 U3586 ( .A(n5321), .B(n5209), .Y(n3759) );
  INVX1 U3587 ( .A(n3759), .Y(n3760) );
  OR2X2 U3588 ( .A(n5999), .B(n5998), .Y(n3761) );
  INVX1 U3589 ( .A(n3761), .Y(n3762) );
  AND2X2 U3590 ( .A(N178), .B(n5757), .Y(n3763) );
  INVX1 U3591 ( .A(n3763), .Y(n3764) );
  AND2X2 U3592 ( .A(n919), .B(n76), .Y(n3765) );
  INVX1 U3593 ( .A(n3765), .Y(n3766) );
  AND2X2 U3594 ( .A(\mem<48><0> ), .B(n6402), .Y(n3767) );
  INVX1 U3595 ( .A(n3767), .Y(n3768) );
  AND2X2 U3596 ( .A(\mem<48><1> ), .B(n6402), .Y(n3769) );
  INVX1 U3597 ( .A(n3769), .Y(n3770) );
  AND2X2 U3598 ( .A(\mem<48><2> ), .B(n6402), .Y(n3771) );
  INVX1 U3599 ( .A(n3771), .Y(n3772) );
  AND2X2 U3600 ( .A(\data_in<3> ), .B(n3914), .Y(n3773) );
  INVX1 U3601 ( .A(n3773), .Y(n3774) );
  AND2X2 U3602 ( .A(n108), .B(\data_in<4> ), .Y(n3775) );
  INVX1 U3603 ( .A(n3775), .Y(n3776) );
  AND2X2 U3604 ( .A(n108), .B(\data_in<5> ), .Y(n3777) );
  INVX1 U3605 ( .A(n3777), .Y(n3778) );
  AND2X2 U3606 ( .A(n3915), .B(\data_in<6> ), .Y(n3779) );
  INVX1 U3607 ( .A(n3779), .Y(n3780) );
  AND2X2 U3608 ( .A(n3915), .B(\data_in<7> ), .Y(n3781) );
  INVX1 U3609 ( .A(n3781), .Y(n3782) );
  AND2X2 U3610 ( .A(\data_in<0> ), .B(n1574), .Y(n3783) );
  INVX1 U3611 ( .A(n3783), .Y(n3784) );
  AND2X2 U3612 ( .A(\data_in<1> ), .B(n1574), .Y(n3785) );
  INVX1 U3613 ( .A(n3785), .Y(n3786) );
  AND2X2 U3614 ( .A(\data_in<2> ), .B(n1574), .Y(n3787) );
  INVX1 U3615 ( .A(n3787), .Y(n3788) );
  AND2X2 U3616 ( .A(\data_in<3> ), .B(n1574), .Y(n3789) );
  INVX1 U3617 ( .A(n3789), .Y(n3790) );
  AND2X2 U3618 ( .A(\data_in<4> ), .B(n1574), .Y(n3791) );
  INVX1 U3619 ( .A(n3791), .Y(n3792) );
  AND2X2 U3620 ( .A(\data_in<5> ), .B(n1574), .Y(n3793) );
  INVX1 U3621 ( .A(n3793), .Y(n3794) );
  AND2X2 U3622 ( .A(\data_in<6> ), .B(n1574), .Y(n3795) );
  INVX1 U3623 ( .A(n3795), .Y(n3796) );
  AND2X2 U3624 ( .A(\data_in<7> ), .B(n1574), .Y(n3797) );
  INVX1 U3625 ( .A(n3797), .Y(n3798) );
  AND2X2 U3626 ( .A(\data_in<0> ), .B(n1620), .Y(n3799) );
  INVX1 U3627 ( .A(n3799), .Y(n3800) );
  AND2X2 U3628 ( .A(\data_in<1> ), .B(n1620), .Y(n3801) );
  INVX1 U3629 ( .A(n3801), .Y(n3802) );
  AND2X2 U3630 ( .A(\data_in<2> ), .B(n1620), .Y(n3803) );
  INVX1 U3631 ( .A(n3803), .Y(n3804) );
  AND2X2 U3632 ( .A(\data_in<3> ), .B(n1620), .Y(n3805) );
  INVX1 U3633 ( .A(n3805), .Y(n3806) );
  AND2X2 U3634 ( .A(\data_in<4> ), .B(n1620), .Y(n3807) );
  INVX1 U3635 ( .A(n3807), .Y(n3808) );
  AND2X2 U3636 ( .A(\data_in<5> ), .B(n1620), .Y(n3809) );
  INVX1 U3637 ( .A(n3809), .Y(n3810) );
  AND2X2 U3638 ( .A(\data_in<6> ), .B(n1620), .Y(n3811) );
  INVX1 U3639 ( .A(n3811), .Y(n3812) );
  AND2X2 U3640 ( .A(\data_in<7> ), .B(n1620), .Y(n3813) );
  INVX1 U3641 ( .A(n3813), .Y(n3814) );
  AND2X2 U3642 ( .A(\mem<13><0> ), .B(n5055), .Y(n3815) );
  INVX1 U3643 ( .A(n3815), .Y(n3816) );
  AND2X2 U3644 ( .A(\mem<13><1> ), .B(n5056), .Y(n3817) );
  INVX1 U3645 ( .A(n3817), .Y(n3818) );
  AND2X2 U3646 ( .A(\mem<13><2> ), .B(n5055), .Y(n3819) );
  INVX1 U3647 ( .A(n3819), .Y(n3820) );
  AND2X2 U3648 ( .A(\mem<13><3> ), .B(n5056), .Y(n3821) );
  INVX1 U3649 ( .A(n3821), .Y(n3822) );
  AND2X2 U3650 ( .A(\mem<13><4> ), .B(n5055), .Y(n3823) );
  INVX1 U3651 ( .A(n3823), .Y(n3824) );
  AND2X2 U3652 ( .A(\mem<13><5> ), .B(n5056), .Y(n3825) );
  INVX1 U3653 ( .A(n3825), .Y(n3826) );
  AND2X2 U3654 ( .A(\mem<13><6> ), .B(n5055), .Y(n3827) );
  INVX1 U3655 ( .A(n3827), .Y(n3828) );
  AND2X2 U3656 ( .A(\mem<13><7> ), .B(n5056), .Y(n3829) );
  INVX1 U3657 ( .A(n3829), .Y(n3830) );
  AND2X2 U3658 ( .A(\mem<9><0> ), .B(n5061), .Y(n3831) );
  INVX1 U3659 ( .A(n3831), .Y(n3832) );
  AND2X2 U3660 ( .A(\mem<9><1> ), .B(n5062), .Y(n3833) );
  INVX1 U3661 ( .A(n3833), .Y(n3834) );
  AND2X2 U3662 ( .A(\mem<9><3> ), .B(n5062), .Y(n3835) );
  INVX1 U3663 ( .A(n3835), .Y(n3836) );
  AND2X2 U3664 ( .A(\mem<9><4> ), .B(n5061), .Y(n3837) );
  INVX1 U3665 ( .A(n3837), .Y(n3838) );
  AND2X2 U3666 ( .A(\mem<9><6> ), .B(n5061), .Y(n3839) );
  INVX1 U3667 ( .A(n3839), .Y(n3840) );
  AND2X2 U3668 ( .A(\mem<9><7> ), .B(n5062), .Y(n3841) );
  INVX1 U3669 ( .A(n3841), .Y(n3842) );
  AND2X2 U3670 ( .A(n782), .B(n3670), .Y(n3843) );
  AND2X2 U3671 ( .A(n6430), .B(n24), .Y(n3844) );
  AND2X2 U3672 ( .A(n911), .B(n3928), .Y(n3845) );
  INVX1 U3673 ( .A(n3845), .Y(n3846) );
  AND2X2 U3674 ( .A(n913), .B(n3927), .Y(n3847) );
  INVX1 U3675 ( .A(n3847), .Y(n3848) );
  OR2X2 U3676 ( .A(n5791), .B(n5790), .Y(n3849) );
  OR2X2 U3677 ( .A(n5887), .B(n5886), .Y(n3850) );
  OR2X2 U3678 ( .A(n5967), .B(n5966), .Y(n3851) );
  OR2X2 U3679 ( .A(n6107), .B(n6108), .Y(n3852) );
  OR2X2 U3680 ( .A(n6211), .B(n6210), .Y(n3853) );
  OR2X2 U3681 ( .A(n6258), .B(n6257), .Y(n3854) );
  OR2X2 U3682 ( .A(n6268), .B(n6267), .Y(n3855) );
  OR2X2 U3683 ( .A(n6337), .B(n6336), .Y(n3856) );
  OR2X2 U3684 ( .A(n6357), .B(n6356), .Y(n3857) );
  INVX1 U3685 ( .A(n714), .Y(n3858) );
  INVX1 U3686 ( .A(n715), .Y(n3859) );
  INVX1 U3687 ( .A(n729), .Y(n3860) );
  INVX1 U3688 ( .A(n743), .Y(n3861) );
  INVX1 U3689 ( .A(n766), .Y(n3862) );
  AND2X2 U3690 ( .A(\data_in<8> ), .B(n1573), .Y(n3863) );
  INVX1 U3691 ( .A(n3863), .Y(n3864) );
  AND2X2 U3692 ( .A(\data_in<9> ), .B(n1573), .Y(n3865) );
  INVX1 U3693 ( .A(n3865), .Y(n3866) );
  AND2X2 U3694 ( .A(\data_in<11> ), .B(n1573), .Y(n3867) );
  INVX1 U3695 ( .A(n3867), .Y(n3868) );
  AND2X2 U3696 ( .A(\data_in<12> ), .B(n1573), .Y(n3869) );
  INVX1 U3697 ( .A(n3869), .Y(n3870) );
  AND2X2 U3698 ( .A(\data_in<14> ), .B(n1573), .Y(n3871) );
  INVX1 U3699 ( .A(n3871), .Y(n3872) );
  AND2X2 U3700 ( .A(\data_in<15> ), .B(n1573), .Y(n3873) );
  INVX1 U3701 ( .A(n3873), .Y(n3874) );
  AND2X2 U3702 ( .A(n907), .B(n76), .Y(n3875) );
  INVX1 U3703 ( .A(n3875), .Y(n3876) );
  AND2X2 U3704 ( .A(n534), .B(n76), .Y(n3877) );
  INVX1 U3705 ( .A(n3877), .Y(n3878) );
  AND2X2 U3706 ( .A(n3914), .B(\data_in<0> ), .Y(n3879) );
  INVX1 U3707 ( .A(n3879), .Y(n3880) );
  AND2X2 U3708 ( .A(n108), .B(\data_in<1> ), .Y(n3881) );
  INVX1 U3709 ( .A(n3881), .Y(n3882) );
  AND2X2 U3710 ( .A(\data_in<2> ), .B(n3914), .Y(n3883) );
  INVX1 U3711 ( .A(n3883), .Y(n3884) );
  AND2X2 U3712 ( .A(\mem<39><2> ), .B(n5013), .Y(n3885) );
  INVX1 U3713 ( .A(n3885), .Y(n3886) );
  AND2X2 U3714 ( .A(\mem<39><5> ), .B(n5013), .Y(n3887) );
  INVX1 U3715 ( .A(n3887), .Y(n3888) );
  AND2X2 U3716 ( .A(\mem<35><2> ), .B(n5021), .Y(n3889) );
  INVX1 U3717 ( .A(n3889), .Y(n3890) );
  AND2X2 U3718 ( .A(\mem<35><5> ), .B(n5020), .Y(n3891) );
  INVX1 U3719 ( .A(n3891), .Y(n3892) );
  AND2X2 U3720 ( .A(\data_in<0> ), .B(n10), .Y(n3893) );
  INVX1 U3721 ( .A(n3893), .Y(n3894) );
  AND2X2 U3722 ( .A(\data_in<1> ), .B(n1635), .Y(n3895) );
  INVX1 U3723 ( .A(n3895), .Y(n3896) );
  AND2X2 U3724 ( .A(\data_in<2> ), .B(n1635), .Y(n3897) );
  INVX1 U3725 ( .A(n3897), .Y(n3898) );
  AND2X2 U3726 ( .A(\data_in<3> ), .B(n10), .Y(n3899) );
  INVX1 U3727 ( .A(n3899), .Y(n3900) );
  AND2X2 U3728 ( .A(\data_in<4> ), .B(n10), .Y(n3901) );
  INVX1 U3729 ( .A(n3901), .Y(n3902) );
  AND2X2 U3730 ( .A(\data_in<5> ), .B(n10), .Y(n3903) );
  INVX1 U3731 ( .A(n3903), .Y(n3904) );
  AND2X2 U3732 ( .A(\data_in<6> ), .B(n1635), .Y(n3905) );
  INVX1 U3733 ( .A(n3905), .Y(n3906) );
  AND2X2 U3734 ( .A(\data_in<7> ), .B(n1635), .Y(n3907) );
  INVX1 U3735 ( .A(n3907), .Y(n3908) );
  INVX1 U3736 ( .A(n5752), .Y(n3909) );
  INVX1 U3737 ( .A(n3659), .Y(n5754) );
  INVX1 U3738 ( .A(n904), .Y(n3910) );
  INVX1 U3739 ( .A(n3910), .Y(n3911) );
  INVX1 U3740 ( .A(n3910), .Y(n3912) );
  INVX1 U3741 ( .A(n497), .Y(n3913) );
  INVX1 U3742 ( .A(n517), .Y(n3914) );
  INVX1 U3743 ( .A(n517), .Y(n3915) );
  MUX2X1 U3744 ( .B(n5515), .A(n5514), .S(n5659), .Y(n5513) );
  INVX1 U3745 ( .A(n3948), .Y(n3917) );
  INVX1 U3746 ( .A(n3994), .Y(n3988) );
  INVX1 U3747 ( .A(n3919), .Y(n3918) );
  INVX1 U3748 ( .A(n5657), .Y(n3919) );
  MUX2X1 U3749 ( .B(\mem<23><7> ), .A(\mem<22><7> ), .S(n3988), .Y(n5627) );
  NAND2X1 U3750 ( .A(\mem<28><7> ), .B(n3920), .Y(n3921) );
  NAND2X1 U3751 ( .A(\mem<29><7> ), .B(n5690), .Y(n3922) );
  INVX1 U3752 ( .A(n106), .Y(n3920) );
  NAND2X1 U3753 ( .A(\mem<6><2> ), .B(n3954), .Y(n3923) );
  NAND2X1 U3754 ( .A(\mem<7><2> ), .B(n5680), .Y(n3924) );
  INVX1 U3755 ( .A(\addr<15> ), .Y(n3925) );
  INVX1 U3756 ( .A(n5183), .Y(n3926) );
  AND2X2 U3757 ( .A(n5711), .B(n3675), .Y(n3927) );
  AND2X2 U3758 ( .A(n3675), .B(n5157), .Y(n3928) );
  NAND2X1 U3759 ( .A(\mem<4><4> ), .B(n5170), .Y(n3929) );
  NAND2X1 U3760 ( .A(\mem<5><4> ), .B(n5689), .Y(n3930) );
  MUX2X1 U3761 ( .B(n5380), .A(n500), .S(n72), .Y(n5379) );
  MUX2X1 U3762 ( .B(n5327), .A(n5328), .S(n5665), .Y(n5326) );
  NAND2X1 U3763 ( .A(\mem<18><1> ), .B(n3931), .Y(n3932) );
  NAND2X1 U3764 ( .A(\mem<19><1> ), .B(n5687), .Y(n3933) );
  INVX1 U3765 ( .A(n5691), .Y(n3931) );
  INVX1 U3766 ( .A(n3940), .Y(n3935) );
  NAND2X1 U3767 ( .A(\mem<24><7> ), .B(n3988), .Y(n3936) );
  NAND2X1 U3768 ( .A(\mem<25><7> ), .B(n5686), .Y(n3937) );
  INVX2 U3769 ( .A(n5738), .Y(n5737) );
  INVX1 U3770 ( .A(n5705), .Y(n5738) );
  NAND2X1 U3771 ( .A(\mem<48><7> ), .B(n3947), .Y(n3938) );
  NAND2X1 U3772 ( .A(\mem<49><7> ), .B(n3935), .Y(n3939) );
  INVX1 U3773 ( .A(n5698), .Y(n3940) );
  NAND2X1 U3774 ( .A(\mem<46><3> ), .B(n3947), .Y(n3941) );
  NAND2X1 U3775 ( .A(\mem<47><3> ), .B(n5691), .Y(n3942) );
  MUX2X1 U3776 ( .B(n5598), .A(n5597), .S(n5658), .Y(n5596) );
  INVX1 U3777 ( .A(n5219), .Y(n3943) );
  NAND2X1 U3778 ( .A(\mem<26><1> ), .B(n3954), .Y(n3945) );
  NAND2X1 U3779 ( .A(\mem<27><1> ), .B(n5694), .Y(n3946) );
  MUX2X1 U3780 ( .B(\mem<61><3> ), .A(\mem<60><3> ), .S(n91), .Y(n5382) );
  MUX2X1 U3781 ( .B(\mem<27><2> ), .A(\mem<26><2> ), .S(n5186), .Y(n5359) );
  MUX2X1 U3782 ( .B(n508), .A(n5310), .S(n5661), .Y(n5309) );
  MUX2X1 U3783 ( .B(n510), .A(n5603), .S(n5671), .Y(n5602) );
  INVX1 U3784 ( .A(n5703), .Y(n5727) );
  MUX2X1 U3785 ( .B(n516), .A(n5382), .S(n5660), .Y(n5381) );
  MUX2X1 U3786 ( .B(n5640), .A(n5643), .S(n3949), .Y(n5647) );
  MUX2X1 U3787 ( .B(\mem<1><2> ), .A(\mem<0><2> ), .S(n3972), .Y(n5377) );
  NAND2X1 U3788 ( .A(\mem<62><3> ), .B(n3931), .Y(n3950) );
  NAND2X1 U3789 ( .A(\mem<63><3> ), .B(n5690), .Y(n3951) );
  NAND2X1 U3790 ( .A(\mem<10><4> ), .B(n3947), .Y(n3952) );
  NAND2X1 U3791 ( .A(\mem<11><4> ), .B(n3961), .Y(n3953) );
  INVX4 U3792 ( .A(n3990), .Y(n3954) );
  INVX2 U3793 ( .A(n3990), .Y(n5676) );
  INVX1 U3794 ( .A(n3948), .Y(n3955) );
  INVX1 U3795 ( .A(n5677), .Y(n5691) );
  MUX2X1 U3796 ( .B(\mem<51><4> ), .A(\mem<50><4> ), .S(n3947), .Y(n5438) );
  MUX2X1 U3797 ( .B(n5455), .A(n5458), .S(n3956), .Y(n5468) );
  MUX2X1 U3798 ( .B(n5596), .A(n5594), .S(n5654), .Y(n5606) );
  MUX2X1 U3799 ( .B(n535), .A(n5566), .S(n71), .Y(n5565) );
  INVX4 U3800 ( .A(n5722), .Y(n5726) );
  BUFX2 U3801 ( .A(n5190), .Y(n3958) );
  INVX1 U3802 ( .A(n5153), .Y(n5687) );
  INVX4 U3803 ( .A(n3995), .Y(n3961) );
  INVX4 U3804 ( .A(n3960), .Y(n5682) );
  MUX2X1 U3805 ( .B(n499), .A(n527), .S(n3959), .Y(N190) );
  INVX1 U3806 ( .A(n3964), .Y(n3960) );
  MUX2X1 U3807 ( .B(n5575), .A(n5574), .S(n5658), .Y(n5573) );
  INVX4 U3808 ( .A(n5651), .Y(n5653) );
  NAND2X1 U3809 ( .A(\mem<44><7> ), .B(n3997), .Y(n3962) );
  NAND2X1 U3810 ( .A(\mem<45><7> ), .B(n5686), .Y(n3963) );
  MUX2X1 U3811 ( .B(\mem<27><6> ), .A(\mem<26><6> ), .S(n3934), .Y(n5572) );
  MUX2X1 U3812 ( .B(n5608), .A(n521), .S(n5658), .Y(n5607) );
  MUX2X1 U3813 ( .B(\mem<34><3> ), .A(\mem<35><3> ), .S(n3989), .Y(n5396) );
  INVX1 U3814 ( .A(n5154), .Y(n3964) );
  INVX1 U3815 ( .A(n5756), .Y(n5698) );
  MUX2X1 U3816 ( .B(\mem<42><6> ), .A(\mem<43><6> ), .S(n3966), .Y(n5558) );
  INVX4 U3817 ( .A(n5697), .Y(n5168) );
  INVX1 U3818 ( .A(n5190), .Y(n3966) );
  OAI21X1 U3819 ( .A(n4218), .B(n5182), .C(n63), .Y(n3967) );
  OAI21X1 U3820 ( .A(n4218), .B(n5182), .C(n3912), .Y(n3968) );
  MUX2X1 U3821 ( .B(\mem<1><0> ), .A(\mem<0><0> ), .S(n3947), .Y(n5271) );
  INVX1 U3822 ( .A(\addr<15> ), .Y(n5183) );
  INVX8 U3823 ( .A(n87), .Y(n5751) );
  MUX2X1 U3824 ( .B(n5569), .A(n5568), .S(n5658), .Y(n5567) );
  MUX2X1 U3825 ( .B(n5409), .A(n5408), .S(n3969), .Y(n5407) );
  AND2X2 U3826 ( .A(n76), .B(n944), .Y(n3970) );
  INVX1 U3827 ( .A(n3995), .Y(n3971) );
  INVX1 U3828 ( .A(n3971), .Y(n3972) );
  INVX1 U3829 ( .A(n5173), .Y(n3973) );
  MUX2X1 U3830 ( .B(n5564), .A(n5563), .S(n3974), .Y(n5562) );
  MUX2X1 U3831 ( .B(\mem<21><0> ), .A(\mem<20><0> ), .S(n5170), .Y(n5254) );
  NAND2X1 U3832 ( .A(\mem<56><0> ), .B(n3988), .Y(n3975) );
  NAND2X1 U3833 ( .A(\mem<57><0> ), .B(n106), .Y(n3976) );
  MUX2X1 U3834 ( .B(\mem<45><3> ), .A(\mem<44><3> ), .S(n5676), .Y(n5389) );
  MUX2X1 U3835 ( .B(\mem<55><7> ), .A(\mem<54><7> ), .S(n3954), .Y(n5601) );
  NAND2X1 U3836 ( .A(\mem<60><7> ), .B(n3982), .Y(n3977) );
  NAND2X1 U3837 ( .A(\mem<61><7> ), .B(n5695), .Y(n3978) );
  NAND2X1 U3838 ( .A(\mem<28><1> ), .B(n3931), .Y(n3979) );
  NAND2X1 U3839 ( .A(\mem<29><1> ), .B(n5696), .Y(n3980) );
  INVX1 U3840 ( .A(n55), .Y(n3981) );
  MUX2X1 U3841 ( .B(\mem<53><3> ), .A(\mem<52><3> ), .S(n3954), .Y(n5385) );
  INVX4 U3842 ( .A(n5727), .Y(n5725) );
  INVX1 U3843 ( .A(n3971), .Y(n3982) );
  INVX1 U3844 ( .A(n6427), .Y(n3983) );
  INVX1 U3845 ( .A(n3948), .Y(n3984) );
  INVX1 U3846 ( .A(n5204), .Y(n3985) );
  MUX2X1 U3847 ( .B(\mem<63><7> ), .A(\mem<62><7> ), .S(n3954), .Y(n5595) );
  MUX2X1 U3848 ( .B(\mem<29><0> ), .A(\mem<28><0> ), .S(n3954), .Y(n5248) );
  MUX2X1 U3849 ( .B(n5272), .A(n5271), .S(n5661), .Y(n5270) );
  MUX2X1 U3850 ( .B(n5396), .A(n531), .S(n5660), .Y(n5395) );
  NAND2X1 U3851 ( .A(\mem<32><3> ), .B(n3954), .Y(n3986) );
  NAND2X1 U3852 ( .A(\mem<33><3> ), .B(n3961), .Y(n3987) );
  INVX1 U3853 ( .A(n5155), .Y(n3990) );
  INVX1 U3854 ( .A(n5153), .Y(n3991) );
  OR2X2 U3855 ( .A(n6083), .B(n5674), .Y(n5199) );
  INVX1 U3856 ( .A(n107), .Y(n5755) );
  MUX2X1 U3857 ( .B(n5555), .A(n5554), .S(n5659), .Y(n5553) );
  INVX1 U3858 ( .A(n107), .Y(n3993) );
  MUX2X1 U3859 ( .B(\mem<59><0> ), .A(\mem<58><0> ), .S(n3972), .Y(n5225) );
  INVX1 U3860 ( .A(n5666), .Y(n5195) );
  INVX1 U3861 ( .A(n5155), .Y(n3994) );
  INVX1 U3862 ( .A(n5755), .Y(n3995) );
  INVX1 U3863 ( .A(n5152), .Y(n5674) );
  INVX1 U3864 ( .A(n5653), .Y(n3996) );
  NAND2X1 U3865 ( .A(\mem<10><2> ), .B(n3997), .Y(n3998) );
  NAND2X1 U3866 ( .A(\mem<11><2> ), .B(n5692), .Y(n3999) );
  INVX1 U3867 ( .A(n3971), .Y(n3997) );
  AND2X2 U3868 ( .A(\mem<12><0> ), .B(n5057), .Y(n4000) );
  INVX1 U3869 ( .A(n4000), .Y(n4001) );
  AND2X2 U3870 ( .A(\mem<12><1> ), .B(n5058), .Y(n4002) );
  INVX1 U3871 ( .A(n4002), .Y(n4003) );
  AND2X2 U3872 ( .A(\mem<12><2> ), .B(n5057), .Y(n4004) );
  INVX1 U3873 ( .A(n4004), .Y(n4005) );
  AND2X2 U3874 ( .A(\mem<12><3> ), .B(n5058), .Y(n4006) );
  INVX1 U3875 ( .A(n4006), .Y(n4007) );
  AND2X2 U3876 ( .A(\mem<12><4> ), .B(n5057), .Y(n4008) );
  INVX1 U3877 ( .A(n4008), .Y(n4009) );
  AND2X2 U3878 ( .A(\mem<12><5> ), .B(n5058), .Y(n4010) );
  INVX1 U3879 ( .A(n4010), .Y(n4011) );
  AND2X2 U3880 ( .A(\mem<12><6> ), .B(n5057), .Y(n4012) );
  INVX1 U3881 ( .A(n4012), .Y(n4013) );
  AND2X2 U3882 ( .A(\mem<12><7> ), .B(n5058), .Y(n4014) );
  INVX1 U3883 ( .A(n4014), .Y(n4015) );
  AND2X2 U3884 ( .A(\mem<11><0> ), .B(n5059), .Y(n4016) );
  INVX1 U3885 ( .A(n4016), .Y(n4017) );
  AND2X2 U3886 ( .A(\mem<11><1> ), .B(n67), .Y(n4018) );
  INVX1 U3887 ( .A(n4018), .Y(n4019) );
  AND2X2 U3888 ( .A(\mem<11><2> ), .B(n67), .Y(n4020) );
  INVX1 U3889 ( .A(n4020), .Y(n4021) );
  AND2X2 U3890 ( .A(\mem<11><3> ), .B(n5059), .Y(n4022) );
  INVX1 U3891 ( .A(n4022), .Y(n4023) );
  AND2X2 U3892 ( .A(\mem<11><4> ), .B(n5059), .Y(n4024) );
  INVX1 U3893 ( .A(n4024), .Y(n4025) );
  AND2X2 U3894 ( .A(\mem<11><5> ), .B(n67), .Y(n4026) );
  INVX1 U3895 ( .A(n4026), .Y(n4027) );
  AND2X2 U3896 ( .A(\mem<11><6> ), .B(n5059), .Y(n4028) );
  INVX1 U3897 ( .A(n4028), .Y(n4029) );
  AND2X2 U3898 ( .A(\mem<11><7> ), .B(n67), .Y(n4030) );
  INVX1 U3899 ( .A(n4030), .Y(n4031) );
  AND2X2 U3900 ( .A(\mem<9><2> ), .B(n5061), .Y(n4032) );
  INVX1 U3901 ( .A(n4032), .Y(n4033) );
  AND2X2 U3902 ( .A(\mem<9><5> ), .B(n5062), .Y(n4034) );
  INVX1 U3903 ( .A(n4034), .Y(n4035) );
  OR2X2 U3904 ( .A(n5876), .B(n5877), .Y(n4036) );
  OR2X2 U3905 ( .A(n6119), .B(n6118), .Y(n4037) );
  OR2X2 U3906 ( .A(n6191), .B(n6190), .Y(n4038) );
  INVX1 U3907 ( .A(n813), .Y(n4039) );
  INVX1 U3908 ( .A(n844), .Y(n4040) );
  AND2X2 U3909 ( .A(\mem<29><3> ), .B(n233), .Y(n4041) );
  INVX1 U3910 ( .A(n4041), .Y(n4042) );
  AND2X2 U3911 ( .A(\mem<29><1> ), .B(n233), .Y(n4043) );
  INVX1 U3912 ( .A(n4043), .Y(n4044) );
  AND2X2 U3913 ( .A(\mem<61><0> ), .B(n5741), .Y(n4045) );
  INVX1 U3914 ( .A(n4045), .Y(n4046) );
  AND2X2 U3915 ( .A(\mem<2><0> ), .B(n5146), .Y(n4047) );
  INVX1 U3916 ( .A(n4047), .Y(n4048) );
  AND2X2 U3917 ( .A(\mem<42><0> ), .B(n5148), .Y(n4049) );
  INVX1 U3918 ( .A(n4049), .Y(n4050) );
  AND2X2 U3919 ( .A(\mem<2><1> ), .B(n5133), .Y(n4051) );
  INVX1 U3920 ( .A(n4051), .Y(n4052) );
  AND2X2 U3921 ( .A(\mem<42><1> ), .B(n5147), .Y(n4053) );
  INVX1 U3922 ( .A(n4053), .Y(n4054) );
  AND2X2 U3923 ( .A(\mem<43><1> ), .B(n196), .Y(n4055) );
  INVX1 U3924 ( .A(n4055), .Y(n4056) );
  AND2X2 U3925 ( .A(\mem<2><2> ), .B(n82), .Y(n4057) );
  INVX1 U3926 ( .A(n4057), .Y(n4058) );
  AND2X2 U3927 ( .A(\mem<42><2> ), .B(n166), .Y(n4059) );
  INVX1 U3928 ( .A(n4059), .Y(n4060) );
  AND2X2 U3929 ( .A(\mem<2><3> ), .B(n5133), .Y(n4061) );
  INVX1 U3930 ( .A(n4061), .Y(n4062) );
  AND2X2 U3931 ( .A(\mem<3><3> ), .B(n192), .Y(n4063) );
  INVX1 U3932 ( .A(n4063), .Y(n4064) );
  AND2X2 U3933 ( .A(\mem<42><3> ), .B(n5146), .Y(n4065) );
  INVX1 U3934 ( .A(n4065), .Y(n4066) );
  AND2X2 U3935 ( .A(\mem<2><4> ), .B(n5132), .Y(n4067) );
  INVX1 U3936 ( .A(n4067), .Y(n4068) );
  AND2X2 U3937 ( .A(\mem<42><4> ), .B(n5134), .Y(n4069) );
  INVX1 U3938 ( .A(n4069), .Y(n4070) );
  AND2X2 U3939 ( .A(\mem<43><4> ), .B(n192), .Y(n4071) );
  INVX1 U3940 ( .A(n4071), .Y(n4072) );
  AND2X2 U3941 ( .A(\mem<2><5> ), .B(n5142), .Y(n4073) );
  INVX1 U3942 ( .A(n4073), .Y(n4074) );
  AND2X2 U3943 ( .A(\mem<3><5> ), .B(n187), .Y(n4075) );
  INVX1 U3944 ( .A(n4075), .Y(n4076) );
  AND2X2 U3945 ( .A(\mem<42><5> ), .B(n166), .Y(n4077) );
  INVX1 U3946 ( .A(n4077), .Y(n4078) );
  AND2X2 U3947 ( .A(\mem<2><6> ), .B(n5126), .Y(n4079) );
  INVX1 U3948 ( .A(n4079), .Y(n4080) );
  AND2X2 U3949 ( .A(\mem<42><6> ), .B(n5131), .Y(n4081) );
  INVX1 U3950 ( .A(n4081), .Y(n4082) );
  AND2X2 U3951 ( .A(\mem<2><7> ), .B(n5137), .Y(n4083) );
  INVX1 U3952 ( .A(n4083), .Y(n4084) );
  AND2X2 U3953 ( .A(\mem<42><7> ), .B(n5131), .Y(n4085) );
  INVX1 U3954 ( .A(n4085), .Y(n4086) );
  AND2X2 U3955 ( .A(n5247), .B(n5657), .Y(n4087) );
  INVX1 U3956 ( .A(n4087), .Y(n4088) );
  AND2X2 U3957 ( .A(n5634), .B(n5652), .Y(n4089) );
  INVX1 U3958 ( .A(n4089), .Y(n4090) );
  AND2X2 U3959 ( .A(n5392), .B(n5655), .Y(n4091) );
  INVX1 U3960 ( .A(n4091), .Y(n4092) );
  AND2X2 U3961 ( .A(n5261), .B(n5657), .Y(n4093) );
  INVX1 U3962 ( .A(n4093), .Y(n4094) );
  AND2X2 U3963 ( .A(n5398), .B(n5655), .Y(n4095) );
  INVX1 U3964 ( .A(n4095), .Y(n4096) );
  AND2X2 U3965 ( .A(n5412), .B(n5655), .Y(n4097) );
  INVX1 U3966 ( .A(n4097), .Y(n4098) );
  AND2X2 U3967 ( .A(n5539), .B(n5653), .Y(n4099) );
  INVX1 U3968 ( .A(n4099), .Y(n4100) );
  AND2X2 U3969 ( .A(n5587), .B(n5653), .Y(n4101) );
  INVX1 U3970 ( .A(n4101), .Y(n4102) );
  AND2X2 U3971 ( .A(n5444), .B(n5217), .Y(n4103) );
  INVX1 U3972 ( .A(n4103), .Y(n4104) );
  OR2X2 U3973 ( .A(n5908), .B(n5907), .Y(n4105) );
  INVX1 U3974 ( .A(n4105), .Y(n4106) );
  OR2X2 U3975 ( .A(n6071), .B(n6070), .Y(n4107) );
  INVX1 U3976 ( .A(n4107), .Y(n4108) );
  OR2X2 U3977 ( .A(n6136), .B(n6135), .Y(n4109) );
  INVX1 U3978 ( .A(n4109), .Y(n4110) );
  AND2X2 U3979 ( .A(\mem<0><5> ), .B(n549), .Y(n4111) );
  INVX1 U3980 ( .A(n4111), .Y(n4112) );
  OR2X2 U3981 ( .A(n5716), .B(n5750), .Y(n4113) );
  INVX1 U3982 ( .A(n4113), .Y(n4114) );
  AND2X2 U3983 ( .A(n5250), .B(n5217), .Y(n4115) );
  INVX1 U3984 ( .A(n4115), .Y(n4116) );
  AND2X2 U3985 ( .A(n5301), .B(n5091), .Y(n4117) );
  INVX1 U3986 ( .A(n4117), .Y(n4118) );
  AND2X2 U3987 ( .A(n5295), .B(n5657), .Y(n4119) );
  INVX1 U3988 ( .A(n4119), .Y(n4120) );
  AND2X2 U3989 ( .A(n5298), .B(n5165), .Y(n4121) );
  INVX1 U3990 ( .A(n4121), .Y(n4122) );
  AND2X2 U3991 ( .A(n5289), .B(n5657), .Y(n4123) );
  INVX1 U3992 ( .A(n4123), .Y(n4124) );
  AND2X2 U3993 ( .A(n5292), .B(n5165), .Y(n4125) );
  INVX1 U3994 ( .A(n4125), .Y(n4126) );
  AND2X2 U3995 ( .A(n5582), .B(n5653), .Y(n4127) );
  INVX1 U3996 ( .A(n4127), .Y(n4128) );
  AND2X2 U3997 ( .A(n5585), .B(n5173), .Y(n4129) );
  INVX1 U3998 ( .A(n4129), .Y(n4130) );
  AND2X2 U3999 ( .A(n5637), .B(n5175), .Y(n4131) );
  INVX1 U4000 ( .A(n4131), .Y(n4132) );
  INVX1 U4001 ( .A(n4133), .Y(n4134) );
  AND2X2 U4002 ( .A(n5229), .B(n5191), .Y(n4135) );
  INVX1 U4003 ( .A(n4135), .Y(n4136) );
  AND2X2 U4004 ( .A(n5234), .B(n5657), .Y(n4137) );
  INVX1 U4005 ( .A(n4137), .Y(n4138) );
  AND2X2 U4006 ( .A(n5237), .B(n5191), .Y(n4139) );
  INVX1 U4007 ( .A(n4139), .Y(n4140) );
  AND2X2 U4008 ( .A(n5264), .B(n5191), .Y(n4141) );
  INVX1 U4009 ( .A(n4141), .Y(n4142) );
  AND2X2 U4010 ( .A(n5430), .B(n5208), .Y(n4143) );
  INVX1 U4011 ( .A(n4143), .Y(n4144) );
  INVX1 U4012 ( .A(n4145), .Y(n4146) );
  AND2X2 U4013 ( .A(n5401), .B(n5175), .Y(n4147) );
  INVX1 U4014 ( .A(n4147), .Y(n4148) );
  AND2X2 U4015 ( .A(n5415), .B(n5204), .Y(n4149) );
  INVX1 U4016 ( .A(n4149), .Y(n4150) );
  AND2X2 U4017 ( .A(n5542), .B(n5206), .Y(n4151) );
  INVX1 U4018 ( .A(n4151), .Y(n4152) );
  AND2X2 U4019 ( .A(n5590), .B(n5209), .Y(n4153) );
  INVX1 U4020 ( .A(n4153), .Y(n4154) );
  AND2X2 U4021 ( .A(n5441), .B(n3973), .Y(n4155) );
  INVX1 U4022 ( .A(n4155), .Y(n4156) );
  AND2X2 U4023 ( .A(n5424), .B(n5084), .Y(n4157) );
  INVX1 U4024 ( .A(n4157), .Y(n4158) );
  AND2X2 U4025 ( .A(\mem<0><1> ), .B(n549), .Y(n4159) );
  INVX1 U4026 ( .A(n4159), .Y(n4160) );
  AND2X2 U4027 ( .A(\mem<0><3> ), .B(n549), .Y(n4161) );
  INVX1 U4028 ( .A(n4161), .Y(n4162) );
  AND2X2 U4029 ( .A(\mem<61><7> ), .B(n233), .Y(n4163) );
  INVX1 U4030 ( .A(n4163), .Y(n4164) );
  INVX1 U4031 ( .A(\addr<6> ), .Y(n4165) );
  INVX1 U4032 ( .A(\addr<8> ), .Y(n4166) );
  BUFX2 U4033 ( .A(n5774), .Y(n4167) );
  INVX1 U4034 ( .A(n5844), .Y(n4168) );
  INVX1 U4035 ( .A(n4168), .Y(n4169) );
  AND2X2 U4036 ( .A(n5843), .B(n629), .Y(n4170) );
  INVX1 U4037 ( .A(n4170), .Y(n4171) );
  INVX1 U4038 ( .A(n4173), .Y(n4172) );
  AND2X2 U4039 ( .A(n5843), .B(n630), .Y(n4173) );
  AND2X2 U4040 ( .A(N181), .B(n630), .Y(n4174) );
  INVX1 U4041 ( .A(n4174), .Y(n4175) );
  INVX1 U4042 ( .A(n5725), .Y(n5724) );
  INVX1 U4043 ( .A(n3970), .Y(n4176) );
  AND2X2 U4044 ( .A(\mem<61><1> ), .B(n5741), .Y(n4177) );
  AND2X2 U4045 ( .A(\mem<61><2> ), .B(n5741), .Y(n4178) );
  INVX1 U4046 ( .A(n4178), .Y(n4179) );
  AND2X2 U4047 ( .A(\mem<61><3> ), .B(n5741), .Y(n4180) );
  AND2X2 U4048 ( .A(\mem<60><3> ), .B(n163), .Y(n4181) );
  AND2X2 U4049 ( .A(\mem<61><4> ), .B(n5741), .Y(n4182) );
  INVX1 U4050 ( .A(n4182), .Y(n4183) );
  AND2X2 U4051 ( .A(\mem<61><5> ), .B(n5741), .Y(n4184) );
  AND2X2 U4052 ( .A(\mem<60><5> ), .B(n151), .Y(n4185) );
  AND2X2 U4053 ( .A(\mem<61><6> ), .B(n233), .Y(n4186) );
  INVX1 U4054 ( .A(n4186), .Y(n4187) );
  AND2X2 U4055 ( .A(\mem<0><6> ), .B(n549), .Y(n4188) );
  INVX1 U4056 ( .A(n4188), .Y(n4189) );
  AND2X2 U4057 ( .A(\mem<0><7> ), .B(n549), .Y(n4190) );
  INVX1 U4058 ( .A(n4190), .Y(n4191) );
  INVX1 U4059 ( .A(n883), .Y(n4192) );
  AND2X2 U4060 ( .A(\data_in<0> ), .B(n1647), .Y(n4193) );
  INVX1 U4061 ( .A(n4193), .Y(n4194) );
  AND2X2 U4062 ( .A(\data_in<1> ), .B(n1647), .Y(n4195) );
  INVX1 U4063 ( .A(n4195), .Y(n4196) );
  AND2X2 U4064 ( .A(\data_in<2> ), .B(n1647), .Y(n4197) );
  INVX1 U4065 ( .A(n4197), .Y(n4198) );
  AND2X2 U4066 ( .A(\data_in<3> ), .B(n1647), .Y(n4199) );
  INVX1 U4067 ( .A(n4199), .Y(n4200) );
  AND2X2 U4068 ( .A(\data_in<4> ), .B(n1647), .Y(n4201) );
  INVX1 U4069 ( .A(n4201), .Y(n4202) );
  AND2X2 U4070 ( .A(\data_in<5> ), .B(n1647), .Y(n4203) );
  INVX1 U4071 ( .A(n4203), .Y(n4204) );
  AND2X2 U4072 ( .A(\data_in<6> ), .B(n1647), .Y(n4205) );
  INVX1 U4073 ( .A(n4205), .Y(n4206) );
  AND2X2 U4074 ( .A(\data_in<7> ), .B(n1647), .Y(n4207) );
  INVX1 U4075 ( .A(n4207), .Y(n4208) );
  AND2X2 U4076 ( .A(n20), .B(n6440), .Y(n4209) );
  INVX1 U4077 ( .A(n6163), .Y(n4210) );
  INVX1 U4078 ( .A(n4210), .Y(n4211) );
  INVX1 U4079 ( .A(n5941), .Y(n4212) );
  INVX1 U4080 ( .A(n4212), .Y(n4213) );
  INVX1 U4081 ( .A(n6093), .Y(n4214) );
  INVX1 U4082 ( .A(n4214), .Y(n4215) );
  INVX1 U4083 ( .A(n6244), .Y(n4216) );
  AND2X2 U4084 ( .A(n5141), .B(n6457), .Y(n4217) );
  INVX1 U4085 ( .A(n4217), .Y(n4218) );
  INVX1 U4086 ( .A(n5830), .Y(n4219) );
  INVX1 U4087 ( .A(n4219), .Y(n4220) );
  OR2X2 U4088 ( .A(n5773), .B(N182), .Y(n4221) );
  OR2X2 U4089 ( .A(n5802), .B(n5801), .Y(n4222) );
  AND2X2 U4090 ( .A(\mem<59><2> ), .B(n194), .Y(n4223) );
  INVX1 U4091 ( .A(n4223), .Y(n4224) );
  OR2X2 U4092 ( .A(n6041), .B(n6042), .Y(n4225) );
  AND2X2 U4093 ( .A(\mem<59><4> ), .B(n191), .Y(n4226) );
  INVX1 U4094 ( .A(n4226), .Y(n4227) );
  AND2X2 U4095 ( .A(\mem<0><4> ), .B(n549), .Y(n4228) );
  INVX1 U4096 ( .A(n4228), .Y(n4229) );
  AND2X2 U4097 ( .A(\mem<59><6> ), .B(n190), .Y(n4230) );
  INVX1 U4098 ( .A(n4230), .Y(n4231) );
  OR2X2 U4099 ( .A(n6288), .B(n6287), .Y(n4232) );
  OR2X2 U4100 ( .A(n6347), .B(n6346), .Y(n4233) );
  OR2X2 U4101 ( .A(n6368), .B(n6367), .Y(n4234) );
  AND2X2 U4102 ( .A(\data_in<8> ), .B(n1648), .Y(n4235) );
  INVX1 U4103 ( .A(n4235), .Y(n4236) );
  AND2X2 U4104 ( .A(\data_in<9> ), .B(n1648), .Y(n4237) );
  INVX1 U4105 ( .A(n4237), .Y(n4238) );
  AND2X2 U4106 ( .A(\data_in<10> ), .B(n1648), .Y(n4239) );
  INVX1 U4107 ( .A(n4239), .Y(n4240) );
  AND2X2 U4108 ( .A(\data_in<11> ), .B(n1648), .Y(n4241) );
  INVX1 U4109 ( .A(n4241), .Y(n4242) );
  AND2X2 U4110 ( .A(\data_in<12> ), .B(n1648), .Y(n4243) );
  INVX1 U4111 ( .A(n4243), .Y(n4244) );
  AND2X2 U4112 ( .A(\data_in<13> ), .B(n1648), .Y(n4245) );
  INVX1 U4113 ( .A(n4245), .Y(n4246) );
  AND2X2 U4114 ( .A(\data_in<14> ), .B(n1648), .Y(n4247) );
  INVX1 U4115 ( .A(n4247), .Y(n4248) );
  AND2X2 U4116 ( .A(\data_in<15> ), .B(n1648), .Y(n4249) );
  INVX1 U4117 ( .A(n4249), .Y(n4250) );
  OR2X2 U4118 ( .A(n5824), .B(n5823), .Y(n4251) );
  AND2X2 U4119 ( .A(\mem<0><2> ), .B(n549), .Y(n4252) );
  INVX1 U4120 ( .A(n4252), .Y(n4253) );
  AND2X2 U4121 ( .A(\mem<63><0> ), .B(n4970), .Y(n4254) );
  INVX1 U4122 ( .A(n4254), .Y(n4255) );
  AND2X2 U4123 ( .A(\mem<63><1> ), .B(n4969), .Y(n4256) );
  INVX1 U4124 ( .A(n4256), .Y(n4257) );
  AND2X2 U4125 ( .A(\mem<63><2> ), .B(n4969), .Y(n4258) );
  INVX1 U4126 ( .A(n4258), .Y(n4259) );
  AND2X2 U4127 ( .A(\mem<63><3> ), .B(n4969), .Y(n4260) );
  INVX1 U4128 ( .A(n4260), .Y(n4261) );
  AND2X2 U4129 ( .A(\mem<63><4> ), .B(n4969), .Y(n4262) );
  INVX1 U4130 ( .A(n4262), .Y(n4263) );
  AND2X2 U4131 ( .A(\mem<63><5> ), .B(n4970), .Y(n4264) );
  INVX1 U4132 ( .A(n4264), .Y(n4265) );
  AND2X2 U4133 ( .A(\mem<63><6> ), .B(n4970), .Y(n4266) );
  INVX1 U4134 ( .A(n4266), .Y(n4267) );
  AND2X2 U4135 ( .A(\mem<63><7> ), .B(n4970), .Y(n4268) );
  INVX1 U4136 ( .A(n4268), .Y(n4269) );
  AND2X2 U4137 ( .A(\mem<62><0> ), .B(n4972), .Y(n4270) );
  INVX1 U4138 ( .A(n4270), .Y(n4271) );
  AND2X2 U4139 ( .A(\mem<62><1> ), .B(n4971), .Y(n4272) );
  INVX1 U4140 ( .A(n4272), .Y(n4273) );
  AND2X2 U4141 ( .A(\mem<62><2> ), .B(n4971), .Y(n4274) );
  INVX1 U4142 ( .A(n4274), .Y(n4275) );
  AND2X2 U4143 ( .A(\mem<62><3> ), .B(n4971), .Y(n4276) );
  INVX1 U4144 ( .A(n4276), .Y(n4277) );
  AND2X2 U4145 ( .A(\mem<62><4> ), .B(n4971), .Y(n4278) );
  INVX1 U4146 ( .A(n4278), .Y(n4279) );
  AND2X2 U4147 ( .A(\mem<62><5> ), .B(n4972), .Y(n4280) );
  INVX1 U4148 ( .A(n4280), .Y(n4281) );
  AND2X2 U4149 ( .A(\mem<62><6> ), .B(n4972), .Y(n4282) );
  INVX1 U4150 ( .A(n4282), .Y(n4283) );
  AND2X2 U4151 ( .A(\mem<62><7> ), .B(n4972), .Y(n4284) );
  INVX1 U4152 ( .A(n4284), .Y(n4285) );
  AND2X2 U4153 ( .A(\mem<61><0> ), .B(n4973), .Y(n4286) );
  INVX1 U4154 ( .A(n4286), .Y(n4287) );
  AND2X2 U4155 ( .A(\mem<61><1> ), .B(n4974), .Y(n4288) );
  INVX1 U4156 ( .A(n4288), .Y(n4289) );
  AND2X2 U4157 ( .A(\mem<61><2> ), .B(n4973), .Y(n4290) );
  INVX1 U4158 ( .A(n4290), .Y(n4291) );
  AND2X2 U4159 ( .A(\mem<61><3> ), .B(n4974), .Y(n4292) );
  INVX1 U4160 ( .A(n4292), .Y(n4293) );
  AND2X2 U4161 ( .A(\mem<61><4> ), .B(n4973), .Y(n4294) );
  INVX1 U4162 ( .A(n4294), .Y(n4295) );
  AND2X2 U4163 ( .A(\mem<61><5> ), .B(n4974), .Y(n4296) );
  INVX1 U4164 ( .A(n4296), .Y(n4297) );
  AND2X2 U4165 ( .A(\mem<61><6> ), .B(n4973), .Y(n4298) );
  INVX1 U4166 ( .A(n4298), .Y(n4299) );
  AND2X2 U4167 ( .A(\mem<61><7> ), .B(n4974), .Y(n4300) );
  INVX1 U4168 ( .A(n4300), .Y(n4301) );
  AND2X2 U4169 ( .A(\mem<60><0> ), .B(n4975), .Y(n4302) );
  INVX1 U4170 ( .A(n4302), .Y(n4303) );
  AND2X2 U4171 ( .A(\mem<60><1> ), .B(n4976), .Y(n4304) );
  INVX1 U4172 ( .A(n4304), .Y(n4305) );
  AND2X2 U4173 ( .A(\mem<60><2> ), .B(n4975), .Y(n4306) );
  INVX1 U4174 ( .A(n4306), .Y(n4307) );
  AND2X2 U4175 ( .A(\mem<60><3> ), .B(n4976), .Y(n4308) );
  INVX1 U4176 ( .A(n4308), .Y(n4309) );
  AND2X2 U4177 ( .A(\mem<60><4> ), .B(n4975), .Y(n4310) );
  INVX1 U4178 ( .A(n4310), .Y(n4311) );
  AND2X2 U4179 ( .A(\mem<60><5> ), .B(n4976), .Y(n4312) );
  INVX1 U4180 ( .A(n4312), .Y(n4313) );
  AND2X2 U4181 ( .A(\mem<60><6> ), .B(n4975), .Y(n4314) );
  INVX1 U4182 ( .A(n4314), .Y(n4315) );
  AND2X2 U4183 ( .A(\mem<60><7> ), .B(n4976), .Y(n4316) );
  INVX1 U4184 ( .A(n4316), .Y(n4317) );
  AND2X2 U4185 ( .A(\mem<59><0> ), .B(n4977), .Y(n4318) );
  INVX1 U4186 ( .A(n4318), .Y(n4319) );
  AND2X2 U4187 ( .A(\mem<59><1> ), .B(n4978), .Y(n4320) );
  INVX1 U4188 ( .A(n4320), .Y(n4321) );
  AND2X2 U4189 ( .A(\mem<59><2> ), .B(n4977), .Y(n4322) );
  INVX1 U4190 ( .A(n4322), .Y(n4323) );
  AND2X2 U4191 ( .A(\mem<59><3> ), .B(n4978), .Y(n4324) );
  INVX1 U4192 ( .A(n4324), .Y(n4325) );
  AND2X2 U4193 ( .A(\mem<59><4> ), .B(n4977), .Y(n4326) );
  INVX1 U4194 ( .A(n4326), .Y(n4327) );
  AND2X2 U4195 ( .A(\mem<59><5> ), .B(n4978), .Y(n4328) );
  INVX1 U4196 ( .A(n4328), .Y(n4329) );
  AND2X2 U4197 ( .A(\mem<59><6> ), .B(n4977), .Y(n4330) );
  INVX1 U4198 ( .A(n4330), .Y(n4331) );
  AND2X2 U4199 ( .A(\mem<59><7> ), .B(n4978), .Y(n4332) );
  INVX1 U4200 ( .A(n4332), .Y(n4333) );
  AND2X2 U4201 ( .A(\mem<58><0> ), .B(n4979), .Y(n4334) );
  INVX1 U4202 ( .A(n4334), .Y(n4335) );
  AND2X2 U4203 ( .A(\mem<58><1> ), .B(n4980), .Y(n4336) );
  INVX1 U4204 ( .A(n4336), .Y(n4337) );
  AND2X2 U4205 ( .A(\mem<58><2> ), .B(n4979), .Y(n4338) );
  INVX1 U4206 ( .A(n4338), .Y(n4339) );
  AND2X2 U4207 ( .A(\mem<58><3> ), .B(n4979), .Y(n4340) );
  INVX1 U4208 ( .A(n4340), .Y(n4341) );
  AND2X2 U4209 ( .A(\mem<58><4> ), .B(n4980), .Y(n4342) );
  INVX1 U4210 ( .A(n4342), .Y(n4343) );
  AND2X2 U4211 ( .A(\mem<58><5> ), .B(n4980), .Y(n4344) );
  INVX1 U4212 ( .A(n4344), .Y(n4345) );
  AND2X2 U4213 ( .A(\mem<58><6> ), .B(n4979), .Y(n4346) );
  INVX1 U4214 ( .A(n4346), .Y(n4347) );
  AND2X2 U4215 ( .A(\mem<58><7> ), .B(n4980), .Y(n4348) );
  INVX1 U4216 ( .A(n4348), .Y(n4349) );
  AND2X2 U4217 ( .A(\mem<57><0> ), .B(n4981), .Y(n4350) );
  INVX1 U4218 ( .A(n4350), .Y(n4351) );
  AND2X2 U4219 ( .A(\mem<57><1> ), .B(n4982), .Y(n4352) );
  INVX1 U4220 ( .A(n4352), .Y(n4353) );
  AND2X2 U4221 ( .A(\mem<57><2> ), .B(n4981), .Y(n4354) );
  INVX1 U4222 ( .A(n4354), .Y(n4355) );
  AND2X2 U4223 ( .A(\mem<57><3> ), .B(n4982), .Y(n4356) );
  INVX1 U4224 ( .A(n4356), .Y(n4357) );
  AND2X2 U4225 ( .A(\mem<57><4> ), .B(n4981), .Y(n4358) );
  INVX1 U4226 ( .A(n4358), .Y(n4359) );
  AND2X2 U4227 ( .A(\mem<57><5> ), .B(n4982), .Y(n4360) );
  INVX1 U4228 ( .A(n4360), .Y(n4361) );
  AND2X2 U4229 ( .A(\mem<57><6> ), .B(n4981), .Y(n4362) );
  INVX1 U4230 ( .A(n4362), .Y(n4363) );
  AND2X2 U4231 ( .A(\mem<57><7> ), .B(n4982), .Y(n4364) );
  INVX1 U4232 ( .A(n4364), .Y(n4365) );
  AND2X2 U4233 ( .A(\mem<55><0> ), .B(n4986), .Y(n4366) );
  INVX1 U4234 ( .A(n4366), .Y(n4367) );
  AND2X2 U4235 ( .A(\mem<55><1> ), .B(n4987), .Y(n4368) );
  INVX1 U4236 ( .A(n4368), .Y(n4369) );
  AND2X2 U4237 ( .A(\mem<55><2> ), .B(n4987), .Y(n4370) );
  INVX1 U4238 ( .A(n4370), .Y(n4371) );
  AND2X2 U4239 ( .A(\mem<55><3> ), .B(n4986), .Y(n4372) );
  INVX1 U4240 ( .A(n4372), .Y(n4373) );
  AND2X2 U4241 ( .A(\mem<55><4> ), .B(n4987), .Y(n4374) );
  INVX1 U4242 ( .A(n4374), .Y(n4375) );
  AND2X2 U4243 ( .A(\mem<55><5> ), .B(n4986), .Y(n4376) );
  INVX1 U4244 ( .A(n4376), .Y(n4377) );
  AND2X2 U4245 ( .A(\mem<55><6> ), .B(n4986), .Y(n4378) );
  INVX1 U4246 ( .A(n4378), .Y(n4379) );
  AND2X2 U4247 ( .A(\mem<55><7> ), .B(n4987), .Y(n4380) );
  INVX1 U4248 ( .A(n4380), .Y(n4381) );
  AND2X2 U4249 ( .A(\mem<54><0> ), .B(n4988), .Y(n4382) );
  INVX1 U4250 ( .A(n4382), .Y(n4383) );
  AND2X2 U4251 ( .A(\mem<54><1> ), .B(n4989), .Y(n4384) );
  INVX1 U4252 ( .A(n4384), .Y(n4385) );
  AND2X2 U4253 ( .A(\mem<54><2> ), .B(n4988), .Y(n4386) );
  INVX1 U4254 ( .A(n4386), .Y(n4387) );
  AND2X2 U4255 ( .A(\mem<54><3> ), .B(n4989), .Y(n4388) );
  INVX1 U4256 ( .A(n4388), .Y(n4389) );
  AND2X2 U4257 ( .A(\mem<54><4> ), .B(n4988), .Y(n4390) );
  INVX1 U4258 ( .A(n4390), .Y(n4391) );
  AND2X2 U4259 ( .A(\mem<54><5> ), .B(n4989), .Y(n4392) );
  INVX1 U4260 ( .A(n4392), .Y(n4393) );
  AND2X2 U4261 ( .A(\mem<54><6> ), .B(n4988), .Y(n4394) );
  INVX1 U4262 ( .A(n4394), .Y(n4395) );
  AND2X2 U4263 ( .A(\mem<54><7> ), .B(n4989), .Y(n4396) );
  INVX1 U4264 ( .A(n4396), .Y(n4397) );
  AND2X2 U4265 ( .A(\mem<53><0> ), .B(n4990), .Y(n4398) );
  INVX1 U4266 ( .A(n4398), .Y(n4399) );
  AND2X2 U4267 ( .A(\mem<53><1> ), .B(n4991), .Y(n4400) );
  INVX1 U4268 ( .A(n4400), .Y(n4401) );
  AND2X2 U4269 ( .A(\mem<53><2> ), .B(n4990), .Y(n4402) );
  INVX1 U4270 ( .A(n4402), .Y(n4403) );
  AND2X2 U4271 ( .A(\mem<53><3> ), .B(n4991), .Y(n4404) );
  INVX1 U4272 ( .A(n4404), .Y(n4405) );
  AND2X2 U4273 ( .A(\mem<53><4> ), .B(n4990), .Y(n4406) );
  INVX1 U4274 ( .A(n4406), .Y(n4407) );
  AND2X2 U4275 ( .A(\mem<53><5> ), .B(n4991), .Y(n4408) );
  INVX1 U4276 ( .A(n4408), .Y(n4409) );
  AND2X2 U4277 ( .A(\mem<53><6> ), .B(n4990), .Y(n4410) );
  INVX1 U4278 ( .A(n4410), .Y(n4411) );
  AND2X2 U4279 ( .A(\mem<53><7> ), .B(n4991), .Y(n4412) );
  INVX1 U4280 ( .A(n4412), .Y(n4413) );
  AND2X2 U4281 ( .A(\mem<52><0> ), .B(n4992), .Y(n4414) );
  INVX1 U4282 ( .A(n4414), .Y(n4415) );
  AND2X2 U4283 ( .A(\mem<52><1> ), .B(n4993), .Y(n4416) );
  INVX1 U4284 ( .A(n4416), .Y(n4417) );
  AND2X2 U4285 ( .A(\mem<52><2> ), .B(n4993), .Y(n4418) );
  INVX1 U4286 ( .A(n4418), .Y(n4419) );
  AND2X2 U4287 ( .A(\mem<52><3> ), .B(n4992), .Y(n4420) );
  INVX1 U4288 ( .A(n4420), .Y(n4421) );
  AND2X2 U4289 ( .A(\mem<52><4> ), .B(n4993), .Y(n4422) );
  INVX1 U4290 ( .A(n4422), .Y(n4423) );
  AND2X2 U4291 ( .A(\mem<52><5> ), .B(n4992), .Y(n4424) );
  INVX1 U4292 ( .A(n4424), .Y(n4425) );
  AND2X2 U4293 ( .A(\mem<52><6> ), .B(n4992), .Y(n4426) );
  INVX1 U4294 ( .A(n4426), .Y(n4427) );
  AND2X2 U4295 ( .A(\mem<52><7> ), .B(n4993), .Y(n4428) );
  INVX1 U4296 ( .A(n4428), .Y(n4429) );
  AND2X2 U4297 ( .A(\mem<51><0> ), .B(n60), .Y(n4430) );
  INVX1 U4298 ( .A(n4430), .Y(n4431) );
  AND2X2 U4299 ( .A(\mem<51><1> ), .B(n60), .Y(n4432) );
  INVX1 U4300 ( .A(n4432), .Y(n4433) );
  AND2X2 U4301 ( .A(\mem<51><2> ), .B(n60), .Y(n4434) );
  INVX1 U4302 ( .A(n4434), .Y(n4435) );
  AND2X2 U4303 ( .A(\mem<51><3> ), .B(n60), .Y(n4436) );
  INVX1 U4304 ( .A(n4436), .Y(n4437) );
  AND2X2 U4305 ( .A(\mem<51><4> ), .B(n60), .Y(n4438) );
  INVX1 U4306 ( .A(n4438), .Y(n4439) );
  AND2X2 U4307 ( .A(\mem<51><5> ), .B(n60), .Y(n4440) );
  INVX1 U4308 ( .A(n4440), .Y(n4441) );
  AND2X2 U4309 ( .A(\mem<51><6> ), .B(n60), .Y(n4442) );
  INVX1 U4310 ( .A(n4442), .Y(n4443) );
  AND2X2 U4311 ( .A(\mem<51><7> ), .B(n60), .Y(n4444) );
  INVX1 U4312 ( .A(n4444), .Y(n4445) );
  AND2X2 U4313 ( .A(\mem<50><0> ), .B(n4994), .Y(n4446) );
  INVX1 U4314 ( .A(n4446), .Y(n4447) );
  AND2X2 U4315 ( .A(\mem<50><1> ), .B(n4995), .Y(n4448) );
  INVX1 U4316 ( .A(n4448), .Y(n4449) );
  AND2X2 U4317 ( .A(\mem<50><2> ), .B(n4994), .Y(n4450) );
  INVX1 U4318 ( .A(n4450), .Y(n4451) );
  AND2X2 U4319 ( .A(\mem<50><3> ), .B(n4995), .Y(n4452) );
  INVX1 U4320 ( .A(n4452), .Y(n4453) );
  AND2X2 U4321 ( .A(\mem<50><4> ), .B(n4994), .Y(n4454) );
  INVX1 U4322 ( .A(n4454), .Y(n4455) );
  AND2X2 U4323 ( .A(\mem<50><5> ), .B(n4995), .Y(n4456) );
  INVX1 U4324 ( .A(n4456), .Y(n4457) );
  AND2X2 U4325 ( .A(\mem<50><6> ), .B(n4994), .Y(n4458) );
  INVX1 U4326 ( .A(n4458), .Y(n4459) );
  AND2X2 U4327 ( .A(\mem<50><7> ), .B(n4995), .Y(n4460) );
  INVX1 U4328 ( .A(n4460), .Y(n4461) );
  AND2X2 U4329 ( .A(\mem<49><0> ), .B(n4996), .Y(n4462) );
  INVX1 U4330 ( .A(n4462), .Y(n4463) );
  AND2X2 U4331 ( .A(\mem<49><1> ), .B(n4997), .Y(n4464) );
  INVX1 U4332 ( .A(n4464), .Y(n4465) );
  AND2X2 U4333 ( .A(\mem<49><2> ), .B(n4996), .Y(n4466) );
  INVX1 U4334 ( .A(n4466), .Y(n4467) );
  AND2X2 U4335 ( .A(\mem<49><3> ), .B(n4997), .Y(n4468) );
  INVX1 U4336 ( .A(n4468), .Y(n4469) );
  AND2X2 U4337 ( .A(\mem<49><4> ), .B(n4996), .Y(n4470) );
  INVX1 U4338 ( .A(n4470), .Y(n4471) );
  AND2X2 U4339 ( .A(\mem<49><5> ), .B(n4997), .Y(n4472) );
  INVX1 U4340 ( .A(n4472), .Y(n4473) );
  AND2X2 U4341 ( .A(\mem<49><6> ), .B(n4996), .Y(n4474) );
  INVX1 U4342 ( .A(n4474), .Y(n4475) );
  AND2X2 U4343 ( .A(\mem<49><7> ), .B(n4997), .Y(n4476) );
  INVX1 U4344 ( .A(n4476), .Y(n4477) );
  AND2X2 U4345 ( .A(\mem<40><0> ), .B(n5012), .Y(n4478) );
  INVX1 U4346 ( .A(n4478), .Y(n4479) );
  AND2X2 U4347 ( .A(\mem<40><1> ), .B(n5012), .Y(n4480) );
  INVX1 U4348 ( .A(n4480), .Y(n4481) );
  AND2X2 U4349 ( .A(\mem<40><2> ), .B(n5012), .Y(n4482) );
  INVX1 U4350 ( .A(n4482), .Y(n4483) );
  AND2X2 U4351 ( .A(\mem<40><3> ), .B(n5012), .Y(n4484) );
  INVX1 U4352 ( .A(n4484), .Y(n4485) );
  AND2X2 U4353 ( .A(\mem<40><4> ), .B(n5012), .Y(n4486) );
  INVX1 U4354 ( .A(n4486), .Y(n4487) );
  AND2X2 U4355 ( .A(\mem<40><5> ), .B(n5012), .Y(n4488) );
  INVX1 U4356 ( .A(n4488), .Y(n4489) );
  AND2X2 U4357 ( .A(\mem<40><6> ), .B(n5012), .Y(n4490) );
  INVX1 U4358 ( .A(n4490), .Y(n4491) );
  AND2X2 U4359 ( .A(\mem<40><7> ), .B(n5012), .Y(n4492) );
  INVX1 U4360 ( .A(n4492), .Y(n4493) );
  AND2X2 U4361 ( .A(\mem<39><0> ), .B(n5013), .Y(n4494) );
  INVX1 U4362 ( .A(n4494), .Y(n4495) );
  AND2X2 U4363 ( .A(\mem<39><1> ), .B(n5013), .Y(n4496) );
  INVX1 U4364 ( .A(n4496), .Y(n4497) );
  AND2X2 U4365 ( .A(\mem<39><3> ), .B(n5013), .Y(n4498) );
  INVX1 U4366 ( .A(n4498), .Y(n4499) );
  AND2X2 U4367 ( .A(\mem<39><4> ), .B(n5013), .Y(n4500) );
  INVX1 U4368 ( .A(n4500), .Y(n4501) );
  AND2X2 U4369 ( .A(\mem<39><6> ), .B(n5013), .Y(n4502) );
  INVX1 U4370 ( .A(n4502), .Y(n4503) );
  AND2X2 U4371 ( .A(\mem<39><7> ), .B(n5013), .Y(n4504) );
  INVX1 U4372 ( .A(n4504), .Y(n4505) );
  AND2X2 U4373 ( .A(\mem<38><0> ), .B(n5014), .Y(n4506) );
  INVX1 U4374 ( .A(n4506), .Y(n4507) );
  AND2X2 U4375 ( .A(\mem<38><1> ), .B(n5015), .Y(n4508) );
  INVX1 U4376 ( .A(n4508), .Y(n4509) );
  AND2X2 U4377 ( .A(\mem<38><2> ), .B(n5014), .Y(n4510) );
  INVX1 U4378 ( .A(n4510), .Y(n4511) );
  AND2X2 U4379 ( .A(\mem<38><3> ), .B(n5015), .Y(n4512) );
  INVX1 U4380 ( .A(n4512), .Y(n4513) );
  AND2X2 U4381 ( .A(\mem<38><4> ), .B(n5014), .Y(n4514) );
  INVX1 U4382 ( .A(n4514), .Y(n4515) );
  AND2X2 U4383 ( .A(\mem<38><5> ), .B(n5015), .Y(n4516) );
  INVX1 U4384 ( .A(n4516), .Y(n4517) );
  AND2X2 U4385 ( .A(\mem<38><6> ), .B(n5014), .Y(n4518) );
  INVX1 U4386 ( .A(n4518), .Y(n4519) );
  AND2X2 U4387 ( .A(\mem<38><7> ), .B(n5015), .Y(n4520) );
  INVX1 U4388 ( .A(n4520), .Y(n4521) );
  AND2X2 U4389 ( .A(\mem<37><0> ), .B(n5016), .Y(n4522) );
  INVX1 U4390 ( .A(n4522), .Y(n4523) );
  AND2X2 U4391 ( .A(\mem<37><1> ), .B(n5017), .Y(n4524) );
  INVX1 U4392 ( .A(n4524), .Y(n4525) );
  AND2X2 U4393 ( .A(\mem<37><2> ), .B(n5016), .Y(n4526) );
  INVX1 U4394 ( .A(n4526), .Y(n4527) );
  AND2X2 U4395 ( .A(\mem<37><3> ), .B(n5017), .Y(n4528) );
  INVX1 U4396 ( .A(n4528), .Y(n4529) );
  AND2X2 U4397 ( .A(\mem<37><4> ), .B(n5016), .Y(n4530) );
  INVX1 U4398 ( .A(n4530), .Y(n4531) );
  AND2X2 U4399 ( .A(\mem<37><5> ), .B(n5017), .Y(n4532) );
  INVX1 U4400 ( .A(n4532), .Y(n4533) );
  AND2X2 U4401 ( .A(\mem<37><6> ), .B(n5016), .Y(n4534) );
  INVX1 U4402 ( .A(n4534), .Y(n4535) );
  AND2X2 U4403 ( .A(\mem<37><7> ), .B(n5017), .Y(n4536) );
  INVX1 U4404 ( .A(n4536), .Y(n4537) );
  AND2X2 U4405 ( .A(\mem<36><0> ), .B(n5018), .Y(n4538) );
  INVX1 U4406 ( .A(n4538), .Y(n4539) );
  AND2X2 U4407 ( .A(\mem<36><1> ), .B(n5019), .Y(n4540) );
  INVX1 U4408 ( .A(n4540), .Y(n4541) );
  AND2X2 U4409 ( .A(\mem<36><2> ), .B(n5018), .Y(n4542) );
  INVX1 U4410 ( .A(n4542), .Y(n4543) );
  AND2X2 U4411 ( .A(\mem<36><3> ), .B(n5019), .Y(n4544) );
  INVX1 U4412 ( .A(n4544), .Y(n4545) );
  AND2X2 U4413 ( .A(\mem<36><4> ), .B(n5018), .Y(n4546) );
  INVX1 U4414 ( .A(n4546), .Y(n4547) );
  AND2X2 U4415 ( .A(\mem<36><5> ), .B(n5019), .Y(n4548) );
  INVX1 U4416 ( .A(n4548), .Y(n4549) );
  AND2X2 U4417 ( .A(\mem<36><6> ), .B(n5018), .Y(n4550) );
  INVX1 U4418 ( .A(n4550), .Y(n4551) );
  AND2X2 U4419 ( .A(\mem<36><7> ), .B(n5019), .Y(n4552) );
  INVX1 U4420 ( .A(n4552), .Y(n4553) );
  AND2X2 U4421 ( .A(\mem<33><0> ), .B(n5024), .Y(n4554) );
  INVX1 U4422 ( .A(n4554), .Y(n4555) );
  AND2X2 U4423 ( .A(\mem<33><1> ), .B(n5025), .Y(n4556) );
  INVX1 U4424 ( .A(n4556), .Y(n4557) );
  AND2X2 U4425 ( .A(\mem<33><2> ), .B(n5024), .Y(n4558) );
  INVX1 U4426 ( .A(n4558), .Y(n4559) );
  AND2X2 U4427 ( .A(\mem<33><3> ), .B(n5025), .Y(n4560) );
  INVX1 U4428 ( .A(n4560), .Y(n4561) );
  AND2X2 U4429 ( .A(\mem<33><4> ), .B(n5024), .Y(n4562) );
  INVX1 U4430 ( .A(n4562), .Y(n4563) );
  AND2X2 U4431 ( .A(\mem<33><5> ), .B(n5025), .Y(n4564) );
  INVX1 U4432 ( .A(n4564), .Y(n4565) );
  AND2X2 U4433 ( .A(\mem<33><6> ), .B(n5024), .Y(n4566) );
  INVX1 U4434 ( .A(n4566), .Y(n4567) );
  AND2X2 U4435 ( .A(\mem<33><7> ), .B(n5025), .Y(n4568) );
  INVX1 U4436 ( .A(n4568), .Y(n4569) );
  AND2X2 U4437 ( .A(\mem<32><0> ), .B(n6426), .Y(n4570) );
  INVX1 U4438 ( .A(n4570), .Y(n4571) );
  AND2X2 U4439 ( .A(\mem<32><1> ), .B(n6426), .Y(n4572) );
  INVX1 U4440 ( .A(n4572), .Y(n4573) );
  AND2X2 U4441 ( .A(\mem<32><2> ), .B(n6426), .Y(n4574) );
  INVX1 U4442 ( .A(n4574), .Y(n4575) );
  AND2X2 U4443 ( .A(\mem<32><3> ), .B(n6426), .Y(n4576) );
  INVX1 U4444 ( .A(n4576), .Y(n4577) );
  AND2X2 U4445 ( .A(\mem<32><4> ), .B(n6426), .Y(n4578) );
  INVX1 U4446 ( .A(n4578), .Y(n4579) );
  AND2X2 U4447 ( .A(\mem<32><5> ), .B(n6426), .Y(n4580) );
  INVX1 U4448 ( .A(n4580), .Y(n4581) );
  AND2X2 U4449 ( .A(\mem<32><6> ), .B(n6426), .Y(n4582) );
  INVX1 U4450 ( .A(n4582), .Y(n4583) );
  AND2X2 U4451 ( .A(\mem<32><7> ), .B(n6426), .Y(n4584) );
  INVX1 U4452 ( .A(n4584), .Y(n4585) );
  AND2X2 U4453 ( .A(\mem<31><0> ), .B(n5026), .Y(n4586) );
  INVX1 U4454 ( .A(n4586), .Y(n4587) );
  AND2X2 U4455 ( .A(\mem<31><1> ), .B(n5027), .Y(n4588) );
  INVX1 U4456 ( .A(n4588), .Y(n4589) );
  AND2X2 U4457 ( .A(\mem<31><2> ), .B(n5026), .Y(n4590) );
  INVX1 U4458 ( .A(n4590), .Y(n4591) );
  AND2X2 U4459 ( .A(\mem<31><3> ), .B(n5027), .Y(n4592) );
  INVX1 U4460 ( .A(n4592), .Y(n4593) );
  AND2X2 U4461 ( .A(\mem<31><4> ), .B(n5027), .Y(n4594) );
  INVX1 U4462 ( .A(n4594), .Y(n4595) );
  AND2X2 U4463 ( .A(\mem<31><5> ), .B(n5026), .Y(n4596) );
  INVX1 U4464 ( .A(n4596), .Y(n4597) );
  AND2X2 U4465 ( .A(\mem<31><6> ), .B(n5026), .Y(n4598) );
  INVX1 U4466 ( .A(n4598), .Y(n4599) );
  AND2X2 U4467 ( .A(\mem<31><7> ), .B(n5027), .Y(n4600) );
  INVX1 U4468 ( .A(n4600), .Y(n4601) );
  AND2X2 U4469 ( .A(\mem<30><0> ), .B(n827), .Y(n4602) );
  INVX1 U4470 ( .A(n4602), .Y(n4603) );
  AND2X2 U4471 ( .A(\mem<30><1> ), .B(n827), .Y(n4604) );
  INVX1 U4472 ( .A(n4604), .Y(n4605) );
  AND2X2 U4473 ( .A(\mem<30><2> ), .B(n827), .Y(n4606) );
  INVX1 U4474 ( .A(n4606), .Y(n4607) );
  AND2X2 U4475 ( .A(\mem<30><3> ), .B(n827), .Y(n4608) );
  INVX1 U4476 ( .A(n4608), .Y(n4609) );
  AND2X2 U4477 ( .A(\mem<30><4> ), .B(n827), .Y(n4610) );
  INVX1 U4478 ( .A(n4610), .Y(n4611) );
  AND2X2 U4479 ( .A(\mem<30><5> ), .B(n827), .Y(n4612) );
  INVX1 U4480 ( .A(n4612), .Y(n4613) );
  AND2X2 U4481 ( .A(\mem<30><6> ), .B(n827), .Y(n4614) );
  INVX1 U4482 ( .A(n4614), .Y(n4615) );
  AND2X2 U4483 ( .A(\mem<30><7> ), .B(n827), .Y(n4616) );
  INVX1 U4484 ( .A(n4616), .Y(n4617) );
  AND2X2 U4485 ( .A(\mem<29><0> ), .B(n5028), .Y(n4618) );
  INVX1 U4486 ( .A(n4618), .Y(n4619) );
  AND2X2 U4487 ( .A(\mem<29><1> ), .B(n5029), .Y(n4620) );
  INVX1 U4488 ( .A(n4620), .Y(n4621) );
  AND2X2 U4489 ( .A(\mem<29><2> ), .B(n5028), .Y(n4622) );
  INVX1 U4490 ( .A(n4622), .Y(n4623) );
  AND2X2 U4491 ( .A(\mem<29><3> ), .B(n5029), .Y(n4624) );
  INVX1 U4492 ( .A(n4624), .Y(n4625) );
  AND2X2 U4493 ( .A(\mem<29><4> ), .B(n5028), .Y(n4626) );
  INVX1 U4494 ( .A(n4626), .Y(n4627) );
  AND2X2 U4495 ( .A(\mem<29><5> ), .B(n5029), .Y(n4628) );
  INVX1 U4496 ( .A(n4628), .Y(n4629) );
  AND2X2 U4497 ( .A(\mem<29><6> ), .B(n5028), .Y(n4630) );
  INVX1 U4498 ( .A(n4630), .Y(n4631) );
  AND2X2 U4499 ( .A(\mem<29><7> ), .B(n5029), .Y(n4632) );
  INVX1 U4500 ( .A(n4632), .Y(n4633) );
  AND2X2 U4501 ( .A(\mem<28><0> ), .B(n5031), .Y(n4634) );
  INVX1 U4502 ( .A(n4634), .Y(n4635) );
  AND2X2 U4503 ( .A(\mem<28><1> ), .B(n5031), .Y(n4636) );
  INVX1 U4504 ( .A(n4636), .Y(n4637) );
  AND2X2 U4505 ( .A(\mem<28><2> ), .B(n5030), .Y(n4638) );
  INVX1 U4506 ( .A(n4638), .Y(n4639) );
  AND2X2 U4507 ( .A(\mem<28><3> ), .B(n5030), .Y(n4640) );
  INVX1 U4508 ( .A(n4640), .Y(n4641) );
  AND2X2 U4509 ( .A(\mem<28><4> ), .B(n5030), .Y(n4642) );
  INVX1 U4510 ( .A(n4642), .Y(n4643) );
  AND2X2 U4511 ( .A(\mem<28><5> ), .B(n5031), .Y(n4644) );
  INVX1 U4512 ( .A(n4644), .Y(n4645) );
  AND2X2 U4513 ( .A(\mem<28><6> ), .B(n5031), .Y(n4646) );
  INVX1 U4514 ( .A(n4646), .Y(n4647) );
  AND2X2 U4515 ( .A(\mem<28><7> ), .B(n5030), .Y(n4648) );
  INVX1 U4516 ( .A(n4648), .Y(n4649) );
  AND2X2 U4517 ( .A(\mem<27><0> ), .B(n5032), .Y(n4650) );
  INVX1 U4518 ( .A(n4650), .Y(n4651) );
  AND2X2 U4519 ( .A(\mem<27><1> ), .B(n5032), .Y(n4652) );
  INVX1 U4520 ( .A(n4652), .Y(n4653) );
  AND2X2 U4521 ( .A(\mem<27><2> ), .B(n5032), .Y(n4654) );
  INVX1 U4522 ( .A(n4654), .Y(n4655) );
  AND2X2 U4523 ( .A(\mem<27><3> ), .B(n5032), .Y(n4656) );
  INVX1 U4524 ( .A(n4656), .Y(n4657) );
  AND2X2 U4525 ( .A(\mem<27><4> ), .B(n5032), .Y(n4658) );
  INVX1 U4526 ( .A(n4658), .Y(n4659) );
  AND2X2 U4527 ( .A(\mem<27><5> ), .B(n5032), .Y(n4660) );
  INVX1 U4528 ( .A(n4660), .Y(n4661) );
  AND2X2 U4529 ( .A(\mem<27><6> ), .B(n5032), .Y(n4662) );
  INVX1 U4530 ( .A(n4662), .Y(n4663) );
  AND2X2 U4531 ( .A(\mem<27><7> ), .B(n5032), .Y(n4664) );
  INVX1 U4532 ( .A(n4664), .Y(n4665) );
  AND2X2 U4533 ( .A(\mem<26><0> ), .B(n5033), .Y(n4666) );
  INVX1 U4534 ( .A(n4666), .Y(n4667) );
  AND2X2 U4535 ( .A(\mem<26><1> ), .B(n5034), .Y(n4668) );
  INVX1 U4536 ( .A(n4668), .Y(n4669) );
  AND2X2 U4537 ( .A(\mem<26><2> ), .B(n5033), .Y(n4670) );
  INVX1 U4538 ( .A(n4670), .Y(n4671) );
  AND2X2 U4539 ( .A(\mem<26><3> ), .B(n5034), .Y(n4672) );
  INVX1 U4540 ( .A(n4672), .Y(n4673) );
  AND2X2 U4541 ( .A(\mem<26><4> ), .B(n5033), .Y(n4674) );
  INVX1 U4542 ( .A(n4674), .Y(n4675) );
  AND2X2 U4543 ( .A(\mem<26><5> ), .B(n5034), .Y(n4676) );
  INVX1 U4544 ( .A(n4676), .Y(n4677) );
  AND2X2 U4545 ( .A(\mem<26><6> ), .B(n5033), .Y(n4678) );
  INVX1 U4546 ( .A(n4678), .Y(n4679) );
  AND2X2 U4547 ( .A(\mem<26><7> ), .B(n5034), .Y(n4680) );
  INVX1 U4548 ( .A(n4680), .Y(n4681) );
  AND2X2 U4549 ( .A(\mem<25><0> ), .B(n5035), .Y(n4682) );
  INVX1 U4550 ( .A(n4682), .Y(n4683) );
  AND2X2 U4551 ( .A(\mem<25><1> ), .B(n5035), .Y(n4684) );
  INVX1 U4552 ( .A(n4684), .Y(n4685) );
  AND2X2 U4553 ( .A(\mem<25><2> ), .B(n5035), .Y(n4686) );
  INVX1 U4554 ( .A(n4686), .Y(n4687) );
  AND2X2 U4555 ( .A(\mem<25><3> ), .B(n5035), .Y(n4688) );
  INVX1 U4556 ( .A(n4688), .Y(n4689) );
  AND2X2 U4557 ( .A(\mem<25><4> ), .B(n5035), .Y(n4690) );
  INVX1 U4558 ( .A(n4690), .Y(n4691) );
  AND2X2 U4559 ( .A(\mem<25><5> ), .B(n5035), .Y(n4692) );
  INVX1 U4560 ( .A(n4692), .Y(n4693) );
  AND2X2 U4561 ( .A(\mem<25><6> ), .B(n5035), .Y(n4694) );
  INVX1 U4562 ( .A(n4694), .Y(n4695) );
  AND2X2 U4563 ( .A(\mem<25><7> ), .B(n5035), .Y(n4696) );
  INVX1 U4564 ( .A(n4696), .Y(n4697) );
  AND2X2 U4565 ( .A(\mem<24><0> ), .B(n5036), .Y(n4698) );
  INVX1 U4566 ( .A(n4698), .Y(n4699) );
  AND2X2 U4567 ( .A(\mem<24><1> ), .B(n5037), .Y(n4700) );
  INVX1 U4568 ( .A(n4700), .Y(n4701) );
  AND2X2 U4569 ( .A(\mem<24><2> ), .B(n74), .Y(n4702) );
  INVX1 U4570 ( .A(n4702), .Y(n4703) );
  AND2X2 U4571 ( .A(\mem<24><3> ), .B(n5036), .Y(n4704) );
  INVX1 U4572 ( .A(n4704), .Y(n4705) );
  AND2X2 U4573 ( .A(\mem<24><4> ), .B(n5037), .Y(n4706) );
  INVX1 U4574 ( .A(n4706), .Y(n4707) );
  AND2X2 U4575 ( .A(\mem<24><5> ), .B(n74), .Y(n4708) );
  INVX1 U4576 ( .A(n4708), .Y(n4709) );
  AND2X2 U4577 ( .A(\mem<24><6> ), .B(n5036), .Y(n4710) );
  INVX1 U4578 ( .A(n4710), .Y(n4711) );
  AND2X2 U4579 ( .A(\mem<24><7> ), .B(n5037), .Y(n4712) );
  INVX1 U4580 ( .A(n4712), .Y(n4713) );
  AND2X2 U4581 ( .A(\mem<23><0> ), .B(n5038), .Y(n4714) );
  INVX1 U4582 ( .A(n4714), .Y(n4715) );
  AND2X2 U4583 ( .A(\mem<23><1> ), .B(n5039), .Y(n4716) );
  INVX1 U4584 ( .A(n4716), .Y(n4717) );
  AND2X2 U4585 ( .A(\mem<23><2> ), .B(n5038), .Y(n4718) );
  INVX1 U4586 ( .A(n4718), .Y(n4719) );
  AND2X2 U4587 ( .A(\mem<23><3> ), .B(n5039), .Y(n4720) );
  INVX1 U4588 ( .A(n4720), .Y(n4721) );
  AND2X2 U4589 ( .A(\mem<23><4> ), .B(n5038), .Y(n4722) );
  INVX1 U4590 ( .A(n4722), .Y(n4723) );
  AND2X2 U4591 ( .A(\mem<23><5> ), .B(n5039), .Y(n4724) );
  INVX1 U4592 ( .A(n4724), .Y(n4725) );
  AND2X2 U4593 ( .A(\mem<23><6> ), .B(n5038), .Y(n4726) );
  INVX1 U4594 ( .A(n4726), .Y(n4727) );
  AND2X2 U4595 ( .A(\mem<23><7> ), .B(n5039), .Y(n4728) );
  INVX1 U4596 ( .A(n4728), .Y(n4729) );
  AND2X2 U4597 ( .A(\mem<22><0> ), .B(n5040), .Y(n4730) );
  INVX1 U4598 ( .A(n4730), .Y(n4731) );
  AND2X2 U4599 ( .A(\mem<22><1> ), .B(n5041), .Y(n4732) );
  INVX1 U4600 ( .A(n4732), .Y(n4733) );
  AND2X2 U4601 ( .A(\mem<22><2> ), .B(n5040), .Y(n4734) );
  INVX1 U4602 ( .A(n4734), .Y(n4735) );
  AND2X2 U4603 ( .A(\mem<22><3> ), .B(n5041), .Y(n4736) );
  INVX1 U4604 ( .A(n4736), .Y(n4737) );
  AND2X2 U4605 ( .A(\mem<22><4> ), .B(n5040), .Y(n4738) );
  INVX1 U4606 ( .A(n4738), .Y(n4739) );
  AND2X2 U4607 ( .A(\mem<22><5> ), .B(n5041), .Y(n4740) );
  INVX1 U4608 ( .A(n4740), .Y(n4741) );
  AND2X2 U4609 ( .A(\mem<22><6> ), .B(n5040), .Y(n4742) );
  INVX1 U4610 ( .A(n4742), .Y(n4743) );
  AND2X2 U4611 ( .A(\mem<22><7> ), .B(n5041), .Y(n4744) );
  INVX1 U4612 ( .A(n4744), .Y(n4745) );
  AND2X2 U4613 ( .A(\mem<21><0> ), .B(n5042), .Y(n4746) );
  INVX1 U4614 ( .A(n4746), .Y(n4747) );
  AND2X2 U4615 ( .A(\mem<21><1> ), .B(n5043), .Y(n4748) );
  INVX1 U4616 ( .A(n4748), .Y(n4749) );
  AND2X2 U4617 ( .A(\mem<21><2> ), .B(n5042), .Y(n4750) );
  INVX1 U4618 ( .A(n4750), .Y(n4751) );
  AND2X2 U4619 ( .A(\mem<21><3> ), .B(n5043), .Y(n4752) );
  INVX1 U4620 ( .A(n4752), .Y(n4753) );
  AND2X2 U4621 ( .A(\mem<21><4> ), .B(n5042), .Y(n4754) );
  INVX1 U4622 ( .A(n4754), .Y(n4755) );
  AND2X2 U4623 ( .A(\mem<21><5> ), .B(n5043), .Y(n4756) );
  INVX1 U4624 ( .A(n4756), .Y(n4757) );
  AND2X2 U4625 ( .A(\mem<21><6> ), .B(n5042), .Y(n4758) );
  INVX1 U4626 ( .A(n4758), .Y(n4759) );
  AND2X2 U4627 ( .A(\mem<21><7> ), .B(n5043), .Y(n4760) );
  INVX1 U4628 ( .A(n4760), .Y(n4761) );
  AND2X2 U4629 ( .A(\mem<20><0> ), .B(n5045), .Y(n4762) );
  INVX1 U4630 ( .A(n4762), .Y(n4763) );
  AND2X2 U4631 ( .A(\mem<20><1> ), .B(n5044), .Y(n4764) );
  INVX1 U4632 ( .A(n4764), .Y(n4765) );
  AND2X2 U4633 ( .A(\mem<20><2> ), .B(n5045), .Y(n4766) );
  INVX1 U4634 ( .A(n4766), .Y(n4767) );
  AND2X2 U4635 ( .A(\mem<20><3> ), .B(n5044), .Y(n4768) );
  INVX1 U4636 ( .A(n4768), .Y(n4769) );
  AND2X2 U4637 ( .A(\mem<20><4> ), .B(n5045), .Y(n4770) );
  INVX1 U4638 ( .A(n4770), .Y(n4771) );
  AND2X2 U4639 ( .A(\mem<20><5> ), .B(n5044), .Y(n4772) );
  INVX1 U4640 ( .A(n4772), .Y(n4773) );
  AND2X2 U4641 ( .A(\mem<20><6> ), .B(n5045), .Y(n4774) );
  INVX1 U4642 ( .A(n4774), .Y(n4775) );
  AND2X2 U4643 ( .A(\mem<20><7> ), .B(n5044), .Y(n4776) );
  INVX1 U4644 ( .A(n4776), .Y(n4777) );
  AND2X2 U4645 ( .A(\mem<19><0> ), .B(n5046), .Y(n4778) );
  INVX1 U4646 ( .A(n4778), .Y(n4779) );
  AND2X2 U4647 ( .A(\mem<19><1> ), .B(n5047), .Y(n4780) );
  INVX1 U4648 ( .A(n4780), .Y(n4781) );
  AND2X2 U4649 ( .A(\mem<19><2> ), .B(n57), .Y(n4782) );
  INVX1 U4650 ( .A(n4782), .Y(n4783) );
  AND2X2 U4651 ( .A(\mem<19><3> ), .B(n5046), .Y(n4784) );
  INVX1 U4652 ( .A(n4784), .Y(n4785) );
  AND2X2 U4653 ( .A(\mem<19><4> ), .B(n5047), .Y(n4786) );
  INVX1 U4654 ( .A(n4786), .Y(n4787) );
  AND2X2 U4655 ( .A(\mem<19><5> ), .B(n57), .Y(n4788) );
  INVX1 U4656 ( .A(n4788), .Y(n4789) );
  AND2X2 U4657 ( .A(\mem<19><6> ), .B(n5046), .Y(n4790) );
  INVX1 U4658 ( .A(n4790), .Y(n4791) );
  AND2X2 U4659 ( .A(\mem<19><7> ), .B(n5047), .Y(n4792) );
  INVX1 U4660 ( .A(n4792), .Y(n4793) );
  AND2X2 U4661 ( .A(\mem<18><0> ), .B(n5049), .Y(n4794) );
  INVX1 U4662 ( .A(n4794), .Y(n4795) );
  AND2X2 U4663 ( .A(\mem<18><1> ), .B(n5048), .Y(n4796) );
  INVX1 U4664 ( .A(n4796), .Y(n4797) );
  AND2X2 U4665 ( .A(\mem<18><2> ), .B(n5048), .Y(n4798) );
  INVX1 U4666 ( .A(n4798), .Y(n4799) );
  AND2X2 U4667 ( .A(\mem<18><3> ), .B(n5048), .Y(n4800) );
  INVX1 U4668 ( .A(n4800), .Y(n4801) );
  AND2X2 U4669 ( .A(\mem<18><4> ), .B(n5048), .Y(n4802) );
  INVX1 U4670 ( .A(n4802), .Y(n4803) );
  AND2X2 U4671 ( .A(\mem<18><5> ), .B(n5049), .Y(n4804) );
  INVX1 U4672 ( .A(n4804), .Y(n4805) );
  AND2X2 U4673 ( .A(\mem<18><6> ), .B(n5049), .Y(n4806) );
  INVX1 U4674 ( .A(n4806), .Y(n4807) );
  AND2X2 U4675 ( .A(\mem<18><7> ), .B(n5049), .Y(n4808) );
  INVX1 U4676 ( .A(n4808), .Y(n4809) );
  AND2X2 U4677 ( .A(\mem<17><0> ), .B(n5050), .Y(n4810) );
  INVX1 U4678 ( .A(n4810), .Y(n4811) );
  AND2X2 U4679 ( .A(\mem<17><1> ), .B(n5051), .Y(n4812) );
  INVX1 U4680 ( .A(n4812), .Y(n4813) );
  AND2X2 U4681 ( .A(\mem<17><2> ), .B(n5050), .Y(n4814) );
  INVX1 U4682 ( .A(n4814), .Y(n4815) );
  AND2X2 U4683 ( .A(\mem<17><3> ), .B(n5051), .Y(n4816) );
  INVX1 U4684 ( .A(n4816), .Y(n4817) );
  AND2X2 U4685 ( .A(\mem<17><4> ), .B(n5050), .Y(n4818) );
  INVX1 U4686 ( .A(n4818), .Y(n4819) );
  AND2X2 U4687 ( .A(\mem<17><5> ), .B(n5051), .Y(n4820) );
  INVX1 U4688 ( .A(n4820), .Y(n4821) );
  AND2X2 U4689 ( .A(\mem<17><6> ), .B(n5050), .Y(n4822) );
  INVX1 U4690 ( .A(n4822), .Y(n4823) );
  AND2X2 U4691 ( .A(\mem<17><7> ), .B(n5051), .Y(n4824) );
  INVX1 U4692 ( .A(n4824), .Y(n4825) );
  AND2X2 U4693 ( .A(\mem<15><0> ), .B(n5053), .Y(n4826) );
  INVX1 U4694 ( .A(n4826), .Y(n4827) );
  AND2X2 U4695 ( .A(\mem<15><1> ), .B(n5054), .Y(n4828) );
  INVX1 U4696 ( .A(n4828), .Y(n4829) );
  AND2X2 U4697 ( .A(\mem<15><2> ), .B(n5053), .Y(n4830) );
  INVX1 U4698 ( .A(n4830), .Y(n4831) );
  AND2X2 U4699 ( .A(\mem<15><3> ), .B(n5054), .Y(n4832) );
  INVX1 U4700 ( .A(n4832), .Y(n4833) );
  AND2X2 U4701 ( .A(\mem<15><4> ), .B(n5053), .Y(n4834) );
  INVX1 U4702 ( .A(n4834), .Y(n4835) );
  AND2X2 U4703 ( .A(\mem<15><5> ), .B(n5054), .Y(n4836) );
  INVX1 U4704 ( .A(n4836), .Y(n4837) );
  AND2X2 U4705 ( .A(\mem<15><6> ), .B(n5053), .Y(n4838) );
  INVX1 U4706 ( .A(n4838), .Y(n4839) );
  AND2X2 U4707 ( .A(\mem<15><7> ), .B(n5054), .Y(n4840) );
  INVX1 U4708 ( .A(n4840), .Y(n4841) );
  AND2X2 U4709 ( .A(\mem<14><0> ), .B(n4967), .Y(n4842) );
  INVX1 U4710 ( .A(n4842), .Y(n4843) );
  AND2X2 U4711 ( .A(\mem<14><1> ), .B(n4968), .Y(n4844) );
  INVX1 U4712 ( .A(n4844), .Y(n4845) );
  AND2X2 U4713 ( .A(\mem<14><2> ), .B(n4967), .Y(n4846) );
  INVX1 U4714 ( .A(n4846), .Y(n4847) );
  AND2X2 U4715 ( .A(\mem<14><3> ), .B(n4968), .Y(n4848) );
  INVX1 U4716 ( .A(n4848), .Y(n4849) );
  AND2X2 U4717 ( .A(\mem<14><4> ), .B(n4967), .Y(n4850) );
  INVX1 U4718 ( .A(n4850), .Y(n4851) );
  AND2X2 U4719 ( .A(\mem<14><5> ), .B(n4968), .Y(n4852) );
  INVX1 U4720 ( .A(n4852), .Y(n4853) );
  AND2X2 U4721 ( .A(\mem<14><6> ), .B(n4967), .Y(n4854) );
  INVX1 U4722 ( .A(n4854), .Y(n4855) );
  AND2X2 U4723 ( .A(\mem<14><7> ), .B(n4968), .Y(n4856) );
  INVX1 U4724 ( .A(n4856), .Y(n4857) );
  AND2X2 U4725 ( .A(\mem<7><0> ), .B(n5063), .Y(n4858) );
  INVX1 U4726 ( .A(n4858), .Y(n4859) );
  AND2X2 U4727 ( .A(\mem<7><1> ), .B(n5064), .Y(n4860) );
  INVX1 U4728 ( .A(n4860), .Y(n4861) );
  AND2X2 U4729 ( .A(\mem<7><2> ), .B(n5063), .Y(n4862) );
  INVX1 U4730 ( .A(n4862), .Y(n4863) );
  AND2X2 U4731 ( .A(\mem<7><3> ), .B(n5064), .Y(n4864) );
  INVX1 U4732 ( .A(n4864), .Y(n4865) );
  AND2X2 U4733 ( .A(\mem<7><4> ), .B(n5063), .Y(n4866) );
  INVX1 U4734 ( .A(n4866), .Y(n4867) );
  AND2X2 U4735 ( .A(\mem<7><5> ), .B(n5064), .Y(n4868) );
  INVX1 U4736 ( .A(n4868), .Y(n4869) );
  AND2X2 U4737 ( .A(\mem<7><6> ), .B(n5063), .Y(n4870) );
  INVX1 U4738 ( .A(n4870), .Y(n4871) );
  AND2X2 U4739 ( .A(\mem<7><7> ), .B(n5064), .Y(n4872) );
  INVX1 U4740 ( .A(n4872), .Y(n4873) );
  AND2X2 U4741 ( .A(\mem<6><0> ), .B(n898), .Y(n4874) );
  INVX1 U4742 ( .A(n4874), .Y(n4875) );
  AND2X2 U4743 ( .A(\mem<6><1> ), .B(n69), .Y(n4876) );
  INVX1 U4744 ( .A(n4876), .Y(n4877) );
  AND2X2 U4745 ( .A(\mem<6><2> ), .B(n69), .Y(n4878) );
  INVX1 U4746 ( .A(n4878), .Y(n4879) );
  AND2X2 U4747 ( .A(\mem<6><3> ), .B(n898), .Y(n4880) );
  INVX1 U4748 ( .A(n4880), .Y(n4881) );
  AND2X2 U4749 ( .A(\mem<6><4> ), .B(n69), .Y(n4882) );
  INVX1 U4750 ( .A(n4882), .Y(n4883) );
  AND2X2 U4751 ( .A(\mem<6><5> ), .B(n69), .Y(n4884) );
  INVX1 U4752 ( .A(n4884), .Y(n4885) );
  AND2X2 U4753 ( .A(\mem<6><6> ), .B(n898), .Y(n4886) );
  INVX1 U4754 ( .A(n4886), .Y(n4887) );
  AND2X2 U4755 ( .A(\mem<6><7> ), .B(n69), .Y(n4888) );
  INVX1 U4756 ( .A(n4888), .Y(n4889) );
  AND2X2 U4757 ( .A(\mem<4><0> ), .B(n5067), .Y(n4890) );
  INVX1 U4758 ( .A(n4890), .Y(n4891) );
  AND2X2 U4759 ( .A(\mem<4><1> ), .B(n5068), .Y(n4892) );
  INVX1 U4760 ( .A(n4892), .Y(n4893) );
  AND2X2 U4761 ( .A(\mem<4><2> ), .B(n5067), .Y(n4894) );
  INVX1 U4762 ( .A(n4894), .Y(n4895) );
  AND2X2 U4763 ( .A(\mem<4><3> ), .B(n5068), .Y(n4896) );
  INVX1 U4764 ( .A(n4896), .Y(n4897) );
  AND2X2 U4765 ( .A(\mem<4><4> ), .B(n5067), .Y(n4898) );
  INVX1 U4766 ( .A(n4898), .Y(n4899) );
  AND2X2 U4767 ( .A(\mem<4><5> ), .B(n5068), .Y(n4900) );
  INVX1 U4768 ( .A(n4900), .Y(n4901) );
  AND2X2 U4769 ( .A(\mem<4><6> ), .B(n5067), .Y(n4902) );
  INVX1 U4770 ( .A(n4902), .Y(n4903) );
  AND2X2 U4771 ( .A(\mem<4><7> ), .B(n5068), .Y(n4904) );
  INVX1 U4772 ( .A(n4904), .Y(n4905) );
  AND2X2 U4773 ( .A(\mem<3><0> ), .B(n5070), .Y(n4906) );
  INVX1 U4774 ( .A(n4906), .Y(n4907) );
  AND2X2 U4775 ( .A(\mem<3><1> ), .B(n5070), .Y(n4908) );
  INVX1 U4776 ( .A(n4908), .Y(n4909) );
  AND2X2 U4777 ( .A(\mem<3><2> ), .B(n5070), .Y(n4910) );
  INVX1 U4778 ( .A(n4910), .Y(n4911) );
  AND2X2 U4779 ( .A(\mem<3><3> ), .B(n5069), .Y(n4912) );
  INVX1 U4780 ( .A(n4912), .Y(n4913) );
  AND2X2 U4781 ( .A(\mem<3><4> ), .B(n5069), .Y(n4914) );
  INVX1 U4782 ( .A(n4914), .Y(n4915) );
  AND2X2 U4783 ( .A(\mem<3><5> ), .B(n5069), .Y(n4916) );
  INVX1 U4784 ( .A(n4916), .Y(n4917) );
  AND2X2 U4785 ( .A(\mem<3><6> ), .B(n5070), .Y(n4918) );
  INVX1 U4786 ( .A(n4918), .Y(n4919) );
  AND2X2 U4787 ( .A(\mem<3><7> ), .B(n5069), .Y(n4920) );
  INVX1 U4788 ( .A(n4920), .Y(n4921) );
  AND2X2 U4789 ( .A(\mem<2><0> ), .B(n5071), .Y(n4922) );
  INVX1 U4790 ( .A(n4922), .Y(n4923) );
  AND2X2 U4791 ( .A(\mem<2><1> ), .B(n5072), .Y(n4924) );
  INVX1 U4792 ( .A(n4924), .Y(n4925) );
  AND2X2 U4793 ( .A(\mem<2><2> ), .B(n5071), .Y(n4926) );
  INVX1 U4794 ( .A(n4926), .Y(n4927) );
  AND2X2 U4795 ( .A(\mem<2><3> ), .B(n5072), .Y(n4928) );
  INVX1 U4796 ( .A(n4928), .Y(n4929) );
  AND2X2 U4797 ( .A(\mem<2><4> ), .B(n5071), .Y(n4930) );
  INVX1 U4798 ( .A(n4930), .Y(n4931) );
  AND2X2 U4799 ( .A(\mem<2><5> ), .B(n5072), .Y(n4932) );
  INVX1 U4800 ( .A(n4932), .Y(n4933) );
  AND2X2 U4801 ( .A(\mem<2><6> ), .B(n5071), .Y(n4934) );
  INVX1 U4802 ( .A(n4934), .Y(n4935) );
  AND2X2 U4803 ( .A(\mem<2><7> ), .B(n5072), .Y(n4936) );
  INVX1 U4804 ( .A(n4936), .Y(n4937) );
  INVX2 U4805 ( .A(n3909), .Y(n5753) );
  AND2X2 U4806 ( .A(n78), .B(n591), .Y(n4938) );
  AND2X2 U4807 ( .A(n5726), .B(n5194), .Y(n4939) );
  INVX1 U4808 ( .A(n4939), .Y(n4940) );
  AND2X2 U4809 ( .A(N182), .B(n5193), .Y(n4941) );
  INVX1 U4810 ( .A(n4941), .Y(n4942) );
  INVX1 U4811 ( .A(n4941), .Y(n4943) );
  INVX1 U4812 ( .A(wr), .Y(n5856) );
  INVX1 U4813 ( .A(n3686), .Y(n4944) );
  INVX1 U4814 ( .A(n3686), .Y(n4945) );
  INVX1 U4815 ( .A(n557), .Y(n4946) );
  INVX1 U4816 ( .A(n557), .Y(n4947) );
  INVX1 U4817 ( .A(n6438), .Y(n4948) );
  INVX1 U4818 ( .A(n4948), .Y(n4950) );
  INVX1 U4819 ( .A(n6449), .Y(n4951) );
  INVX1 U4820 ( .A(n4951), .Y(n4952) );
  INVX1 U4821 ( .A(n4951), .Y(n4953) );
  INVX1 U4822 ( .A(n4951), .Y(n4954) );
  INVX1 U4823 ( .A(n6451), .Y(n4955) );
  INVX2 U4824 ( .A(n4955), .Y(n4956) );
  INVX1 U4825 ( .A(n6450), .Y(n4957) );
  INVX1 U4826 ( .A(n4957), .Y(n4958) );
  INVX1 U4827 ( .A(n4957), .Y(n4959) );
  INVX1 U4828 ( .A(n4957), .Y(n4960) );
  INVX1 U4829 ( .A(n6452), .Y(n4961) );
  INVX2 U4830 ( .A(n4961), .Y(n4962) );
  INVX1 U4831 ( .A(n6453), .Y(n4963) );
  INVX1 U4832 ( .A(n6455), .Y(n4965) );
  INVX2 U4833 ( .A(n4965), .Y(n4966) );
  INVX1 U4834 ( .A(n563), .Y(n4967) );
  INVX1 U4835 ( .A(n563), .Y(n4968) );
  INVX1 U4836 ( .A(n666), .Y(n4969) );
  INVX1 U4837 ( .A(n666), .Y(n4970) );
  INVX1 U4838 ( .A(n667), .Y(n4971) );
  INVX1 U4839 ( .A(n667), .Y(n4972) );
  INVX1 U4840 ( .A(n668), .Y(n4973) );
  INVX1 U4841 ( .A(n668), .Y(n4974) );
  INVX1 U4842 ( .A(n669), .Y(n4975) );
  INVX1 U4843 ( .A(n669), .Y(n4976) );
  INVX1 U4844 ( .A(n670), .Y(n4977) );
  INVX1 U4845 ( .A(n670), .Y(n4978) );
  INVX1 U4846 ( .A(n671), .Y(n4979) );
  INVX1 U4847 ( .A(n671), .Y(n4980) );
  INVX1 U4848 ( .A(n672), .Y(n4981) );
  INVX1 U4849 ( .A(n672), .Y(n4982) );
  INVX1 U4850 ( .A(n674), .Y(n4983) );
  INVX1 U4851 ( .A(n4983), .Y(n4984) );
  INVX1 U4852 ( .A(n4983), .Y(n4985) );
  INVX1 U4853 ( .A(n675), .Y(n4986) );
  INVX1 U4854 ( .A(n675), .Y(n4987) );
  INVX1 U4855 ( .A(n676), .Y(n4988) );
  INVX1 U4856 ( .A(n676), .Y(n4989) );
  INVX1 U4857 ( .A(n677), .Y(n4990) );
  INVX1 U4858 ( .A(n677), .Y(n4991) );
  INVX1 U4859 ( .A(n678), .Y(n4992) );
  INVX1 U4860 ( .A(n678), .Y(n4993) );
  INVX1 U4861 ( .A(n692), .Y(n4994) );
  INVX1 U4862 ( .A(n692), .Y(n4995) );
  INVX1 U4863 ( .A(n693), .Y(n4996) );
  INVX1 U4864 ( .A(n693), .Y(n4997) );
  INVX1 U4865 ( .A(n696), .Y(n4998) );
  INVX1 U4866 ( .A(n696), .Y(n4999) );
  INVX1 U4867 ( .A(n713), .Y(n5000) );
  INVX1 U4868 ( .A(n713), .Y(n5001) );
  INVX1 U4869 ( .A(n728), .Y(n5002) );
  INVX1 U4870 ( .A(n728), .Y(n5003) );
  INVX1 U4871 ( .A(n740), .Y(n5004) );
  INVX1 U4872 ( .A(n740), .Y(n5005) );
  INVX1 U4873 ( .A(n752), .Y(n5006) );
  INVX1 U4874 ( .A(n752), .Y(n5007) );
  INVX1 U4875 ( .A(n765), .Y(n5008) );
  INVX1 U4876 ( .A(n777), .Y(n5010) );
  INVX1 U4877 ( .A(n777), .Y(n5011) );
  INVX1 U4878 ( .A(n782), .Y(n5012) );
  INVX1 U4879 ( .A(n783), .Y(n5013) );
  INVX1 U4880 ( .A(n808), .Y(n5014) );
  INVX1 U4881 ( .A(n808), .Y(n5015) );
  INVX1 U4882 ( .A(n809), .Y(n5016) );
  INVX1 U4883 ( .A(n809), .Y(n5017) );
  INVX1 U4884 ( .A(n810), .Y(n5018) );
  INVX1 U4885 ( .A(n810), .Y(n5019) );
  INVX1 U4886 ( .A(n811), .Y(n5020) );
  INVX1 U4887 ( .A(n811), .Y(n5021) );
  INVX1 U4888 ( .A(n812), .Y(n5022) );
  INVX1 U4889 ( .A(n812), .Y(n5023) );
  INVX1 U4890 ( .A(n824), .Y(n5024) );
  INVX1 U4891 ( .A(n824), .Y(n5025) );
  INVX1 U4892 ( .A(n825), .Y(n5026) );
  INVX1 U4893 ( .A(n825), .Y(n5027) );
  INVX1 U4894 ( .A(n828), .Y(n5028) );
  INVX1 U4895 ( .A(n828), .Y(n5029) );
  INVX1 U4896 ( .A(n829), .Y(n5030) );
  INVX1 U4897 ( .A(n829), .Y(n5031) );
  INVX1 U4898 ( .A(n830), .Y(n5032) );
  INVX1 U4899 ( .A(n831), .Y(n5033) );
  INVX1 U4900 ( .A(n831), .Y(n5034) );
  INVX1 U4901 ( .A(n832), .Y(n5035) );
  INVX1 U4902 ( .A(n833), .Y(n5036) );
  INVX1 U4903 ( .A(n833), .Y(n5037) );
  INVX1 U4904 ( .A(n834), .Y(n5038) );
  INVX1 U4905 ( .A(n834), .Y(n5039) );
  INVX1 U4906 ( .A(n835), .Y(n5040) );
  INVX1 U4907 ( .A(n835), .Y(n5041) );
  INVX1 U4908 ( .A(n836), .Y(n5042) );
  INVX1 U4909 ( .A(n836), .Y(n5043) );
  INVX1 U4910 ( .A(n837), .Y(n5044) );
  INVX1 U4911 ( .A(n837), .Y(n5045) );
  INVX1 U4912 ( .A(n869), .Y(n5046) );
  INVX1 U4913 ( .A(n869), .Y(n5047) );
  INVX1 U4914 ( .A(n870), .Y(n5048) );
  INVX1 U4915 ( .A(n870), .Y(n5049) );
  INVX1 U4916 ( .A(n871), .Y(n5050) );
  INVX1 U4917 ( .A(n871), .Y(n5051) );
  INVX1 U4918 ( .A(n873), .Y(n5053) );
  INVX1 U4919 ( .A(n873), .Y(n5054) );
  INVX1 U4920 ( .A(n874), .Y(n5055) );
  INVX1 U4921 ( .A(n874), .Y(n5056) );
  INVX1 U4922 ( .A(n875), .Y(n5057) );
  INVX1 U4923 ( .A(n875), .Y(n5058) );
  INVX1 U4924 ( .A(n876), .Y(n5059) );
  INVX1 U4925 ( .A(n877), .Y(n5060) );
  INVX1 U4926 ( .A(n878), .Y(n5061) );
  INVX1 U4927 ( .A(n878), .Y(n5062) );
  INVX1 U4928 ( .A(n896), .Y(n5063) );
  INVX1 U4929 ( .A(n896), .Y(n5064) );
  INVX1 U4930 ( .A(n899), .Y(n5065) );
  INVX1 U4931 ( .A(n899), .Y(n5066) );
  INVX1 U4932 ( .A(n900), .Y(n5067) );
  INVX1 U4933 ( .A(n900), .Y(n5068) );
  INVX1 U4934 ( .A(n901), .Y(n5069) );
  INVX1 U4935 ( .A(n901), .Y(n5070) );
  INVX1 U4936 ( .A(n902), .Y(n5071) );
  INVX1 U4937 ( .A(n902), .Y(n5072) );
  INVX1 U4938 ( .A(n5593), .Y(n5073) );
  INVX1 U4939 ( .A(n5273), .Y(n5074) );
  AOI22X1 U4940 ( .A(n5705), .B(\mem<6><3> ), .C(\mem<4><3> ), .D(n149), .Y(
        n5075) );
  INVX2 U4941 ( .A(n5075), .Y(n6070) );
  AND2X2 U4942 ( .A(n6425), .B(n6457), .Y(n5076) );
  OAI21X1 U4943 ( .A(n3909), .B(n5921), .C(n5920), .Y(n5925) );
  INVX1 U4944 ( .A(\mem<1><1> ), .Y(n5921) );
  NAND3X1 U4945 ( .A(n3766), .B(n597), .C(n553), .Y(n5077) );
  INVX1 U4946 ( .A(n5077), .Y(n6088) );
  INVX1 U4947 ( .A(n5246), .Y(n5078) );
  INVX1 U4948 ( .A(n5536), .Y(n5079) );
  INVX1 U4949 ( .A(n5707), .Y(n5080) );
  INVX1 U4950 ( .A(n5492), .Y(n5081) );
  INVX1 U4951 ( .A(n5157), .Y(n5082) );
  INVX1 U4952 ( .A(n5507), .Y(n5083) );
  INVX1 U4953 ( .A(N181), .Y(n5084) );
  INVX1 U4954 ( .A(n5259), .Y(n5085) );
  AND2X2 U4955 ( .A(n5742), .B(n874), .Y(n6437) );
  NAND3X1 U4956 ( .A(n4015), .B(n2890), .C(n3600), .Y(n6574) );
  NAND3X1 U4957 ( .A(n4013), .B(n2888), .C(n3598), .Y(n6575) );
  NAND3X1 U4958 ( .A(n4011), .B(n2886), .C(n3596), .Y(n6576) );
  NAND3X1 U4959 ( .A(n4009), .B(n2884), .C(n3594), .Y(n6577) );
  NAND3X1 U4960 ( .A(n4007), .B(n2882), .C(n3592), .Y(n6578) );
  NAND3X1 U4961 ( .A(n4005), .B(n2880), .C(n3590), .Y(n6579) );
  NAND3X1 U4962 ( .A(n4003), .B(n2878), .C(n3588), .Y(n6580) );
  NAND3X1 U4963 ( .A(n4001), .B(n2876), .C(n3586), .Y(n6581) );
  NAND3X1 U4964 ( .A(n3842), .B(n2938), .C(n3636), .Y(n6550) );
  NAND3X1 U4965 ( .A(n3840), .B(n2936), .C(n3634), .Y(n6551) );
  NAND3X1 U4966 ( .A(n4035), .B(n2934), .C(n3632), .Y(n6552) );
  NAND3X1 U4967 ( .A(n3838), .B(n2932), .C(n3630), .Y(n6553) );
  NAND3X1 U4968 ( .A(n3836), .B(n2930), .C(n3628), .Y(n6554) );
  NAND3X1 U4969 ( .A(n4033), .B(n2928), .C(n3626), .Y(n6555) );
  NAND3X1 U4970 ( .A(n3834), .B(n2926), .C(n3624), .Y(n6556) );
  NAND3X1 U4971 ( .A(n3832), .B(n2924), .C(n3622), .Y(n6557) );
  NAND3X1 U4972 ( .A(n4031), .B(n2906), .C(n3616), .Y(n6566) );
  NAND3X1 U4973 ( .A(n4029), .B(n2904), .C(n3614), .Y(n6567) );
  NAND3X1 U4974 ( .A(n4027), .B(n2902), .C(n3612), .Y(n6568) );
  NAND3X1 U4975 ( .A(n4025), .B(n2900), .C(n3610), .Y(n6569) );
  NAND3X1 U4976 ( .A(n4023), .B(n2898), .C(n3608), .Y(n6570) );
  NAND3X1 U4977 ( .A(n4021), .B(n2896), .C(n3606), .Y(n6571) );
  NAND3X1 U4978 ( .A(n4019), .B(n2894), .C(n3604), .Y(n6572) );
  NAND3X1 U4979 ( .A(n4017), .B(n2892), .C(n3602), .Y(n6573) );
  NAND3X1 U4980 ( .A(n3830), .B(n2874), .C(n3584), .Y(n6582) );
  NAND3X1 U4981 ( .A(n3828), .B(n2872), .C(n3582), .Y(n6583) );
  NAND3X1 U4982 ( .A(n3826), .B(n2870), .C(n3580), .Y(n6584) );
  NAND3X1 U4983 ( .A(n3824), .B(n2868), .C(n3578), .Y(n6585) );
  NAND3X1 U4984 ( .A(n3822), .B(n2866), .C(n3576), .Y(n6586) );
  NAND3X1 U4985 ( .A(n3820), .B(n2864), .C(n3574), .Y(n6587) );
  NAND3X1 U4986 ( .A(n3818), .B(n2862), .C(n3572), .Y(n6588) );
  NAND3X1 U4987 ( .A(n3816), .B(n2860), .C(n3570), .Y(n6589) );
  INVX1 U4988 ( .A(N181), .Y(n5086) );
  INVX1 U4989 ( .A(n5579), .Y(n5087) );
  INVX1 U4990 ( .A(n5565), .Y(n5088) );
  INVX1 U4991 ( .A(n3657), .Y(n6422) );
  INVX1 U4992 ( .A(n5711), .Y(n5089) );
  INVX1 U4993 ( .A(n5551), .Y(n5090) );
  INVX1 U4994 ( .A(N181), .Y(n5091) );
  NAND3X1 U4995 ( .A(n1149), .B(n5092), .C(n1706), .Y(n5093) );
  INVX1 U4996 ( .A(n6375), .Y(n5092) );
  INVX1 U4997 ( .A(n5093), .Y(n6398) );
  NAND3X1 U4998 ( .A(n1705), .B(n5094), .C(n1148), .Y(n5095) );
  INVX1 U4999 ( .A(n6295), .Y(n5094) );
  INVX1 U5000 ( .A(n5095), .Y(n6319) );
  NAND3X1 U5001 ( .A(n4191), .B(n3846), .C(n3878), .Y(n6375) );
  NAND3X1 U5002 ( .A(n4189), .B(n3848), .C(n3033), .Y(n6295) );
  INVX1 U5003 ( .A(N185), .Y(n5096) );
  OAI21X1 U5004 ( .A(n5097), .B(n32), .C(n5188), .Y(n5189) );
  INVX1 U5005 ( .A(n5612), .Y(n5097) );
  INVX1 U5006 ( .A(n5232), .Y(n5098) );
  AND2X2 U5007 ( .A(n909), .B(n6457), .Y(n5099) );
  INVX4 U5008 ( .A(n5099), .Y(n6402) );
  NAND3X1 U5009 ( .A(n581), .B(n596), .C(n655), .Y(n5100) );
  INVX1 U5010 ( .A(n5100), .Y(n6239) );
  NAND3X1 U5011 ( .A(n4176), .B(n602), .C(n554), .Y(n5101) );
  INVX1 U5012 ( .A(n5101), .Y(n5936) );
  AND2X2 U5013 ( .A(n5675), .B(\mem<50><3> ), .Y(n5102) );
  INVX1 U5014 ( .A(n5102), .Y(n5213) );
  AND2X2 U5015 ( .A(n3956), .B(n5615), .Y(n5103) );
  INVX1 U5016 ( .A(n5103), .Y(n5188) );
  INVX1 U5017 ( .A(N188), .Y(n5104) );
  INVX1 U5018 ( .A(N190), .Y(n5105) );
  NAND3X1 U5019 ( .A(n1147), .B(n5106), .C(n1704), .Y(n5107) );
  INVX1 U5020 ( .A(n5995), .Y(n5106) );
  INVX1 U5021 ( .A(n5107), .Y(n6017) );
  NAND3X1 U5022 ( .A(n5108), .B(n1146), .C(n4220), .Y(n5109) );
  INVX1 U5023 ( .A(n5831), .Y(n5108) );
  INVX1 U5024 ( .A(n5109), .Y(n5858) );
  AND2X2 U5025 ( .A(n5679), .B(\mem<40><3> ), .Y(n5110) );
  INVX1 U5026 ( .A(n5110), .Y(n5198) );
  AND2X2 U5027 ( .A(n3988), .B(\mem<56><3> ), .Y(n5111) );
  INVX1 U5028 ( .A(n5111), .Y(n5161) );
  INVX1 U5029 ( .A(n5522), .Y(n5112) );
  INVX1 U5030 ( .A(n5748), .Y(n5114) );
  INVX1 U5031 ( .A(n5114), .Y(n5115) );
  INVX1 U5032 ( .A(n5144), .Y(n5116) );
  INVX1 U5033 ( .A(n3653), .Y(n5117) );
  INVX1 U5034 ( .A(n5116), .Y(n5118) );
  INVX1 U5035 ( .A(n5117), .Y(n5119) );
  INVX1 U5036 ( .A(n6456), .Y(n5120) );
  INVX1 U5037 ( .A(n5134), .Y(n5121) );
  INVX1 U5038 ( .A(n5120), .Y(n5122) );
  INVX1 U5039 ( .A(n5117), .Y(n5123) );
  INVX1 U5040 ( .A(n5117), .Y(n5124) );
  INVX1 U5041 ( .A(n5116), .Y(n5125) );
  INVX1 U5042 ( .A(n5123), .Y(n5127) );
  INVX1 U5043 ( .A(n5124), .Y(n5130) );
  INVX1 U5044 ( .A(n5124), .Y(n5131) );
  INVX1 U5045 ( .A(n5118), .Y(n5134) );
  INVX1 U5046 ( .A(n5146), .Y(n5135) );
  INVX1 U5047 ( .A(n5147), .Y(n5136) );
  INVX1 U5048 ( .A(n165), .Y(n5137) );
  INVX1 U5049 ( .A(n165), .Y(n5139) );
  INVX1 U5050 ( .A(n3653), .Y(n5140) );
  INVX1 U5051 ( .A(n5748), .Y(n5142) );
  INVX1 U5052 ( .A(n5136), .Y(n5143) );
  INVX1 U5053 ( .A(n3654), .Y(n5144) );
  INVX1 U5054 ( .A(n3655), .Y(n5145) );
  INVX1 U5055 ( .A(n5145), .Y(n5146) );
  INVX1 U5056 ( .A(n5145), .Y(n5147) );
  INVX1 U5057 ( .A(n5145), .Y(n5148) );
  INVX1 U5058 ( .A(n5144), .Y(n5149) );
  INVX1 U5059 ( .A(n82), .Y(n5748) );
  INVX1 U5060 ( .A(n5134), .Y(n6456) );
  MUX2X1 U5061 ( .B(\mem<47><2> ), .A(\mem<46><2> ), .S(n3947), .Y(n5342) );
  INVX4 U5062 ( .A(n5218), .Y(n5150) );
  MUX2X1 U5063 ( .B(n507), .A(n5339), .S(n5159), .Y(n5338) );
  INVX1 U5064 ( .A(n5649), .Y(n5159) );
  MUX2X1 U5065 ( .B(\mem<17><7> ), .A(\mem<16><7> ), .S(n5697), .Y(n5629) );
  MUX2X1 U5066 ( .B(n529), .A(n576), .S(n3959), .Y(N191) );
  MUX2X1 U5067 ( .B(\mem<39><7> ), .A(\mem<38><7> ), .S(n3958), .Y(n5614) );
  MUX2X1 U5068 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n5178), .Y(n5630) );
  INVX1 U5069 ( .A(n5154), .Y(n5152) );
  INVX1 U5070 ( .A(N177), .Y(n5155) );
  AND2X2 U5071 ( .A(n3664), .B(n5157), .Y(n5156) );
  MUX2X1 U5072 ( .B(n5426), .A(n619), .S(n5160), .Y(N189) );
  INVX1 U5073 ( .A(N182), .Y(n5160) );
  AND2X2 U5074 ( .A(n90), .B(n5714), .Y(n5157) );
  MUX2X1 U5075 ( .B(n5558), .A(n5557), .S(n5158), .Y(n5556) );
  MUX2X1 U5076 ( .B(n5633), .A(n5632), .S(n5159), .Y(n5631) );
  MUX2X1 U5077 ( .B(\mem<17><1> ), .A(\mem<16><1> ), .S(n3988), .Y(n5310) );
  NAND2X1 U5078 ( .A(\mem<57><3> ), .B(n5685), .Y(n5162) );
  INVX1 U5079 ( .A(n5710), .Y(n5163) );
  INVX1 U5080 ( .A(n5710), .Y(n5164) );
  INVX1 U5081 ( .A(n5710), .Y(n5699) );
  INVX1 U5082 ( .A(n5657), .Y(n5165) );
  INVX1 U5083 ( .A(n5164), .Y(n5176) );
  NAND2X1 U5084 ( .A(\mem<8><1> ), .B(n3997), .Y(n5166) );
  NAND2X1 U5085 ( .A(\mem<9><1> ), .B(n93), .Y(n5167) );
  MUX2X1 U5086 ( .B(\mem<41><7> ), .A(\mem<40><7> ), .S(n5674), .Y(n5610) );
  MUX2X1 U5087 ( .B(\mem<35><1> ), .A(\mem<34><1> ), .S(n3982), .Y(n5300) );
  MUX2X1 U5088 ( .B(\mem<58><7> ), .A(\mem<59><7> ), .S(n3966), .Y(n5598) );
  INVX1 U5089 ( .A(n5163), .Y(n5702) );
  MUX2X1 U5090 ( .B(\mem<41><6> ), .A(\mem<40><6> ), .S(n3934), .Y(n5557) );
  OR2X2 U5091 ( .A(n5169), .B(n176), .Y(n6176) );
  NAND2X1 U5092 ( .A(\mem<8><6> ), .B(n5170), .Y(n5171) );
  NAND2X1 U5093 ( .A(\mem<9><6> ), .B(n3991), .Y(n5172) );
  INVX1 U5094 ( .A(n3991), .Y(n5170) );
  INVX1 U5095 ( .A(n5653), .Y(n5173) );
  MUX2X1 U5096 ( .B(n5233), .A(n598), .S(n5648), .Y(n5232) );
  AND2X2 U5097 ( .A(n107), .B(n5216), .Y(n5174) );
  INVX1 U5098 ( .A(n5652), .Y(n5175) );
  MUX2X1 U5099 ( .B(\mem<43><1> ), .A(\mem<42><1> ), .S(n3988), .Y(n5294) );
  MUX2X1 U5100 ( .B(n532), .A(n520), .S(n5648), .Y(n5387) );
  INVX1 U5101 ( .A(n5164), .Y(n5177) );
  INVX1 U5102 ( .A(n5163), .Y(n5700) );
  MUX2X1 U5103 ( .B(n5620), .A(n5619), .S(n5648), .Y(n5618) );
  MUX2X1 U5104 ( .B(\mem<33><6> ), .A(\mem<32><6> ), .S(n5676), .Y(n5563) );
  MUX2X1 U5105 ( .B(\mem<61><6> ), .A(\mem<60><6> ), .S(n3954), .Y(n5540) );
  MUX2X1 U5106 ( .B(\mem<41><4> ), .A(\mem<40><4> ), .S(n3954), .Y(n5445) );
  INVX1 U5107 ( .A(n5183), .Y(n5184) );
  INVX1 U5108 ( .A(n5192), .Y(n5185) );
  INVX1 U5109 ( .A(n3948), .Y(n5192) );
  MUX2X1 U5110 ( .B(\mem<63><6> ), .A(\mem<62><6> ), .S(n3954), .Y(n5541) );
  MUX2X1 U5111 ( .B(\mem<13><1> ), .A(\mem<12><1> ), .S(n5186), .Y(n5314) );
  AND2X2 U5112 ( .A(n3995), .B(n591), .Y(n5187) );
  INVX1 U5113 ( .A(n5189), .Y(n5619) );
  MUX2X1 U5114 ( .B(\mem<45><6> ), .A(\mem<44><6> ), .S(n3954), .Y(n5554) );
  MUX2X1 U5115 ( .B(\mem<39><6> ), .A(\mem<38><6> ), .S(n3954), .Y(n5561) );
  AND2X2 U5116 ( .A(n4042), .B(n946), .Y(n6020) );
  INVX1 U5117 ( .A(n170), .Y(n5747) );
  MUX2X1 U5118 ( .B(\mem<49><6> ), .A(\mem<48><6> ), .S(n3954), .Y(n5549) );
  MUX2X1 U5119 ( .B(\mem<11><6> ), .A(\mem<10><6> ), .S(n3958), .Y(n5586) );
  INVX1 U5120 ( .A(n5657), .Y(n5191) );
  AND2X2 U5121 ( .A(n4044), .B(n948), .Y(n5863) );
  MUX2X1 U5122 ( .B(\mem<51><6> ), .A(\mem<50><6> ), .S(n5674), .Y(n5550) );
  INVX2 U5123 ( .A(n5742), .Y(n5741) );
  AND2X2 U5124 ( .A(N181), .B(N180), .Y(n5193) );
  INVX1 U5125 ( .A(n5193), .Y(n5773) );
  AND2X2 U5126 ( .A(n121), .B(\mem<20><6> ), .Y(n6273) );
  MUX2X1 U5127 ( .B(n5397), .A(n5387), .S(n3948), .Y(n5426) );
  AND2X2 U5128 ( .A(n5157), .B(n3683), .Y(n5194) );
  MUX2X1 U5129 ( .B(n511), .A(n5389), .S(n5195), .Y(n5388) );
  INVX1 U5130 ( .A(n5208), .Y(n5196) );
  INVX1 U5131 ( .A(n5655), .Y(n5208) );
  OR2X2 U5132 ( .A(n5197), .B(n3991), .Y(n5202) );
  NAND2X1 U5133 ( .A(\mem<54><3> ), .B(n5674), .Y(n5200) );
  NAND2X1 U5134 ( .A(\mem<55><3> ), .B(n3961), .Y(n5201) );
  NAND2X1 U5135 ( .A(\mem<59><3> ), .B(n5692), .Y(n5203) );
  INVX1 U5136 ( .A(n5655), .Y(n5204) );
  INVX4 U5137 ( .A(n5650), .Y(n5655) );
  INVX1 U5138 ( .A(n6439), .Y(n5205) );
  INVX1 U5139 ( .A(n5653), .Y(n5206) );
  MUX2X1 U5140 ( .B(\mem<49><5> ), .A(\mem<48><5> ), .S(n5678), .Y(n5490) );
  INVX1 U5141 ( .A(n6439), .Y(n5207) );
  INVX1 U5142 ( .A(n5219), .Y(n5746) );
  MUX2X1 U5143 ( .B(\mem<43><7> ), .A(\mem<42><7> ), .S(n91), .Y(n5611) );
  OR2X2 U5144 ( .A(N182), .B(N180), .Y(n5807) );
  NAND2X1 U5145 ( .A(\mem<48><3> ), .B(n3947), .Y(n5210) );
  NAND2X1 U5146 ( .A(\mem<49><3> ), .B(n5683), .Y(n5211) );
  MUX2X1 U5147 ( .B(n5494), .A(n5493), .S(n5212), .Y(n5492) );
  MUX2X1 U5148 ( .B(\mem<43><3> ), .A(\mem<42><3> ), .S(n3954), .Y(n5391) );
  INVX1 U5149 ( .A(n5757), .Y(n5651) );
  INVX1 U5150 ( .A(n264), .Y(n5650) );
  INVX1 U5151 ( .A(N182), .Y(n5218) );
  NAND2X1 U5152 ( .A(\mem<51><3> ), .B(n5179), .Y(n5214) );
  AND2X2 U5153 ( .A(n5711), .B(n3683), .Y(n5215) );
  AND2X2 U5154 ( .A(N178), .B(n5180), .Y(n5216) );
  INVX1 U5155 ( .A(n5704), .Y(n5706) );
  INVX1 U5156 ( .A(n3927), .Y(n6400) );
  MUX2X1 U5157 ( .B(n615), .A(n5454), .S(n5212), .Y(n5453) );
  MUX2X1 U5158 ( .B(n5471), .A(n5470), .S(n5658), .Y(n5469) );
  MUX2X1 U5159 ( .B(n614), .A(n584), .S(n5218), .Y(N186) );
  AND2X2 U5160 ( .A(n168), .B(n623), .Y(n5219) );
  MUX2X1 U5161 ( .B(\mem<11><1> ), .A(\mem<10><1> ), .S(n3958), .Y(n5317) );
  INVX1 U5162 ( .A(N182), .Y(n5220) );
  MUX2X1 U5163 ( .B(n5222), .A(n5223), .S(n5662), .Y(n5221) );
  MUX2X1 U5164 ( .B(n524), .A(n5225), .S(n5662), .Y(n5224) );
  MUX2X1 U5165 ( .B(n5227), .A(n5228), .S(n5662), .Y(n5226) );
  MUX2X1 U5166 ( .B(n5230), .A(n5231), .S(n5662), .Y(n5229) );
  MUX2X1 U5167 ( .B(n5235), .A(n5236), .S(n5662), .Y(n5234) );
  MUX2X1 U5168 ( .B(n5238), .A(n5239), .S(n5662), .Y(n5237) );
  MUX2X1 U5169 ( .B(n5241), .A(n5242), .S(n5662), .Y(n5240) );
  MUX2X1 U5170 ( .B(n5244), .A(n5245), .S(n5662), .Y(n5243) );
  MUX2X1 U5171 ( .B(n5248), .A(n5249), .S(n5663), .Y(n5247) );
  MUX2X1 U5172 ( .B(n5251), .A(n5252), .S(n5663), .Y(n5250) );
  MUX2X1 U5173 ( .B(n5254), .A(n5255), .S(n5663), .Y(n5253) );
  MUX2X1 U5174 ( .B(n5257), .A(n5258), .S(n5663), .Y(n5256) );
  MUX2X1 U5175 ( .B(n5260), .A(n574), .S(n5649), .Y(n5259) );
  MUX2X1 U5176 ( .B(n5262), .A(n5263), .S(n5663), .Y(n5261) );
  MUX2X1 U5177 ( .B(n5265), .A(n5266), .S(n5663), .Y(n5264) );
  MUX2X1 U5178 ( .B(n5268), .A(n5269), .S(n5663), .Y(n5267) );
  MUX2X1 U5179 ( .B(n589), .A(n599), .S(n5150), .Y(N192) );
  MUX2X1 U5180 ( .B(n5276), .A(n5277), .S(n5663), .Y(n5275) );
  MUX2X1 U5181 ( .B(n5279), .A(n5280), .S(n5663), .Y(n5278) );
  MUX2X1 U5182 ( .B(n5282), .A(n5283), .S(n5663), .Y(n5281) );
  MUX2X1 U5183 ( .B(n5285), .A(n5286), .S(n5663), .Y(n5284) );
  MUX2X1 U5184 ( .B(n5288), .A(n501), .S(n5649), .Y(n5287) );
  MUX2X1 U5185 ( .B(n5290), .A(n5291), .S(n5664), .Y(n5289) );
  MUX2X1 U5186 ( .B(n5293), .A(n5294), .S(n5664), .Y(n5292) );
  MUX2X1 U5187 ( .B(n5296), .A(n5297), .S(n5664), .Y(n5295) );
  MUX2X1 U5188 ( .B(n5299), .A(n5300), .S(n5664), .Y(n5298) );
  MUX2X1 U5189 ( .B(n577), .A(n579), .S(n5649), .Y(n5301) );
  MUX2X1 U5190 ( .B(n5305), .A(n512), .S(n5664), .Y(n5304) );
  MUX2X1 U5191 ( .B(n5307), .A(n5308), .S(n5664), .Y(n5306) );
  MUX2X1 U5192 ( .B(n5314), .A(n5315), .S(n5664), .Y(n5313) );
  MUX2X1 U5193 ( .B(n578), .A(n5317), .S(n5664), .Y(n5316) );
  MUX2X1 U5194 ( .B(n5319), .A(n5320), .S(n5664), .Y(n5318) );
  MUX2X1 U5195 ( .B(n5322), .A(n5323), .S(n5664), .Y(n5321) );
  MUX2X1 U5196 ( .B(n587), .A(n5325), .S(n5649), .Y(n5324) );
  MUX2X1 U5197 ( .B(n5330), .A(n5331), .S(n5665), .Y(n5329) );
  MUX2X1 U5198 ( .B(n5333), .A(n5334), .S(n5665), .Y(n5332) );
  MUX2X1 U5199 ( .B(n5336), .A(n5337), .S(n5665), .Y(n5335) );
  MUX2X1 U5200 ( .B(n5341), .A(n5342), .S(n5665), .Y(n5340) );
  MUX2X1 U5201 ( .B(n5344), .A(n5345), .S(n5665), .Y(n5343) );
  MUX2X1 U5202 ( .B(n5347), .A(n5348), .S(n5665), .Y(n5346) );
  MUX2X1 U5203 ( .B(n5350), .A(n5351), .S(n5665), .Y(n5349) );
  MUX2X1 U5204 ( .B(n5355), .A(n5356), .S(n5665), .Y(n5354) );
  MUX2X1 U5205 ( .B(n5358), .A(n5359), .S(n5665), .Y(n5357) );
  MUX2X1 U5206 ( .B(n5361), .A(n5362), .S(n5665), .Y(n5360) );
  MUX2X1 U5207 ( .B(n5364), .A(n5365), .S(n5665), .Y(n5363) );
  MUX2X1 U5208 ( .B(n5367), .A(n5368), .S(n5649), .Y(n5366) );
  MUX2X1 U5209 ( .B(n5370), .A(n5371), .S(n5666), .Y(n5369) );
  MUX2X1 U5210 ( .B(n5373), .A(n536), .S(n5666), .Y(n5372) );
  MUX2X1 U5211 ( .B(n5375), .A(n503), .S(n5666), .Y(n5374) );
  MUX2X1 U5212 ( .B(n5377), .A(n5378), .S(n5666), .Y(n5376) );
  MUX2X1 U5213 ( .B(n575), .A(n609), .S(n5666), .Y(n5383) );
  MUX2X1 U5214 ( .B(n613), .A(n618), .S(n5666), .Y(n5386) );
  MUX2X1 U5215 ( .B(n606), .A(n5391), .S(n5666), .Y(n5390) );
  MUX2X1 U5216 ( .B(n5393), .A(n5394), .S(n5666), .Y(n5392) );
  MUX2X1 U5217 ( .B(n586), .A(n522), .S(n5649), .Y(n5397) );
  MUX2X1 U5218 ( .B(n5402), .A(n5403), .S(n5667), .Y(n5401) );
  MUX2X1 U5219 ( .B(n5405), .A(n5406), .S(n5667), .Y(n5404) );
  MUX2X1 U5220 ( .B(n5411), .A(n604), .S(n5649), .Y(n5410) );
  MUX2X1 U5221 ( .B(n5413), .A(n5414), .S(n5667), .Y(n5412) );
  MUX2X1 U5222 ( .B(n5419), .A(n5420), .S(n5667), .Y(n5418) );
  MUX2X1 U5223 ( .B(n5422), .A(n5423), .S(n5667), .Y(n5421) );
  MUX2X1 U5224 ( .B(n5428), .A(n5429), .S(n5667), .Y(n5427) );
  MUX2X1 U5225 ( .B(n5431), .A(n5432), .S(n5667), .Y(n5430) );
  MUX2X1 U5226 ( .B(n5434), .A(n5435), .S(n5667), .Y(n5433) );
  MUX2X1 U5227 ( .B(n5437), .A(n5438), .S(n5667), .Y(n5436) );
  MUX2X1 U5228 ( .B(n5442), .A(n5443), .S(n5668), .Y(n5441) );
  MUX2X1 U5229 ( .B(n5448), .A(n5449), .S(n5668), .Y(n5447) );
  MUX2X1 U5230 ( .B(n5451), .A(n5452), .S(n5668), .Y(n5450) );
  MUX2X1 U5231 ( .B(n5456), .A(n5457), .S(n5668), .Y(n5455) );
  MUX2X1 U5232 ( .B(n5459), .A(n5460), .S(n5668), .Y(n5458) );
  MUX2X1 U5233 ( .B(n5462), .A(n5463), .S(n5668), .Y(n5461) );
  MUX2X1 U5234 ( .B(n5465), .A(n5466), .S(n5668), .Y(n5464) );
  MUX2X1 U5235 ( .B(n514), .A(n5468), .S(n5649), .Y(n5467) );
  MUX2X1 U5236 ( .B(n5473), .A(n518), .S(n5668), .Y(n5472) );
  MUX2X1 U5237 ( .B(n504), .A(n5475), .S(n5668), .Y(n5474) );
  MUX2X1 U5238 ( .B(n5477), .A(n5478), .S(n5668), .Y(n5476) );
  MUX2X1 U5239 ( .B(n506), .A(n513), .S(n5649), .Y(n5479) );
  MUX2X1 U5240 ( .B(n505), .A(n515), .S(n5150), .Y(N188) );
  MUX2X1 U5241 ( .B(n5481), .A(n5482), .S(n5669), .Y(n5480) );
  MUX2X1 U5242 ( .B(n5484), .A(n5485), .S(n5669), .Y(n5483) );
  MUX2X1 U5243 ( .B(n5487), .A(n5488), .S(n5669), .Y(n5486) );
  MUX2X1 U5244 ( .B(n5490), .A(n5491), .S(n5669), .Y(n5489) );
  MUX2X1 U5245 ( .B(n5496), .A(n5497), .S(n5669), .Y(n5495) );
  MUX2X1 U5246 ( .B(n5502), .A(n5503), .S(n5669), .Y(n5501) );
  MUX2X1 U5247 ( .B(n5505), .A(n5506), .S(n5669), .Y(n5504) );
  MUX2X1 U5248 ( .B(n5508), .A(n5509), .S(n5649), .Y(n5507) );
  MUX2X1 U5249 ( .B(n5511), .A(n5512), .S(n5669), .Y(n5510) );
  MUX2X1 U5250 ( .B(n5517), .A(n5518), .S(n5669), .Y(n5516) );
  MUX2X1 U5251 ( .B(n5520), .A(n5521), .S(n5669), .Y(n5519) );
  MUX2X1 U5252 ( .B(n5525), .A(n5526), .S(n5670), .Y(n5524) );
  MUX2X1 U5253 ( .B(n5528), .A(n5529), .S(n5670), .Y(n5527) );
  MUX2X1 U5254 ( .B(n5531), .A(n5532), .S(n5670), .Y(n5530) );
  MUX2X1 U5255 ( .B(n5534), .A(n5535), .S(n5670), .Y(n5533) );
  MUX2X1 U5256 ( .B(n5537), .A(n5538), .S(n5649), .Y(n5536) );
  MUX2X1 U5257 ( .B(n620), .A(n607), .S(n5150), .Y(N187) );
  MUX2X1 U5258 ( .B(n5540), .A(n5541), .S(n5670), .Y(n5539) );
  MUX2X1 U5259 ( .B(n5543), .A(n5544), .S(n5670), .Y(n5542) );
  MUX2X1 U5260 ( .B(n5546), .A(n5547), .S(n5670), .Y(n5545) );
  MUX2X1 U5261 ( .B(n5549), .A(n5550), .S(n5670), .Y(n5548) );
  MUX2X1 U5262 ( .B(n5552), .A(n611), .S(n5649), .Y(n5551) );
  MUX2X1 U5263 ( .B(n5560), .A(n5561), .S(n5670), .Y(n5559) );
  MUX2X1 U5264 ( .B(n5571), .A(n5572), .S(n5671), .Y(n5570) );
  MUX2X1 U5265 ( .B(n5577), .A(n5578), .S(n5671), .Y(n5576) );
  MUX2X1 U5266 ( .B(n5580), .A(n5581), .S(n5649), .Y(n5579) );
  MUX2X1 U5267 ( .B(n5583), .A(n5584), .S(n5671), .Y(n5582) );
  MUX2X1 U5268 ( .B(n582), .A(n5586), .S(n5671), .Y(n5585) );
  MUX2X1 U5269 ( .B(n5588), .A(n5589), .S(n5671), .Y(n5587) );
  MUX2X1 U5270 ( .B(n5591), .A(n5592), .S(n5671), .Y(n5590) );
  MUX2X1 U5271 ( .B(n525), .A(n5595), .S(n5671), .Y(n5594) );
  MUX2X1 U5272 ( .B(n5600), .A(n5601), .S(n5671), .Y(n5599) );
  MUX2X1 U5273 ( .B(n5605), .A(n5606), .S(n5649), .Y(n5604) );
  MUX2X1 U5274 ( .B(n5613), .A(n5614), .S(n5672), .Y(n5612) );
  MUX2X1 U5275 ( .B(n5616), .A(n5617), .S(n5672), .Y(n5615) );
  MUX2X1 U5276 ( .B(n502), .A(n5622), .S(n5672), .Y(n5621) );
  MUX2X1 U5277 ( .B(n509), .A(n5624), .S(n5672), .Y(n5623) );
  MUX2X1 U5278 ( .B(n5626), .A(n5627), .S(n5672), .Y(n5625) );
  MUX2X1 U5279 ( .B(n5629), .A(n5630), .S(n5672), .Y(n5628) );
  MUX2X1 U5280 ( .B(n5635), .A(n5636), .S(n5672), .Y(n5634) );
  MUX2X1 U5281 ( .B(n5638), .A(n5639), .S(n5672), .Y(n5637) );
  MUX2X1 U5282 ( .B(n5641), .A(n5642), .S(n5672), .Y(n5640) );
  MUX2X1 U5283 ( .B(n5644), .A(n5645), .S(n5672), .Y(n5643) );
  MUX2X1 U5284 ( .B(n5647), .A(n585), .S(n5649), .Y(n5646) );
  MUX2X1 U5285 ( .B(\mem<62><0> ), .A(\mem<63><0> ), .S(n5680), .Y(n5223) );
  MUX2X1 U5286 ( .B(\mem<60><0> ), .A(\mem<61><0> ), .S(n5692), .Y(n5222) );
  MUX2X1 U5287 ( .B(n5224), .A(n5221), .S(n5657), .Y(n5233) );
  MUX2X1 U5288 ( .B(\mem<54><0> ), .A(\mem<55><0> ), .S(n3989), .Y(n5228) );
  MUX2X1 U5289 ( .B(\mem<52><0> ), .A(\mem<53><0> ), .S(n106), .Y(n5227) );
  MUX2X1 U5290 ( .B(\mem<50><0> ), .A(\mem<51><0> ), .S(n5692), .Y(n5231) );
  MUX2X1 U5291 ( .B(\mem<48><0> ), .A(\mem<49><0> ), .S(n5687), .Y(n5230) );
  MUX2X1 U5292 ( .B(\mem<46><0> ), .A(\mem<47><0> ), .S(n3961), .Y(n5236) );
  MUX2X1 U5293 ( .B(\mem<44><0> ), .A(\mem<45><0> ), .S(n93), .Y(n5235) );
  MUX2X1 U5294 ( .B(\mem<42><0> ), .A(\mem<43><0> ), .S(n5685), .Y(n5239) );
  MUX2X1 U5295 ( .B(\mem<40><0> ), .A(\mem<41><0> ), .S(n5680), .Y(n5238) );
  MUX2X1 U5296 ( .B(\mem<38><0> ), .A(\mem<39><0> ), .S(n5689), .Y(n5242) );
  MUX2X1 U5297 ( .B(\mem<36><0> ), .A(\mem<37><0> ), .S(n5685), .Y(n5241) );
  MUX2X1 U5298 ( .B(\mem<34><0> ), .A(\mem<35><0> ), .S(n5692), .Y(n5245) );
  MUX2X1 U5299 ( .B(\mem<32><0> ), .A(\mem<33><0> ), .S(n5685), .Y(n5244) );
  MUX2X1 U5300 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n3935), .Y(n5249) );
  MUX2X1 U5301 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n5689), .Y(n5252) );
  MUX2X1 U5302 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n5689), .Y(n5251) );
  MUX2X1 U5303 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n167), .Y(n5255) );
  MUX2X1 U5304 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n5689), .Y(n5258) );
  MUX2X1 U5305 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n5689), .Y(n5257) );
  MUX2X1 U5306 ( .B(n5256), .A(n5253), .S(n5657), .Y(n5260) );
  MUX2X1 U5307 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n3957), .Y(n5263) );
  MUX2X1 U5308 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n5689), .Y(n5262) );
  MUX2X1 U5309 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n5689), .Y(n5266) );
  MUX2X1 U5310 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n5689), .Y(n5265) );
  MUX2X1 U5311 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n5681), .Y(n5269) );
  MUX2X1 U5312 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n5683), .Y(n5268) );
  MUX2X1 U5313 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n5689), .Y(n5272) );
  MUX2X1 U5314 ( .B(n5270), .A(n5267), .S(n5657), .Y(n5274) );
  MUX2X1 U5315 ( .B(\mem<60><1> ), .A(\mem<61><1> ), .S(n5683), .Y(n5276) );
  MUX2X1 U5316 ( .B(\mem<58><1> ), .A(\mem<59><1> ), .S(n5683), .Y(n5280) );
  MUX2X1 U5317 ( .B(\mem<56><1> ), .A(\mem<57><1> ), .S(n5683), .Y(n5279) );
  MUX2X1 U5318 ( .B(\mem<54><1> ), .A(\mem<55><1> ), .S(n5696), .Y(n5283) );
  MUX2X1 U5319 ( .B(\mem<52><1> ), .A(\mem<53><1> ), .S(n5683), .Y(n5282) );
  MUX2X1 U5320 ( .B(\mem<50><1> ), .A(\mem<51><1> ), .S(n5696), .Y(n5286) );
  MUX2X1 U5321 ( .B(\mem<48><1> ), .A(\mem<49><1> ), .S(n5694), .Y(n5285) );
  MUX2X1 U5322 ( .B(n5284), .A(n5281), .S(n5657), .Y(n5288) );
  MUX2X1 U5323 ( .B(\mem<46><1> ), .A(\mem<47><1> ), .S(n5683), .Y(n5291) );
  MUX2X1 U5324 ( .B(\mem<44><1> ), .A(\mem<45><1> ), .S(n5696), .Y(n5290) );
  MUX2X1 U5325 ( .B(\mem<40><1> ), .A(\mem<41><1> ), .S(n5694), .Y(n5293) );
  MUX2X1 U5326 ( .B(\mem<38><1> ), .A(\mem<39><1> ), .S(n5681), .Y(n5297) );
  MUX2X1 U5327 ( .B(\mem<36><1> ), .A(\mem<37><1> ), .S(n5695), .Y(n5296) );
  MUX2X1 U5328 ( .B(\mem<32><1> ), .A(\mem<33><1> ), .S(n5694), .Y(n5299) );
  MUX2X1 U5329 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n5695), .Y(n5303) );
  MUX2X1 U5330 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n5681), .Y(n5305) );
  MUX2X1 U5331 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n5694), .Y(n5308) );
  MUX2X1 U5332 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n5681), .Y(n5307) );
  MUX2X1 U5333 ( .B(n5309), .A(n5306), .S(n5656), .Y(n5312) );
  MUX2X1 U5334 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n5686), .Y(n5315) );
  MUX2X1 U5335 ( .B(n5316), .A(n5313), .S(n5656), .Y(n5325) );
  MUX2X1 U5336 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n5179), .Y(n5319) );
  MUX2X1 U5337 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n5686), .Y(n5323) );
  MUX2X1 U5338 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n5694), .Y(n5322) );
  MUX2X1 U5339 ( .B(\mem<62><2> ), .A(\mem<63><2> ), .S(n5693), .Y(n5328) );
  MUX2X1 U5340 ( .B(\mem<60><2> ), .A(\mem<61><2> ), .S(n5692), .Y(n5327) );
  MUX2X1 U5341 ( .B(\mem<58><2> ), .A(\mem<59><2> ), .S(n5680), .Y(n5331) );
  MUX2X1 U5342 ( .B(\mem<56><2> ), .A(\mem<57><2> ), .S(n5685), .Y(n5330) );
  MUX2X1 U5343 ( .B(\mem<54><2> ), .A(\mem<55><2> ), .S(n5168), .Y(n5334) );
  MUX2X1 U5344 ( .B(\mem<52><2> ), .A(\mem<53><2> ), .S(n5684), .Y(n5333) );
  MUX2X1 U5345 ( .B(\mem<50><2> ), .A(\mem<51><2> ), .S(n5168), .Y(n5337) );
  MUX2X1 U5346 ( .B(\mem<48><2> ), .A(\mem<49><2> ), .S(n5681), .Y(n5336) );
  MUX2X1 U5347 ( .B(n5335), .A(n5332), .S(n5656), .Y(n5339) );
  MUX2X1 U5348 ( .B(\mem<44><2> ), .A(\mem<45><2> ), .S(n5684), .Y(n5341) );
  MUX2X1 U5349 ( .B(\mem<42><2> ), .A(\mem<43><2> ), .S(n5684), .Y(n5345) );
  MUX2X1 U5350 ( .B(\mem<40><2> ), .A(\mem<41><2> ), .S(n5689), .Y(n5344) );
  MUX2X1 U5351 ( .B(\mem<38><2> ), .A(\mem<39><2> ), .S(n5684), .Y(n5348) );
  MUX2X1 U5352 ( .B(\mem<36><2> ), .A(\mem<37><2> ), .S(n3935), .Y(n5347) );
  MUX2X1 U5353 ( .B(\mem<34><2> ), .A(\mem<35><2> ), .S(n5684), .Y(n5351) );
  MUX2X1 U5354 ( .B(\mem<32><2> ), .A(\mem<33><2> ), .S(n5684), .Y(n5350) );
  MUX2X1 U5355 ( .B(n5349), .A(n5346), .S(n5656), .Y(n5353) );
  MUX2X1 U5356 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n5684), .Y(n5356) );
  MUX2X1 U5357 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n5684), .Y(n5355) );
  MUX2X1 U5358 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n5684), .Y(n5358) );
  MUX2X1 U5359 ( .B(n5357), .A(n5354), .S(n5656), .Y(n5368) );
  MUX2X1 U5360 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n5684), .Y(n5362) );
  MUX2X1 U5361 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n3935), .Y(n5361) );
  MUX2X1 U5362 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n5684), .Y(n5365) );
  MUX2X1 U5363 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n5684), .Y(n5364) );
  MUX2X1 U5364 ( .B(n5363), .A(n5360), .S(n5656), .Y(n5367) );
  MUX2X1 U5365 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n5685), .Y(n5371) );
  MUX2X1 U5366 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n5680), .Y(n5370) );
  MUX2X1 U5367 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n5685), .Y(n5373) );
  MUX2X1 U5368 ( .B(n5372), .A(n5369), .S(n5656), .Y(n5380) );
  MUX2X1 U5369 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n5680), .Y(n5375) );
  MUX2X1 U5370 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n5178), .Y(n5378) );
  MUX2X1 U5371 ( .B(\mem<38><3> ), .A(\mem<39><3> ), .S(n5686), .Y(n5394) );
  MUX2X1 U5372 ( .B(\mem<36><3> ), .A(\mem<37><3> ), .S(n5696), .Y(n5393) );
  MUX2X1 U5373 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n5681), .Y(n5400) );
  MUX2X1 U5374 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n5694), .Y(n5399) );
  MUX2X1 U5375 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n3961), .Y(n5403) );
  MUX2X1 U5376 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n3961), .Y(n5402) );
  MUX2X1 U5377 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n5683), .Y(n5406) );
  MUX2X1 U5378 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n3961), .Y(n5405) );
  MUX2X1 U5379 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n3961), .Y(n5409) );
  MUX2X1 U5380 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n5696), .Y(n5408) );
  MUX2X1 U5381 ( .B(n5407), .A(n5404), .S(n5655), .Y(n5411) );
  MUX2X1 U5382 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n5696), .Y(n5413) );
  MUX2X1 U5383 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n5681), .Y(n5417) );
  MUX2X1 U5384 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n5683), .Y(n5416) );
  MUX2X1 U5385 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n5688), .Y(n5420) );
  MUX2X1 U5386 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n5681), .Y(n5419) );
  MUX2X1 U5387 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n5682), .Y(n5423) );
  MUX2X1 U5388 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n5682), .Y(n5422) );
  MUX2X1 U5389 ( .B(n5421), .A(n5418), .S(n5655), .Y(n5425) );
  MUX2X1 U5390 ( .B(\mem<62><4> ), .A(\mem<63><4> ), .S(n5683), .Y(n5429) );
  MUX2X1 U5391 ( .B(\mem<60><4> ), .A(\mem<61><4> ), .S(n5694), .Y(n5428) );
  MUX2X1 U5392 ( .B(\mem<58><4> ), .A(\mem<59><4> ), .S(n5688), .Y(n5432) );
  MUX2X1 U5393 ( .B(\mem<56><4> ), .A(\mem<57><4> ), .S(n3989), .Y(n5431) );
  MUX2X1 U5394 ( .B(\mem<54><4> ), .A(\mem<55><4> ), .S(n5688), .Y(n5435) );
  MUX2X1 U5395 ( .B(\mem<52><4> ), .A(\mem<53><4> ), .S(n5694), .Y(n5434) );
  MUX2X1 U5396 ( .B(\mem<48><4> ), .A(\mem<49><4> ), .S(n5688), .Y(n5437) );
  MUX2X1 U5397 ( .B(n5436), .A(n5433), .S(n5655), .Y(n5440) );
  MUX2X1 U5398 ( .B(\mem<46><4> ), .A(\mem<47><4> ), .S(n5695), .Y(n5443) );
  MUX2X1 U5399 ( .B(\mem<44><4> ), .A(\mem<45><4> ), .S(n5696), .Y(n5442) );
  MUX2X1 U5400 ( .B(\mem<42><4> ), .A(\mem<43><4> ), .S(n5690), .Y(n5446) );
  MUX2X1 U5401 ( .B(\mem<38><4> ), .A(\mem<39><4> ), .S(n5689), .Y(n5449) );
  MUX2X1 U5402 ( .B(\mem<36><4> ), .A(\mem<37><4> ), .S(n5689), .Y(n5448) );
  MUX2X1 U5403 ( .B(\mem<34><4> ), .A(\mem<35><4> ), .S(n5688), .Y(n5452) );
  MUX2X1 U5404 ( .B(\mem<32><4> ), .A(\mem<33><4> ), .S(n5695), .Y(n5451) );
  MUX2X1 U5405 ( .B(n5450), .A(n5447), .S(n5655), .Y(n5454) );
  MUX2X1 U5406 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n5696), .Y(n5457) );
  MUX2X1 U5407 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n5168), .Y(n5456) );
  MUX2X1 U5408 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n5689), .Y(n5460) );
  MUX2X1 U5409 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n5689), .Y(n5459) );
  MUX2X1 U5410 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n5689), .Y(n5463) );
  MUX2X1 U5411 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n5689), .Y(n5462) );
  MUX2X1 U5412 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n5689), .Y(n5466) );
  MUX2X1 U5413 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n5689), .Y(n5465) );
  MUX2X1 U5414 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n5685), .Y(n5471) );
  MUX2X1 U5415 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n5680), .Y(n5470) );
  MUX2X1 U5416 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n5689), .Y(n5473) );
  MUX2X1 U5417 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n5696), .Y(n5475) );
  MUX2X1 U5418 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n5689), .Y(n5478) );
  MUX2X1 U5419 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n5689), .Y(n5477) );
  MUX2X1 U5420 ( .B(\mem<62><5> ), .A(\mem<63><5> ), .S(n167), .Y(n5482) );
  MUX2X1 U5421 ( .B(\mem<60><5> ), .A(\mem<61><5> ), .S(n5692), .Y(n5481) );
  MUX2X1 U5422 ( .B(\mem<58><5> ), .A(\mem<59><5> ), .S(n5680), .Y(n5485) );
  MUX2X1 U5423 ( .B(\mem<56><5> ), .A(\mem<57><5> ), .S(n167), .Y(n5484) );
  MUX2X1 U5424 ( .B(n5483), .A(n5480), .S(n5654), .Y(n5494) );
  MUX2X1 U5425 ( .B(\mem<54><5> ), .A(\mem<55><5> ), .S(n167), .Y(n5488) );
  MUX2X1 U5426 ( .B(\mem<52><5> ), .A(\mem<53><5> ), .S(n5683), .Y(n5487) );
  MUX2X1 U5427 ( .B(\mem<50><5> ), .A(\mem<51><5> ), .S(n3966), .Y(n5491) );
  MUX2X1 U5428 ( .B(n5489), .A(n5486), .S(n5654), .Y(n5493) );
  MUX2X1 U5429 ( .B(\mem<46><5> ), .A(\mem<47><5> ), .S(n5692), .Y(n5497) );
  MUX2X1 U5430 ( .B(\mem<44><5> ), .A(\mem<45><5> ), .S(n5681), .Y(n5496) );
  MUX2X1 U5431 ( .B(\mem<42><5> ), .A(\mem<43><5> ), .S(n5692), .Y(n5500) );
  MUX2X1 U5432 ( .B(\mem<40><5> ), .A(\mem<41><5> ), .S(n5692), .Y(n5499) );
  MUX2X1 U5433 ( .B(n5498), .A(n5495), .S(n5654), .Y(n5509) );
  MUX2X1 U5434 ( .B(\mem<38><5> ), .A(\mem<39><5> ), .S(n5693), .Y(n5503) );
  MUX2X1 U5435 ( .B(\mem<36><5> ), .A(\mem<37><5> ), .S(n5680), .Y(n5502) );
  MUX2X1 U5436 ( .B(\mem<34><5> ), .A(\mem<35><5> ), .S(n5692), .Y(n5506) );
  MUX2X1 U5437 ( .B(\mem<32><5> ), .A(\mem<33><5> ), .S(n5680), .Y(n5505) );
  MUX2X1 U5438 ( .B(n5504), .A(n5501), .S(n5654), .Y(n5508) );
  MUX2X1 U5439 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n5693), .Y(n5512) );
  MUX2X1 U5440 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n5692), .Y(n5511) );
  MUX2X1 U5441 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n5693), .Y(n5515) );
  MUX2X1 U5442 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n5685), .Y(n5514) );
  MUX2X1 U5443 ( .B(n5513), .A(n5510), .S(n5654), .Y(n5523) );
  MUX2X1 U5444 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n5693), .Y(n5518) );
  MUX2X1 U5445 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n5693), .Y(n5517) );
  MUX2X1 U5446 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n5680), .Y(n5521) );
  MUX2X1 U5447 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n5693), .Y(n5520) );
  MUX2X1 U5448 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n5693), .Y(n5526) );
  MUX2X1 U5449 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n5693), .Y(n5525) );
  MUX2X1 U5450 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n5690), .Y(n5529) );
  MUX2X1 U5451 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n5685), .Y(n5528) );
  MUX2X1 U5452 ( .B(n5527), .A(n5524), .S(n5654), .Y(n5538) );
  MUX2X1 U5453 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n5692), .Y(n5532) );
  MUX2X1 U5454 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n5685), .Y(n5531) );
  MUX2X1 U5455 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n5685), .Y(n5535) );
  MUX2X1 U5456 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n5685), .Y(n5534) );
  MUX2X1 U5457 ( .B(n5533), .A(n5530), .S(n5654), .Y(n5537) );
  MUX2X1 U5458 ( .B(\mem<58><6> ), .A(\mem<59><6> ), .S(n5692), .Y(n5544) );
  MUX2X1 U5459 ( .B(\mem<56><6> ), .A(\mem<57><6> ), .S(n5680), .Y(n5543) );
  MUX2X1 U5460 ( .B(\mem<54><6> ), .A(\mem<55><6> ), .S(n5685), .Y(n5547) );
  MUX2X1 U5461 ( .B(\mem<52><6> ), .A(\mem<53><6> ), .S(n5680), .Y(n5546) );
  MUX2X1 U5462 ( .B(n5548), .A(n5545), .S(n5653), .Y(n5552) );
  MUX2X1 U5463 ( .B(\mem<46><6> ), .A(\mem<47><6> ), .S(n5692), .Y(n5555) );
  MUX2X1 U5464 ( .B(\mem<36><6> ), .A(\mem<37><6> ), .S(n5690), .Y(n5560) );
  MUX2X1 U5465 ( .B(\mem<34><6> ), .A(\mem<35><6> ), .S(n5685), .Y(n5564) );
  MUX2X1 U5466 ( .B(n5562), .A(n5559), .S(n5653), .Y(n5566) );
  MUX2X1 U5467 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n5694), .Y(n5569) );
  MUX2X1 U5468 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n5692), .Y(n5568) );
  MUX2X1 U5469 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n5682), .Y(n5571) );
  MUX2X1 U5470 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n5683), .Y(n5575) );
  MUX2X1 U5471 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n5680), .Y(n5574) );
  MUX2X1 U5472 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n5682), .Y(n5578) );
  MUX2X1 U5473 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n5680), .Y(n5577) );
  MUX2X1 U5474 ( .B(n5576), .A(n5573), .S(n5653), .Y(n5580) );
  MUX2X1 U5475 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n5694), .Y(n5584) );
  MUX2X1 U5476 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n5683), .Y(n5583) );
  MUX2X1 U5477 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n5696), .Y(n5589) );
  MUX2X1 U5478 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n5168), .Y(n5588) );
  MUX2X1 U5479 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n5696), .Y(n5592) );
  MUX2X1 U5480 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n5168), .Y(n5591) );
  MUX2X1 U5481 ( .B(\mem<56><7> ), .A(\mem<57><7> ), .S(n5682), .Y(n5597) );
  MUX2X1 U5482 ( .B(\mem<52><7> ), .A(\mem<53><7> ), .S(n5695), .Y(n5600) );
  MUX2X1 U5483 ( .B(\mem<50><7> ), .A(\mem<51><7> ), .S(n5682), .Y(n5603) );
  MUX2X1 U5484 ( .B(n5602), .A(n5599), .S(n5653), .Y(n5605) );
  MUX2X1 U5485 ( .B(\mem<46><7> ), .A(\mem<47><7> ), .S(n5686), .Y(n5608) );
  MUX2X1 U5486 ( .B(n5609), .A(n5607), .S(n5653), .Y(n5620) );
  MUX2X1 U5487 ( .B(\mem<36><7> ), .A(\mem<37><7> ), .S(n3957), .Y(n5613) );
  MUX2X1 U5488 ( .B(\mem<34><7> ), .A(\mem<35><7> ), .S(n5686), .Y(n5617) );
  MUX2X1 U5489 ( .B(\mem<32><7> ), .A(\mem<33><7> ), .S(n5686), .Y(n5616) );
  MUX2X1 U5490 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n5686), .Y(n5622) );
  MUX2X1 U5491 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n5178), .Y(n5624) );
  MUX2X1 U5492 ( .B(n5623), .A(n5621), .S(n5652), .Y(n5633) );
  MUX2X1 U5493 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n5696), .Y(n5626) );
  MUX2X1 U5494 ( .B(n5628), .A(n5625), .S(n5652), .Y(n5632) );
  MUX2X1 U5495 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n5695), .Y(n5636) );
  MUX2X1 U5496 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n5695), .Y(n5635) );
  MUX2X1 U5497 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n5696), .Y(n5639) );
  MUX2X1 U5498 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n5695), .Y(n5638) );
  MUX2X1 U5499 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n5696), .Y(n5642) );
  MUX2X1 U5500 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n5695), .Y(n5641) );
  MUX2X1 U5501 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n5695), .Y(n5645) );
  MUX2X1 U5502 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n5695), .Y(n5644) );
  INVX8 U5503 ( .A(n5673), .Y(n5658) );
  INVX8 U5504 ( .A(n5673), .Y(n5659) );
  INVX8 U5505 ( .A(n5673), .Y(n5660) );
  INVX8 U5506 ( .A(n5673), .Y(n5661) );
  INVX8 U5507 ( .A(n5661), .Y(n5662) );
  INVX8 U5508 ( .A(n5661), .Y(n5663) );
  INVX8 U5509 ( .A(n5661), .Y(n5664) );
  INVX8 U5510 ( .A(n5660), .Y(n5665) );
  INVX8 U5511 ( .A(n5660), .Y(n5666) );
  INVX8 U5512 ( .A(n5660), .Y(n5667) );
  INVX8 U5513 ( .A(n5659), .Y(n5668) );
  INVX8 U5514 ( .A(n5659), .Y(n5669) );
  INVX8 U5515 ( .A(n5659), .Y(n5670) );
  INVX8 U5516 ( .A(n5658), .Y(n5671) );
  INVX8 U5517 ( .A(n5658), .Y(n5672) );
  INVX8 U5518 ( .A(n5677), .Y(n5680) );
  INVX8 U5519 ( .A(n5678), .Y(n5681) );
  INVX8 U5520 ( .A(n78), .Y(n5683) );
  INVX8 U5521 ( .A(n3992), .Y(n5684) );
  INVX8 U5522 ( .A(n5677), .Y(n5685) );
  INVX8 U5523 ( .A(n5679), .Y(n5689) );
  INVX8 U5524 ( .A(n5677), .Y(n5692) );
  INVX8 U5525 ( .A(n5676), .Y(n5693) );
  INVX8 U5526 ( .A(n81), .Y(n5695) );
  INVX8 U5527 ( .A(n5675), .Y(n5696) );
  NOR3X1 U5528 ( .A(n5704), .B(n32), .C(n3940), .Y(n5703) );
  NOR3X1 U5529 ( .A(n5706), .B(n5155), .C(n32), .Y(n5705) );
  AND2X2 U5530 ( .A(n5714), .B(n403), .Y(n5707) );
  INVX1 U5531 ( .A(n5708), .Y(n5709) );
  INVX1 U5532 ( .A(n5807), .Y(n5832) );
  AND2X2 U5533 ( .A(n5711), .B(n923), .Y(n5710) );
  AND2X2 U5534 ( .A(n5714), .B(n90), .Y(n5711) );
  INVX1 U5535 ( .A(\addr<11> ), .Y(n5771) );
  BUFX2 U5536 ( .A(\addr<13> ), .Y(n5712) );
  AND2X2 U5537 ( .A(n5157), .B(n3662), .Y(n5713) );
  INVX1 U5538 ( .A(n5194), .Y(n6429) );
  AND2X2 U5539 ( .A(n950), .B(n5771), .Y(n5714) );
  BUFX4 U5540 ( .A(n4944), .Y(n5715) );
  INVX8 U5541 ( .A(n3659), .Y(n5718) );
  INVX8 U5542 ( .A(n5726), .Y(n5720) );
  INVX8 U5543 ( .A(n5726), .Y(n5721) );
  INVX8 U5544 ( .A(n5725), .Y(n5723) );
  INVX8 U5545 ( .A(n5734), .Y(n5730) );
  INVX8 U5546 ( .A(n5733), .Y(n5731) );
  INVX8 U5547 ( .A(n5737), .Y(n5733) );
  INVX8 U5548 ( .A(n5736), .Y(n5734) );
  INVX8 U5549 ( .A(n5736), .Y(n5735) );
  INVX8 U5550 ( .A(n5741), .Y(n5739) );
  INVX8 U5551 ( .A(n5187), .Y(n5740) );
  INVX8 U5552 ( .A(n87), .Y(n5749) );
  AOI22X1 U5553 ( .A(\mem<29><0> ), .B(n233), .C(\mem<31><0> ), .D(n223), .Y(
        n5763) );
  OR2X2 U5554 ( .A(n264), .B(N178), .Y(n5761) );
  AOI22X1 U5555 ( .A(\mem<27><0> ), .B(n188), .C(\mem<25><0> ), .D(n92), .Y(
        n5762) );
  NOR2X1 U5556 ( .A(n118), .B(n5764), .Y(n5765) );
  AOI21X1 U5557 ( .A(\mem<30><0> ), .B(n5731), .C(n5765), .Y(n5770) );
  OR2X2 U5558 ( .A(n5757), .B(N178), .Y(n5766) );
  NOR2X1 U5559 ( .A(n5721), .B(n5767), .Y(n5768) );
  AOI21X1 U5560 ( .A(\mem<26><0> ), .B(n5130), .C(n5768), .Y(n5769) );
  NAND3X1 U5561 ( .A(\addr<14> ), .B(\addr<11> ), .C(n5712), .Y(n5775) );
  NAND3X1 U5562 ( .A(\addr<10> ), .B(\addr<12> ), .C(\addr<9> ), .Y(n5774) );
  NAND2X1 U5563 ( .A(\mem<60><0> ), .B(n149), .Y(n5776) );
  OAI21X1 U5564 ( .A(n5733), .B(n5777), .C(n5776), .Y(n5781) );
  NAND2X1 U5565 ( .A(\mem<63><0> ), .B(n227), .Y(n5778) );
  OAI21X1 U5566 ( .A(n5115), .B(n5779), .C(n5778), .Y(n5780) );
  OAI21X1 U5567 ( .A(n175), .B(n5782), .C(n4046), .Y(n5783) );
  AOI21X1 U5568 ( .A(\mem<57><0> ), .B(n92), .C(n5783), .Y(n5784) );
  AOI22X1 U5569 ( .A(\mem<0><0> ), .B(n549), .C(n58), .D(n3026), .Y(n5785) );
  OAI21X1 U5570 ( .A(n625), .B(n5709), .C(n5785), .Y(n5831) );
  NOR2X1 U5571 ( .A(n131), .B(n5786), .Y(n5787) );
  AOI21X1 U5572 ( .A(\mem<14><0> ), .B(n5731), .C(n5787), .Y(n5795) );
  OAI21X1 U5573 ( .A(n5718), .B(n5788), .C(n972), .Y(n5791) );
  OAI21X1 U5574 ( .A(n259), .B(n5789), .C(n974), .Y(n5790) );
  NOR2X1 U5575 ( .A(n5724), .B(n5792), .Y(n5793) );
  AOI21X1 U5576 ( .A(\mem<10><0> ), .B(n5128), .C(n5793), .Y(n5794) );
  NOR2X1 U5577 ( .A(n125), .B(n5796), .Y(n5797) );
  AOI21X1 U5578 ( .A(\mem<38><0> ), .B(n5732), .C(n5797), .Y(n5806) );
  NAND2X1 U5579 ( .A(\mem<35><0> ), .B(n187), .Y(n5798) );
  OAI21X1 U5580 ( .A(n5719), .B(n5799), .C(n5798), .Y(n5802) );
  OAI21X1 U5581 ( .A(n234), .B(n5800), .C(n976), .Y(n5801) );
  NOR2X1 U5582 ( .A(n5724), .B(n5803), .Y(n5804) );
  AOI21X1 U5583 ( .A(\mem<34><0> ), .B(n5141), .C(n5804), .Y(n5805) );
  AOI22X1 U5584 ( .A(n23), .B(n454), .C(n96), .D(n488), .Y(n5830) );
  NOR2X1 U5585 ( .A(n117), .B(n5808), .Y(n5809) );
  AOI21X1 U5586 ( .A(\mem<22><0> ), .B(n5731), .C(n5809), .Y(n5817) );
  OAI21X1 U5587 ( .A(n5718), .B(n5810), .C(n978), .Y(n5813) );
  OAI21X1 U5588 ( .A(n250), .B(n5811), .C(n980), .Y(n5812) );
  NOR2X1 U5589 ( .A(n5723), .B(n5814), .Y(n5815) );
  AOI21X1 U5590 ( .A(\mem<18><0> ), .B(n5126), .C(n5815), .Y(n5816) );
  NOR2X1 U5591 ( .A(n125), .B(n5818), .Y(n5819) );
  AOI21X1 U5592 ( .A(\mem<54><0> ), .B(n5731), .C(n5819), .Y(n5828) );
  NAND2X1 U5593 ( .A(\mem<51><0> ), .B(n203), .Y(n5820) );
  OAI21X1 U5594 ( .A(n5718), .B(n5821), .C(n5820), .Y(n5824) );
  OAI21X1 U5595 ( .A(n251), .B(n5822), .C(n982), .Y(n5823) );
  NOR2X1 U5596 ( .A(n5723), .B(n5825), .Y(n5826) );
  AOI21X1 U5597 ( .A(\mem<50><0> ), .B(n5148), .C(n5826), .Y(n5827) );
  AOI22X1 U5598 ( .A(n5194), .B(n456), .C(n5701), .D(n410), .Y(n5829) );
  OAI21X1 U5599 ( .A(n5720), .B(n5833), .C(n4048), .Y(n5836) );
  OAI21X1 U5600 ( .A(n5735), .B(n5834), .C(n984), .Y(n5835) );
  NAND2X1 U5601 ( .A(\mem<3><0> ), .B(n195), .Y(n5837) );
  OAI21X1 U5602 ( .A(n5749), .B(n5838), .C(n5837), .Y(n5842) );
  NAND2X1 U5603 ( .A(\mem<7><0> ), .B(n225), .Y(n5839) );
  OAI21X1 U5604 ( .A(n5739), .B(n5840), .C(n5839), .Y(n5841) );
  NAND3X1 U5605 ( .A(n5843), .B(N180), .C(N182), .Y(n5844) );
  OAI21X1 U5606 ( .A(n5720), .B(n5845), .C(n4050), .Y(n5849) );
  NAND2X1 U5607 ( .A(\mem<44><0> ), .B(n156), .Y(n5846) );
  OAI21X1 U5608 ( .A(n5735), .B(n5847), .C(n5846), .Y(n5848) );
  NAND2X1 U5609 ( .A(\mem<43><0> ), .B(n201), .Y(n5850) );
  OAI21X1 U5610 ( .A(n5749), .B(n5851), .C(n5850), .Y(n5855) );
  NAND2X1 U5611 ( .A(\mem<47><0> ), .B(n227), .Y(n5852) );
  OAI21X1 U5612 ( .A(n5740), .B(n5853), .C(n5852), .Y(n5854) );
  AOI22X1 U5613 ( .A(n33), .B(n1680), .C(n3657), .D(n3028), .Y(n5857) );
  AOI21X1 U5614 ( .A(n5858), .B(n1649), .C(n5715), .Y(\data_out<0> ) );
  NAND2X1 U5615 ( .A(\mem<60><1> ), .B(n160), .Y(n5861) );
  NAND2X1 U5616 ( .A(\mem<62><1> ), .B(n5732), .Y(n5860) );
  AOI22X1 U5617 ( .A(\mem<63><1> ), .B(n227), .C(\mem<58><1> ), .D(n5114), .Y(
        n5859) );
  OAI21X1 U5618 ( .A(n414), .B(n3010), .C(n59), .Y(n5870) );
  AOI22X1 U5619 ( .A(\mem<27><1> ), .B(n186), .C(\mem<25><1> ), .D(n92), .Y(
        n5862) );
  NOR2X1 U5620 ( .A(n126), .B(n5864), .Y(n5865) );
  AOI21X1 U5621 ( .A(\mem<30><1> ), .B(n5731), .C(n5865), .Y(n5869) );
  NOR2X1 U5622 ( .A(n5723), .B(n5866), .Y(n5867) );
  AOI21X1 U5623 ( .A(\mem<26><1> ), .B(n5142), .C(n5867), .Y(n5868) );
  NOR2X1 U5624 ( .A(n143), .B(n5871), .Y(n5872) );
  AOI21X1 U5625 ( .A(\mem<14><1> ), .B(n5731), .C(n5872), .Y(n5881) );
  NAND2X1 U5626 ( .A(\mem<11><1> ), .B(n197), .Y(n5873) );
  OAI21X1 U5627 ( .A(n5717), .B(n5874), .C(n5873), .Y(n5877) );
  OAI21X1 U5628 ( .A(n263), .B(n5875), .C(n266), .Y(n5876) );
  NOR2X1 U5629 ( .A(n5723), .B(n5878), .Y(n5879) );
  AOI21X1 U5630 ( .A(\mem<10><1> ), .B(n5149), .C(n5879), .Y(n5880) );
  NOR2X1 U5631 ( .A(n113), .B(n5882), .Y(n5883) );
  AOI21X1 U5632 ( .A(\mem<38><1> ), .B(n5731), .C(n5883), .Y(n5891) );
  OAI21X1 U5633 ( .A(n5719), .B(n5884), .C(n986), .Y(n5887) );
  OAI21X1 U5634 ( .A(n258), .B(n5885), .C(n988), .Y(n5886) );
  NOR2X1 U5635 ( .A(n5723), .B(n5888), .Y(n5889) );
  AOI21X1 U5636 ( .A(\mem<34><1> ), .B(n5138), .C(n5889), .Y(n5890) );
  AOI22X1 U5637 ( .A(n472), .B(n210), .C(n416), .D(n3913), .Y(n5914) );
  NOR2X1 U5638 ( .A(n120), .B(n5892), .Y(n5893) );
  AOI21X1 U5639 ( .A(\mem<22><1> ), .B(n5731), .C(n5893), .Y(n5902) );
  NAND2X1 U5640 ( .A(\mem<19><1> ), .B(n195), .Y(n5894) );
  OAI21X1 U5641 ( .A(n5717), .B(n5895), .C(n5894), .Y(n5898) );
  OAI21X1 U5642 ( .A(n261), .B(n5896), .C(n990), .Y(n5897) );
  NOR2X1 U5643 ( .A(n5723), .B(n5899), .Y(n5900) );
  AOI21X1 U5644 ( .A(\mem<18><1> ), .B(n3655), .C(n5900), .Y(n5901) );
  AOI21X1 U5645 ( .A(\mem<54><1> ), .B(n5731), .C(n5903), .Y(n5912) );
  NAND2X1 U5646 ( .A(\mem<51><1> ), .B(n203), .Y(n5904) );
  OAI21X1 U5647 ( .A(n101), .B(n5905), .C(n5904), .Y(n5908) );
  OAI21X1 U5648 ( .A(n251), .B(n5906), .C(n992), .Y(n5907) );
  NOR2X1 U5649 ( .A(n5723), .B(n5909), .Y(n5910) );
  AOI21X1 U5650 ( .A(\mem<50><1> ), .B(n5139), .C(n5910), .Y(n5911) );
  AOI22X1 U5651 ( .A(n458), .B(n5215), .C(n3024), .D(n5701), .Y(n5913) );
  OAI21X1 U5652 ( .A(n5720), .B(n5915), .C(n4052), .Y(n5919) );
  NAND2X1 U5653 ( .A(\mem<4><1> ), .B(n164), .Y(n5916) );
  OAI21X1 U5654 ( .A(n5735), .B(n5917), .C(n5916), .Y(n5918) );
  NAND2X1 U5655 ( .A(\mem<3><1> ), .B(n202), .Y(n5920) );
  NAND2X1 U5656 ( .A(\mem<7><1> ), .B(n223), .Y(n5922) );
  OAI21X1 U5657 ( .A(n5740), .B(n5923), .C(n5922), .Y(n5924) );
  OAI21X1 U5658 ( .A(n5720), .B(n5926), .C(n4054), .Y(n5930) );
  NAND2X1 U5659 ( .A(\mem<44><1> ), .B(n151), .Y(n5927) );
  OAI21X1 U5660 ( .A(n5735), .B(n5928), .C(n5927), .Y(n5929) );
  OAI21X1 U5661 ( .A(n5749), .B(n5931), .C(n4056), .Y(n5934) );
  OAI21X1 U5662 ( .A(n5740), .B(n5932), .C(n994), .Y(n5933) );
  AOI22X1 U5663 ( .A(n33), .B(n1682), .C(n3657), .D(n638), .Y(n5935) );
  AOI21X1 U5664 ( .A(n5936), .B(n1650), .C(n5715), .Y(\data_out<1> ) );
  NAND2X1 U5665 ( .A(\mem<57><2> ), .B(n5753), .Y(n5937) );
  NAND3X1 U5666 ( .A(n5937), .B(n4224), .C(n4179), .Y(n5941) );
  NAND2X1 U5667 ( .A(\mem<60><2> ), .B(n152), .Y(n5940) );
  NAND2X1 U5668 ( .A(\mem<62><2> ), .B(n5732), .Y(n5939) );
  AOI22X1 U5669 ( .A(\mem<63><2> ), .B(n223), .C(\mem<58><2> ), .D(n5131), .Y(
        n5938) );
  OAI21X1 U5670 ( .A(n4213), .B(n3012), .C(n3928), .Y(n5950) );
  AOI22X1 U5671 ( .A(\mem<29><2> ), .B(n233), .C(\mem<31><2> ), .D(n226), .Y(
        n5943) );
  AOI22X1 U5672 ( .A(\mem<27><2> ), .B(n172), .C(\mem<25><2> ), .D(n103), .Y(
        n5942) );
  NOR2X1 U5673 ( .A(n112), .B(n5944), .Y(n5945) );
  AOI21X1 U5674 ( .A(\mem<30><2> ), .B(n5731), .C(n5945), .Y(n5949) );
  NOR2X1 U5675 ( .A(n5723), .B(n5946), .Y(n5947) );
  AOI21X1 U5676 ( .A(\mem<26><2> ), .B(n5130), .C(n5947), .Y(n5948) );
  NAND3X1 U5677 ( .A(n1151), .B(n4253), .C(n5950), .Y(n5995) );
  NOR2X1 U5678 ( .A(n133), .B(n5951), .Y(n5952) );
  AOI21X1 U5679 ( .A(\mem<14><2> ), .B(n5731), .C(n5952), .Y(n5961) );
  OAI21X1 U5680 ( .A(n5718), .B(n5953), .C(n996), .Y(n5957) );
  NAND2X1 U5681 ( .A(\mem<15><2> ), .B(n77), .Y(n5954) );
  OAI21X1 U5682 ( .A(n262), .B(n5955), .C(n5954), .Y(n5956) );
  NOR2X1 U5683 ( .A(n5723), .B(n5958), .Y(n5959) );
  AOI21X1 U5684 ( .A(\mem<10><2> ), .B(n5126), .C(n5959), .Y(n5960) );
  NOR2X1 U5685 ( .A(n123), .B(n5962), .Y(n5963) );
  AOI21X1 U5686 ( .A(\mem<38><2> ), .B(n5731), .C(n5963), .Y(n5971) );
  OAI21X1 U5687 ( .A(n5719), .B(n5964), .C(n998), .Y(n5967) );
  OAI21X1 U5688 ( .A(n237), .B(n5965), .C(n1000), .Y(n5966) );
  NOR2X1 U5689 ( .A(n5723), .B(n5968), .Y(n5969) );
  AOI21X1 U5690 ( .A(\mem<34><2> ), .B(n5133), .C(n5969), .Y(n5970) );
  AOI22X1 U5691 ( .A(n474), .B(n204), .C(n420), .D(n212), .Y(n5994) );
  NOR2X1 U5692 ( .A(n118), .B(n5972), .Y(n5973) );
  AOI21X1 U5693 ( .A(\mem<22><2> ), .B(n5731), .C(n5973), .Y(n5981) );
  OAI21X1 U5694 ( .A(n5719), .B(n5974), .C(n1002), .Y(n5977) );
  OAI21X1 U5695 ( .A(n239), .B(n5975), .C(n1004), .Y(n5976) );
  NOR2X1 U5696 ( .A(n5723), .B(n5978), .Y(n5979) );
  AOI21X1 U5697 ( .A(\mem<18><2> ), .B(n5127), .C(n5979), .Y(n5980) );
  NOR2X1 U5698 ( .A(n115), .B(n5982), .Y(n5983) );
  AOI21X1 U5699 ( .A(\mem<54><2> ), .B(n5731), .C(n5983), .Y(n5992) );
  NAND2X1 U5700 ( .A(\mem<51><2> ), .B(n199), .Y(n5984) );
  OAI21X1 U5701 ( .A(n5718), .B(n5985), .C(n5984), .Y(n5988) );
  OAI21X1 U5702 ( .A(n240), .B(n5986), .C(n1006), .Y(n5987) );
  NOR2X1 U5703 ( .A(n5723), .B(n5989), .Y(n5990) );
  AOI21X1 U5704 ( .A(\mem<50><2> ), .B(n82), .C(n5990), .Y(n5991) );
  AOI22X1 U5705 ( .A(n5194), .B(n460), .C(n5701), .D(n490), .Y(n5993) );
  OAI21X1 U5706 ( .A(n5721), .B(n5996), .C(n4058), .Y(n5999) );
  OAI21X1 U5707 ( .A(n5735), .B(n5997), .C(n1008), .Y(n5998) );
  NAND2X1 U5708 ( .A(\mem<3><2> ), .B(n199), .Y(n6000) );
  OAI21X1 U5709 ( .A(n5750), .B(n6001), .C(n6000), .Y(n6005) );
  NAND2X1 U5710 ( .A(\mem<7><2> ), .B(n224), .Y(n6002) );
  OAI21X1 U5711 ( .A(n5740), .B(n6003), .C(n6002), .Y(n6004) );
  OAI21X1 U5712 ( .A(n5720), .B(n6006), .C(n4060), .Y(n6010) );
  NAND2X1 U5713 ( .A(\mem<44><2> ), .B(n164), .Y(n6007) );
  OAI21X1 U5714 ( .A(n5735), .B(n6008), .C(n6007), .Y(n6009) );
  NAND2X1 U5715 ( .A(\mem<43><2> ), .B(n185), .Y(n6011) );
  OAI21X1 U5716 ( .A(n5749), .B(n6012), .C(n6011), .Y(n6015) );
  OAI21X1 U5717 ( .A(n5739), .B(n6013), .C(n1010), .Y(n6014) );
  AOI22X1 U5718 ( .A(n6459), .B(n1684), .C(n3657), .D(n3030), .Y(n6016) );
  AOI21X1 U5719 ( .A(n6017), .B(n1651), .C(n5715), .Y(\data_out<2> ) );
  AOI22X1 U5720 ( .A(\mem<63><3> ), .B(n223), .C(\mem<58><3> ), .D(n166), .Y(
        n6018) );
  OAI21X1 U5721 ( .A(n424), .B(n484), .C(n58), .Y(n6027) );
  AOI22X1 U5722 ( .A(\mem<27><3> ), .B(n203), .C(\mem<25><3> ), .D(n92), .Y(
        n6019) );
  NOR2X1 U5723 ( .A(n124), .B(n6021), .Y(n6022) );
  AOI21X1 U5724 ( .A(\mem<30><3> ), .B(n5731), .C(n6022), .Y(n6026) );
  NOR2X1 U5725 ( .A(n5723), .B(n6023), .Y(n6024) );
  AOI21X1 U5726 ( .A(\mem<26><3> ), .B(n5137), .C(n6024), .Y(n6025) );
  NOR2X1 U5727 ( .A(n128), .B(n6028), .Y(n6029) );
  AOI21X1 U5728 ( .A(\mem<14><3> ), .B(n5731), .C(n6029), .Y(n6036) );
  NAND2X1 U5729 ( .A(\mem<11><3> ), .B(n169), .Y(n6030) );
  OAI21X1 U5730 ( .A(n5717), .B(n6031), .C(n6030), .Y(n6034) );
  OAI21X1 U5731 ( .A(n246), .B(n6032), .C(n268), .Y(n6033) );
  NOR2X1 U5732 ( .A(n139), .B(n6037), .Y(n6038) );
  AOI21X1 U5733 ( .A(\mem<38><3> ), .B(n5731), .C(n6038), .Y(n6044) );
  OAI21X1 U5734 ( .A(n5717), .B(n6039), .C(n34), .Y(n6042) );
  OAI21X1 U5735 ( .A(n247), .B(n6040), .C(n1012), .Y(n6041) );
  AOI22X1 U5736 ( .A(n476), .B(n45), .C(n4947), .D(n426), .Y(n6068) );
  NOR2X1 U5737 ( .A(n145), .B(n6045), .Y(n6046) );
  AOI21X1 U5738 ( .A(\mem<22><3> ), .B(n5731), .C(n6046), .Y(n6055) );
  NAND2X1 U5739 ( .A(\mem<19><3> ), .B(n188), .Y(n6047) );
  OAI21X1 U5740 ( .A(n5718), .B(n6048), .C(n6047), .Y(n6051) );
  OAI21X1 U5741 ( .A(n245), .B(n6049), .C(n1014), .Y(n6050) );
  NOR2X1 U5742 ( .A(n5722), .B(n6052), .Y(n6053) );
  AOI21X1 U5743 ( .A(\mem<18><3> ), .B(n5140), .C(n6053), .Y(n6054) );
  NOR2X1 U5744 ( .A(n115), .B(n6056), .Y(n6057) );
  AOI21X1 U5745 ( .A(\mem<54><3> ), .B(n5731), .C(n6057), .Y(n6066) );
  NAND2X1 U5746 ( .A(\mem<51><3> ), .B(n189), .Y(n6058) );
  OAI21X1 U5747 ( .A(n5717), .B(n6059), .C(n6058), .Y(n6062) );
  OAI21X1 U5748 ( .A(n257), .B(n6060), .C(n1016), .Y(n6061) );
  NOR2X1 U5749 ( .A(n5722), .B(n6063), .Y(n6064) );
  AOI21X1 U5750 ( .A(\mem<50><3> ), .B(n5116), .C(n6064), .Y(n6065) );
  AOI22X1 U5751 ( .A(n5215), .B(n462), .C(n211), .D(n492), .Y(n6067) );
  OAI21X1 U5752 ( .A(n5720), .B(n6069), .C(n4062), .Y(n6071) );
  OAI21X1 U5753 ( .A(n5749), .B(n6072), .C(n4064), .Y(n6076) );
  NAND2X1 U5754 ( .A(\mem<7><3> ), .B(n224), .Y(n6073) );
  OAI21X1 U5755 ( .A(n5739), .B(n6074), .C(n6073), .Y(n6075) );
  OAI21X1 U5756 ( .A(n5721), .B(n6077), .C(n4066), .Y(n6081) );
  NAND2X1 U5757 ( .A(\mem<44><3> ), .B(n153), .Y(n6078) );
  OAI21X1 U5758 ( .A(n5735), .B(n6079), .C(n6078), .Y(n6080) );
  NAND2X1 U5759 ( .A(\mem<43><3> ), .B(n197), .Y(n6082) );
  OAI21X1 U5760 ( .A(n5749), .B(n6083), .C(n6082), .Y(n6086) );
  OAI21X1 U5761 ( .A(n5739), .B(n6084), .C(n1018), .Y(n6085) );
  AOI22X1 U5762 ( .A(n6459), .B(n1678), .C(n68), .D(n646), .Y(n6087) );
  AOI21X1 U5763 ( .A(n6088), .B(n1652), .C(n5715), .Y(\data_out<3> ) );
  NAND2X1 U5764 ( .A(\mem<57><4> ), .B(n5753), .Y(n6089) );
  NAND3X1 U5765 ( .A(n6089), .B(n4227), .C(n4183), .Y(n6093) );
  NAND2X1 U5766 ( .A(\mem<60><4> ), .B(n163), .Y(n6092) );
  NAND2X1 U5767 ( .A(\mem<62><4> ), .B(n5732), .Y(n6091) );
  AOI22X1 U5768 ( .A(\mem<63><4> ), .B(n224), .C(\mem<58><4> ), .D(n5140), .Y(
        n6090) );
  OAI21X1 U5769 ( .A(n4215), .B(n3014), .C(n3928), .Y(n6102) );
  AOI22X1 U5770 ( .A(\mem<29><4> ), .B(n233), .C(\mem<31><4> ), .D(n227), .Y(
        n6095) );
  AOI22X1 U5771 ( .A(\mem<27><4> ), .B(n194), .C(\mem<25><4> ), .D(n92), .Y(
        n6094) );
  NOR2X1 U5772 ( .A(n119), .B(n6096), .Y(n6097) );
  AOI21X1 U5773 ( .A(\mem<30><4> ), .B(n5731), .C(n6097), .Y(n6101) );
  NOR2X1 U5774 ( .A(n5722), .B(n6098), .Y(n6099) );
  AOI21X1 U5775 ( .A(\mem<26><4> ), .B(n5143), .C(n6099), .Y(n6100) );
  NAND3X1 U5776 ( .A(n6102), .B(n4229), .C(n3876), .Y(n6143) );
  NOR2X1 U5777 ( .A(n141), .B(n6103), .Y(n6104) );
  AOI21X1 U5778 ( .A(\mem<14><4> ), .B(n5731), .C(n6104), .Y(n6112) );
  OAI21X1 U5779 ( .A(n5717), .B(n6105), .C(n1020), .Y(n6108) );
  OAI21X1 U5780 ( .A(n248), .B(n6106), .C(n1022), .Y(n6107) );
  NOR2X1 U5781 ( .A(n5722), .B(n6109), .Y(n6110) );
  AOI21X1 U5782 ( .A(\mem<10><4> ), .B(n5129), .C(n6110), .Y(n6111) );
  NOR2X1 U5783 ( .A(n135), .B(n6113), .Y(n6114) );
  AOI21X1 U5784 ( .A(\mem<38><4> ), .B(n5731), .C(n6114), .Y(n6121) );
  NAND2X1 U5785 ( .A(\mem<35><4> ), .B(n187), .Y(n6115) );
  OAI21X1 U5786 ( .A(n5718), .B(n6116), .C(n6115), .Y(n6119) );
  OAI21X1 U5787 ( .A(n5740), .B(n6117), .C(n1024), .Y(n6118) );
  AOI22X1 U5788 ( .A(n478), .B(n7), .C(n29), .D(n429), .Y(n6142) );
  NOR2X1 U5789 ( .A(n142), .B(n6122), .Y(n6123) );
  AOI21X1 U5790 ( .A(\mem<22><4> ), .B(n5731), .C(n6123), .Y(n6129) );
  OAI21X1 U5791 ( .A(n5717), .B(n6124), .C(n1026), .Y(n6127) );
  OAI21X1 U5792 ( .A(n252), .B(n6125), .C(n1028), .Y(n6126) );
  NOR2X1 U5793 ( .A(n114), .B(n6130), .Y(n6131) );
  AOI21X1 U5794 ( .A(\mem<54><4> ), .B(n5731), .C(n6131), .Y(n6140) );
  NAND2X1 U5795 ( .A(\mem<51><4> ), .B(n189), .Y(n6132) );
  OAI21X1 U5796 ( .A(n95), .B(n6133), .C(n6132), .Y(n6136) );
  OAI21X1 U5797 ( .A(n234), .B(n6134), .C(n1030), .Y(n6135) );
  NOR2X1 U5798 ( .A(n5722), .B(n6137), .Y(n6138) );
  AOI21X1 U5799 ( .A(\mem<50><4> ), .B(n5127), .C(n6138), .Y(n6139) );
  AOI22X1 U5800 ( .A(n5215), .B(n464), .C(n211), .D(n595), .Y(n6141) );
  OAI21X1 U5801 ( .A(n5720), .B(n6144), .C(n4068), .Y(n6148) );
  NAND2X1 U5802 ( .A(\mem<4><4> ), .B(n152), .Y(n6145) );
  OAI21X1 U5803 ( .A(n5734), .B(n6146), .C(n6145), .Y(n6147) );
  NAND2X1 U5804 ( .A(\mem<3><4> ), .B(n193), .Y(n6149) );
  OAI21X1 U5805 ( .A(n5751), .B(n6150), .C(n6149), .Y(n6153) );
  OAI21X1 U5806 ( .A(n5739), .B(n6151), .C(n1032), .Y(n6152) );
  OAI21X1 U5807 ( .A(n5721), .B(n6154), .C(n4070), .Y(n6158) );
  NAND2X1 U5808 ( .A(\mem<44><4> ), .B(n153), .Y(n6155) );
  OAI21X1 U5809 ( .A(n5734), .B(n6156), .C(n6155), .Y(n6157) );
  OAI21X1 U5810 ( .A(n5750), .B(n6159), .C(n4072), .Y(n6162) );
  OAI21X1 U5811 ( .A(n5739), .B(n6160), .C(n1034), .Y(n6161) );
  AOI22X1 U5812 ( .A(n33), .B(n1686), .C(n61), .D(n651), .Y(n6163) );
  AOI21X1 U5813 ( .A(n1657), .B(n4211), .C(n5715), .Y(\data_out<4> ) );
  AOI22X1 U5814 ( .A(\mem<63><5> ), .B(n3685), .C(\mem<58><5> ), .D(n5128), 
        .Y(n6164) );
  OAI21X1 U5815 ( .A(n432), .B(n486), .C(n3928), .Y(n6173) );
  AOI22X1 U5816 ( .A(\mem<29><5> ), .B(n233), .C(\mem<31><5> ), .D(n225), .Y(
        n6166) );
  AOI22X1 U5817 ( .A(\mem<27><5> ), .B(n173), .C(\mem<25><5> ), .D(n92), .Y(
        n6165) );
  NOR2X1 U5818 ( .A(n119), .B(n6167), .Y(n6168) );
  AOI21X1 U5819 ( .A(\mem<30><5> ), .B(n5731), .C(n6168), .Y(n6172) );
  NOR2X1 U5820 ( .A(n5722), .B(n6169), .Y(n6170) );
  AOI21X1 U5821 ( .A(\mem<26><5> ), .B(n5142), .C(n6170), .Y(n6171) );
  NOR2X1 U5822 ( .A(n134), .B(n6174), .Y(n6175) );
  AOI21X1 U5823 ( .A(\mem<14><5> ), .B(n5731), .C(n6175), .Y(n6184) );
  OAI21X1 U5824 ( .A(n5751), .B(n6177), .C(n6176), .Y(n6180) );
  OAI21X1 U5825 ( .A(n241), .B(n6178), .C(n1036), .Y(n6179) );
  NOR2X1 U5826 ( .A(n5722), .B(n6181), .Y(n6182) );
  AOI21X1 U5827 ( .A(\mem<10><5> ), .B(n5128), .C(n6182), .Y(n6183) );
  NOR2X1 U5828 ( .A(n123), .B(n6185), .Y(n6186) );
  AOI21X1 U5829 ( .A(\mem<38><5> ), .B(n5730), .C(n6186), .Y(n6195) );
  NAND2X1 U5830 ( .A(\mem<35><5> ), .B(n183), .Y(n6187) );
  OAI21X1 U5831 ( .A(n5719), .B(n6188), .C(n6187), .Y(n6191) );
  OAI21X1 U5832 ( .A(n236), .B(n6189), .C(n1038), .Y(n6190) );
  NOR2X1 U5833 ( .A(n5722), .B(n6192), .Y(n6193) );
  AOI21X1 U5834 ( .A(\mem<34><5> ), .B(n5148), .C(n6193), .Y(n6194) );
  AOI22X1 U5835 ( .A(n204), .B(n1676), .C(n434), .D(n212), .Y(n6217) );
  NOR2X1 U5836 ( .A(n112), .B(n6196), .Y(n6197) );
  AOI21X1 U5837 ( .A(\mem<22><5> ), .B(n5730), .C(n6197), .Y(n6205) );
  OAI21X1 U5838 ( .A(n101), .B(n6198), .C(n1040), .Y(n6201) );
  OAI21X1 U5839 ( .A(n260), .B(n6199), .C(n1042), .Y(n6200) );
  NOR2X1 U5840 ( .A(n5722), .B(n6202), .Y(n6203) );
  AOI21X1 U5841 ( .A(\mem<18><5> ), .B(n5146), .C(n6203), .Y(n6204) );
  NOR2X1 U5842 ( .A(n124), .B(n6206), .Y(n6207) );
  AOI21X1 U5843 ( .A(\mem<54><5> ), .B(n5730), .C(n6207), .Y(n6215) );
  OAI21X1 U5844 ( .A(n5719), .B(n6208), .C(n1044), .Y(n6211) );
  OAI21X1 U5845 ( .A(n262), .B(n6209), .C(n1046), .Y(n6210) );
  NOR2X1 U5846 ( .A(n5722), .B(n6212), .Y(n6213) );
  AOI21X1 U5847 ( .A(\mem<50><5> ), .B(n5137), .C(n6213), .Y(n6214) );
  AOI22X1 U5848 ( .A(n466), .B(n5215), .C(n5176), .D(n438), .Y(n6216) );
  OAI21X1 U5849 ( .A(n5721), .B(n6218), .C(n4074), .Y(n6222) );
  NAND2X1 U5850 ( .A(\mem<4><5> ), .B(n154), .Y(n6219) );
  OAI21X1 U5851 ( .A(n5734), .B(n6220), .C(n6219), .Y(n6221) );
  OAI21X1 U5852 ( .A(n5751), .B(n6223), .C(n4076), .Y(n6227) );
  NAND2X1 U5853 ( .A(\mem<7><5> ), .B(n226), .Y(n6224) );
  OAI21X1 U5854 ( .A(n5739), .B(n6225), .C(n6224), .Y(n6226) );
  OAI21X1 U5855 ( .A(n5720), .B(n6228), .C(n4078), .Y(n6232) );
  NAND2X1 U5856 ( .A(\mem<44><5> ), .B(n150), .Y(n6229) );
  OAI21X1 U5857 ( .A(n5734), .B(n6230), .C(n6229), .Y(n6231) );
  NAND2X1 U5858 ( .A(\mem<43><5> ), .B(n189), .Y(n6233) );
  OAI21X1 U5859 ( .A(n5749), .B(n6234), .C(n6233), .Y(n6237) );
  OAI21X1 U5860 ( .A(n5739), .B(n6235), .C(n1048), .Y(n6236) );
  AOI22X1 U5861 ( .A(n33), .B(n1688), .C(n3657), .D(n657), .Y(n6238) );
  AOI21X1 U5862 ( .A(n6239), .B(n1653), .C(n5715), .Y(\data_out<5> ) );
  NAND2X1 U5863 ( .A(\mem<57><6> ), .B(n5753), .Y(n6240) );
  NAND3X1 U5864 ( .A(n6240), .B(n4231), .C(n4187), .Y(n6244) );
  NAND2X1 U5865 ( .A(\mem<60><6> ), .B(n154), .Y(n6243) );
  NAND2X1 U5866 ( .A(\mem<62><6> ), .B(n5732), .Y(n6242) );
  AOI22X1 U5867 ( .A(\mem<63><6> ), .B(n226), .C(\mem<58><6> ), .D(n5127), .Y(
        n6241) );
  AOI22X1 U5868 ( .A(\mem<29><6> ), .B(n233), .C(\mem<31><6> ), .D(n226), .Y(
        n6246) );
  AOI22X1 U5869 ( .A(\mem<27><6> ), .B(n173), .C(\mem<25><6> ), .D(n92), .Y(
        n6245) );
  NOR2X1 U5870 ( .A(n117), .B(n6247), .Y(n6248) );
  AOI21X1 U5871 ( .A(\mem<30><6> ), .B(n5730), .C(n6248), .Y(n6252) );
  NOR2X1 U5872 ( .A(n5721), .B(n6249), .Y(n6250) );
  AOI21X1 U5873 ( .A(\mem<26><6> ), .B(n5130), .C(n6250), .Y(n6251) );
  NOR2X1 U5874 ( .A(n113), .B(n6253), .Y(n6254) );
  AOI21X1 U5875 ( .A(\mem<14><6> ), .B(n5730), .C(n6254), .Y(n6262) );
  OAI21X1 U5876 ( .A(n86), .B(n6255), .C(n1050), .Y(n6258) );
  OAI21X1 U5877 ( .A(n249), .B(n6256), .C(n1052), .Y(n6257) );
  NOR2X1 U5878 ( .A(n5722), .B(n6259), .Y(n6260) );
  AOI21X1 U5879 ( .A(\mem<10><6> ), .B(n5130), .C(n6260), .Y(n6261) );
  NOR2X1 U5880 ( .A(n129), .B(n6263), .Y(n6264) );
  AOI21X1 U5881 ( .A(\mem<38><6> ), .B(n5730), .C(n6264), .Y(n6272) );
  OAI21X1 U5882 ( .A(n5718), .B(n6265), .C(n1054), .Y(n6268) );
  OAI21X1 U5883 ( .A(n253), .B(n6266), .C(n1056), .Y(n6267) );
  NOR2X1 U5884 ( .A(n5721), .B(n6269), .Y(n6270) );
  AOI21X1 U5885 ( .A(\mem<34><6> ), .B(n5137), .C(n6270), .Y(n6271) );
  AOI22X1 U5886 ( .A(n480), .B(n204), .C(n5156), .D(n442), .Y(n6294) );
  AOI21X1 U5887 ( .A(\mem<22><6> ), .B(n5730), .C(n6273), .Y(n6281) );
  OAI21X1 U5888 ( .A(n86), .B(n6274), .C(n1058), .Y(n6277) );
  OAI21X1 U5889 ( .A(n260), .B(n6275), .C(n1060), .Y(n6276) );
  NOR2X1 U5890 ( .A(n5721), .B(n6278), .Y(n6279) );
  AOI21X1 U5891 ( .A(\mem<18><6> ), .B(n5147), .C(n6279), .Y(n6280) );
  NOR2X1 U5892 ( .A(n114), .B(n6282), .Y(n6283) );
  AOI21X1 U5893 ( .A(\mem<54><6> ), .B(n5730), .C(n6283), .Y(n6292) );
  NAND2X1 U5894 ( .A(\mem<51><6> ), .B(n186), .Y(n6284) );
  OAI21X1 U5895 ( .A(n86), .B(n6285), .C(n6284), .Y(n6288) );
  OAI21X1 U5896 ( .A(n235), .B(n6286), .C(n1062), .Y(n6287) );
  NOR2X1 U5897 ( .A(n5721), .B(n6289), .Y(n6290) );
  AOI21X1 U5898 ( .A(\mem<50><6> ), .B(n5128), .C(n6290), .Y(n6291) );
  AOI22X1 U5899 ( .A(n56), .B(n468), .C(n5702), .D(n494), .Y(n6293) );
  OAI21X1 U5900 ( .A(n5720), .B(n6296), .C(n4080), .Y(n6300) );
  NAND2X1 U5901 ( .A(\mem<4><6> ), .B(n162), .Y(n6297) );
  OAI21X1 U5902 ( .A(n5734), .B(n6298), .C(n6297), .Y(n6299) );
  NAND2X1 U5903 ( .A(\mem<3><6> ), .B(n183), .Y(n6301) );
  OAI21X1 U5904 ( .A(n5749), .B(n6302), .C(n6301), .Y(n6306) );
  NAND2X1 U5905 ( .A(\mem<7><6> ), .B(n224), .Y(n6303) );
  OAI21X1 U5906 ( .A(n5739), .B(n6304), .C(n6303), .Y(n6305) );
  OAI21X1 U5907 ( .A(n5720), .B(n6307), .C(n4082), .Y(n6311) );
  NAND2X1 U5908 ( .A(\mem<44><6> ), .B(n150), .Y(n6308) );
  OAI21X1 U5909 ( .A(n5734), .B(n6309), .C(n6308), .Y(n6310) );
  NAND2X1 U5910 ( .A(\mem<43><6> ), .B(n184), .Y(n6312) );
  OAI21X1 U5911 ( .A(n5749), .B(n6313), .C(n6312), .Y(n6317) );
  NAND2X1 U5912 ( .A(\mem<47><6> ), .B(n226), .Y(n6314) );
  OAI21X1 U5913 ( .A(n5739), .B(n6315), .C(n6314), .Y(n6316) );
  AOI22X1 U5914 ( .A(n33), .B(n1690), .C(n3657), .D(n661), .Y(n6318) );
  AOI21X1 U5915 ( .A(n6319), .B(n1654), .C(n5715), .Y(\data_out<6> ) );
  NAND2X1 U5916 ( .A(\mem<59><7> ), .B(n191), .Y(n6320) );
  NAND2X1 U5917 ( .A(\mem<60><7> ), .B(n158), .Y(n6323) );
  NAND2X1 U5918 ( .A(\mem<62><7> ), .B(n5732), .Y(n6322) );
  AOI22X1 U5919 ( .A(\mem<63><7> ), .B(n226), .C(\mem<58><7> ), .D(n5127), .Y(
        n6321) );
  AOI22X1 U5920 ( .A(\mem<29><7> ), .B(n233), .C(\mem<31><7> ), .D(n225), .Y(
        n6325) );
  AOI22X1 U5921 ( .A(\mem<27><7> ), .B(n193), .C(\mem<25><7> ), .D(n103), .Y(
        n6324) );
  NOR2X1 U5922 ( .A(n138), .B(n6326), .Y(n6327) );
  AOI21X1 U5923 ( .A(\mem<30><7> ), .B(n5730), .C(n6327), .Y(n6331) );
  NOR2X1 U5924 ( .A(n5721), .B(n6328), .Y(n6329) );
  AOI21X1 U5925 ( .A(\mem<26><7> ), .B(n5131), .C(n6329), .Y(n6330) );
  NOR2X1 U5926 ( .A(n130), .B(n6332), .Y(n6333) );
  AOI21X1 U5927 ( .A(\mem<14><7> ), .B(n5730), .C(n6333), .Y(n6341) );
  OAI21X1 U5928 ( .A(n5718), .B(n6334), .C(n1064), .Y(n6337) );
  OAI21X1 U5929 ( .A(n238), .B(n6335), .C(n1066), .Y(n6336) );
  NOR2X1 U5930 ( .A(n5721), .B(n6338), .Y(n6339) );
  AOI21X1 U5931 ( .A(\mem<10><7> ), .B(n5132), .C(n6339), .Y(n6340) );
  NOR2X1 U5932 ( .A(n136), .B(n6342), .Y(n6343) );
  AOI21X1 U5933 ( .A(\mem<38><7> ), .B(n5730), .C(n6343), .Y(n6351) );
  OAI21X1 U5934 ( .A(n5719), .B(n6344), .C(n270), .Y(n6347) );
  OAI21X1 U5935 ( .A(n241), .B(n6345), .C(n1068), .Y(n6346) );
  NOR2X1 U5936 ( .A(n5722), .B(n6348), .Y(n6349) );
  AOI21X1 U5937 ( .A(\mem<34><7> ), .B(n5139), .C(n6349), .Y(n6350) );
  AOI22X1 U5938 ( .A(n482), .B(n210), .C(n5156), .D(n446), .Y(n6374) );
  NOR2X1 U5939 ( .A(n126), .B(n6352), .Y(n6353) );
  AOI21X1 U5940 ( .A(\mem<22><7> ), .B(n5730), .C(n6353), .Y(n6361) );
  OAI21X1 U5941 ( .A(n5718), .B(n6354), .C(n1070), .Y(n6357) );
  OAI21X1 U5942 ( .A(n259), .B(n6355), .C(n1072), .Y(n6356) );
  NOR2X1 U5943 ( .A(n5721), .B(n6358), .Y(n6359) );
  AOI21X1 U5944 ( .A(\mem<18><7> ), .B(n5131), .C(n6359), .Y(n6360) );
  NOR2X1 U5945 ( .A(n115), .B(n6362), .Y(n6363) );
  AOI21X1 U5946 ( .A(\mem<54><7> ), .B(n5730), .C(n6363), .Y(n6372) );
  NAND2X1 U5947 ( .A(\mem<51><7> ), .B(n203), .Y(n6364) );
  OAI21X1 U5948 ( .A(n86), .B(n6365), .C(n6364), .Y(n6368) );
  OAI21X1 U5949 ( .A(n253), .B(n6366), .C(n1074), .Y(n6367) );
  NOR2X1 U5950 ( .A(n5722), .B(n6369), .Y(n6370) );
  AOI21X1 U5951 ( .A(\mem<50><7> ), .B(n5126), .C(n6370), .Y(n6371) );
  AOI22X1 U5952 ( .A(n5215), .B(n470), .C(n5701), .D(n450), .Y(n6373) );
  OAI21X1 U5953 ( .A(n5720), .B(n6376), .C(n4084), .Y(n6380) );
  NAND2X1 U5954 ( .A(\mem<4><7> ), .B(n157), .Y(n6377) );
  OAI21X1 U5955 ( .A(n5734), .B(n6378), .C(n6377), .Y(n6379) );
  NAND2X1 U5956 ( .A(\mem<3><7> ), .B(n198), .Y(n6381) );
  OAI21X1 U5957 ( .A(n5749), .B(n6382), .C(n6381), .Y(n6385) );
  OAI21X1 U5958 ( .A(n5739), .B(n6383), .C(n1076), .Y(n6384) );
  OAI21X1 U5959 ( .A(n5720), .B(n6386), .C(n4086), .Y(n6390) );
  NAND2X1 U5960 ( .A(\mem<44><7> ), .B(n152), .Y(n6387) );
  OAI21X1 U5961 ( .A(n5734), .B(n6388), .C(n6387), .Y(n6389) );
  NAND2X1 U5962 ( .A(\mem<43><7> ), .B(n200), .Y(n6391) );
  OAI21X1 U5963 ( .A(n5749), .B(n6392), .C(n6391), .Y(n6396) );
  NAND2X1 U5964 ( .A(\mem<47><7> ), .B(n227), .Y(n6393) );
  OAI21X1 U5965 ( .A(n5739), .B(n6394), .C(n6393), .Y(n6395) );
  AOI22X1 U5966 ( .A(n33), .B(n1692), .C(n3657), .D(n665), .Y(n6397) );
  AOI21X1 U5967 ( .A(n6398), .B(n1655), .C(n5715), .Y(\data_out<7> ) );
  INVX2 U5968 ( .A(n5715), .Y(n6399) );
  AND2X2 U5969 ( .A(N192), .B(n6399), .Y(\data_out<8> ) );
  AND2X2 U5970 ( .A(N191), .B(n6399), .Y(\data_out<9> ) );
  AND2X2 U5971 ( .A(N189), .B(n6399), .Y(\data_out<11> ) );
  AND2X2 U5972 ( .A(N187), .B(n6399), .Y(\data_out<13> ) );
  AND2X2 U5973 ( .A(N186), .B(n6399), .Y(\data_out<14> ) );
  NAND3X1 U5974 ( .A(enable), .B(wr), .C(n5760), .Y(n6458) );
  NAND3X1 U5975 ( .A(n4255), .B(n1712), .C(n3038), .Y(n6989) );
  NAND3X1 U5976 ( .A(n4257), .B(n1714), .C(n3040), .Y(n6988) );
  NAND3X1 U5977 ( .A(n4259), .B(n1716), .C(n3042), .Y(n6987) );
  NAND3X1 U5978 ( .A(n4261), .B(n1718), .C(n3044), .Y(n6986) );
  NAND3X1 U5979 ( .A(n4263), .B(n1720), .C(n3046), .Y(n6985) );
  NAND3X1 U5980 ( .A(n4265), .B(n1722), .C(n3048), .Y(n6984) );
  NAND3X1 U5981 ( .A(n4267), .B(n1724), .C(n3050), .Y(n6983) );
  NAND3X1 U5982 ( .A(n4269), .B(n1726), .C(n3052), .Y(n6982) );
  AOI21X1 U5983 ( .A(n5735), .B(n218), .C(n5716), .Y(n6450) );
  NAND3X1 U5984 ( .A(n4271), .B(n1728), .C(n3054), .Y(n6981) );
  NAND3X1 U5985 ( .A(n4273), .B(n1730), .C(n3056), .Y(n6980) );
  NAND3X1 U5986 ( .A(n4275), .B(n1732), .C(n3058), .Y(n6979) );
  NAND3X1 U5987 ( .A(n4277), .B(n1734), .C(n3060), .Y(n6978) );
  NAND3X1 U5988 ( .A(n4279), .B(n1736), .C(n3062), .Y(n6977) );
  NAND3X1 U5989 ( .A(n4281), .B(n1738), .C(n3064), .Y(n6976) );
  NAND3X1 U5990 ( .A(n4283), .B(n1740), .C(n3066), .Y(n6975) );
  NAND3X1 U5991 ( .A(n4285), .B(n1742), .C(n3068), .Y(n6974) );
  AOI21X1 U5992 ( .A(n5735), .B(n5740), .C(n5716), .Y(n6451) );
  NAND3X1 U5993 ( .A(n4287), .B(n1744), .C(n3070), .Y(n6973) );
  NAND3X1 U5994 ( .A(n4289), .B(n1746), .C(n3072), .Y(n6972) );
  NAND3X1 U5995 ( .A(n4291), .B(n1748), .C(n3074), .Y(n6971) );
  NAND3X1 U5996 ( .A(n4293), .B(n1750), .C(n3076), .Y(n6970) );
  NAND3X1 U5997 ( .A(n4295), .B(n1752), .C(n3078), .Y(n6969) );
  NAND3X1 U5998 ( .A(n4297), .B(n1754), .C(n3080), .Y(n6968) );
  NAND3X1 U5999 ( .A(n4299), .B(n1756), .C(n3082), .Y(n6967) );
  NAND3X1 U6000 ( .A(n4301), .B(n1758), .C(n3084), .Y(n6966) );
  AOI21X1 U6001 ( .A(n136), .B(n5740), .C(n5716), .Y(n6452) );
  NAND3X1 U6002 ( .A(n4303), .B(n1760), .C(n3086), .Y(n6965) );
  NAND3X1 U6003 ( .A(n4305), .B(n1762), .C(n3088), .Y(n6964) );
  NAND3X1 U6004 ( .A(n4307), .B(n1764), .C(n3090), .Y(n6963) );
  NAND3X1 U6005 ( .A(n4309), .B(n1766), .C(n3092), .Y(n6962) );
  NAND3X1 U6006 ( .A(n4311), .B(n1768), .C(n3094), .Y(n6961) );
  NAND3X1 U6007 ( .A(n4313), .B(n1770), .C(n3096), .Y(n6960) );
  NAND3X1 U6008 ( .A(n4315), .B(n1772), .C(n3098), .Y(n6959) );
  NAND3X1 U6009 ( .A(n4317), .B(n1774), .C(n3100), .Y(n6958) );
  AOI21X1 U6010 ( .A(n120), .B(n176), .C(n5716), .Y(n6453) );
  NAND3X1 U6011 ( .A(n4319), .B(n1776), .C(n3102), .Y(n6957) );
  NAND3X1 U6012 ( .A(n4321), .B(n1778), .C(n3104), .Y(n6956) );
  NAND3X1 U6013 ( .A(n4323), .B(n1780), .C(n3106), .Y(n6955) );
  NAND3X1 U6014 ( .A(n4325), .B(n1782), .C(n3108), .Y(n6954) );
  NAND3X1 U6015 ( .A(n4327), .B(n1784), .C(n3110), .Y(n6953) );
  NAND3X1 U6016 ( .A(n4329), .B(n1786), .C(n3112), .Y(n6952) );
  NAND3X1 U6017 ( .A(n4331), .B(n1788), .C(n3114), .Y(n6951) );
  NAND3X1 U6018 ( .A(n4333), .B(n1790), .C(n3116), .Y(n6950) );
  AOI21X1 U6019 ( .A(n6456), .B(n174), .C(n5716), .Y(n6455) );
  NAND3X1 U6020 ( .A(n4335), .B(n1792), .C(n3118), .Y(n6949) );
  NAND3X1 U6021 ( .A(n4337), .B(n1794), .C(n3120), .Y(n6948) );
  NAND3X1 U6022 ( .A(n4339), .B(n1796), .C(n3122), .Y(n6947) );
  NAND3X1 U6023 ( .A(n4341), .B(n1798), .C(n3124), .Y(n6946) );
  NAND3X1 U6024 ( .A(n4343), .B(n1800), .C(n3126), .Y(n6945) );
  NAND3X1 U6025 ( .A(n4345), .B(n1802), .C(n3128), .Y(n6944) );
  NAND3X1 U6026 ( .A(n4347), .B(n1804), .C(n3130), .Y(n6943) );
  NAND3X1 U6027 ( .A(n4349), .B(n1806), .C(n3132), .Y(n6942) );
  AOI21X1 U6028 ( .A(n5118), .B(n5750), .C(n5716), .Y(n6438) );
  NAND3X1 U6029 ( .A(n4351), .B(n1808), .C(n3134), .Y(n6941) );
  NAND3X1 U6030 ( .A(n4353), .B(n1810), .C(n3136), .Y(n6940) );
  NAND3X1 U6031 ( .A(n4355), .B(n1812), .C(n3138), .Y(n6939) );
  NAND3X1 U6032 ( .A(n4357), .B(n1814), .C(n3140), .Y(n6938) );
  NAND3X1 U6033 ( .A(n4359), .B(n2328), .C(n3142), .Y(n6937) );
  NAND3X1 U6034 ( .A(n4361), .B(n2330), .C(n3144), .Y(n6936) );
  NAND3X1 U6035 ( .A(n4363), .B(n2332), .C(n3146), .Y(n6935) );
  NAND3X1 U6036 ( .A(n4365), .B(n2334), .C(n3148), .Y(n6934) );
  OAI21X1 U6037 ( .A(n6400), .B(n5751), .C(n3666), .Y(n6401) );
  NAND3X1 U6038 ( .A(n272), .B(n2336), .C(n1154), .Y(n6933) );
  NAND3X1 U6039 ( .A(n274), .B(n2338), .C(n1156), .Y(n6932) );
  NAND3X1 U6040 ( .A(n1158), .B(n2340), .C(n3150), .Y(n6931) );
  NAND3X1 U6041 ( .A(n276), .B(n2342), .C(n1160), .Y(n6930) );
  NAND3X1 U6042 ( .A(n278), .B(n2344), .C(n1162), .Y(n6929) );
  NAND3X1 U6043 ( .A(n1164), .B(n2346), .C(n3152), .Y(n6928) );
  NAND3X1 U6044 ( .A(n280), .B(n2348), .C(n1166), .Y(n6927) );
  NAND3X1 U6045 ( .A(n282), .B(n2350), .C(n1168), .Y(n6926) );
  AOI21X1 U6046 ( .A(n5721), .B(n218), .C(n5716), .Y(n6449) );
  NAND3X1 U6047 ( .A(n4367), .B(n2352), .C(n3154), .Y(n6925) );
  NAND3X1 U6048 ( .A(n4369), .B(n2354), .C(n3156), .Y(n6924) );
  NAND3X1 U6049 ( .A(n4371), .B(n2356), .C(n3158), .Y(n6923) );
  NAND3X1 U6050 ( .A(n4373), .B(n2358), .C(n3160), .Y(n6922) );
  NAND3X1 U6051 ( .A(n4375), .B(n2360), .C(n3162), .Y(n6921) );
  NAND3X1 U6052 ( .A(n4377), .B(n2362), .C(n3164), .Y(n6920) );
  NAND3X1 U6053 ( .A(n4379), .B(n2364), .C(n3166), .Y(n6919) );
  NAND3X1 U6054 ( .A(n4381), .B(n2366), .C(n3168), .Y(n6918) );
  NAND3X1 U6055 ( .A(n4383), .B(n2368), .C(n3170), .Y(n6917) );
  NAND3X1 U6056 ( .A(n4385), .B(n2370), .C(n3172), .Y(n6916) );
  NAND3X1 U6057 ( .A(n4387), .B(n2372), .C(n3174), .Y(n6915) );
  NAND3X1 U6058 ( .A(n4389), .B(n2374), .C(n3176), .Y(n6914) );
  NAND3X1 U6059 ( .A(n4391), .B(n2376), .C(n3178), .Y(n6913) );
  NAND3X1 U6060 ( .A(n4393), .B(n2378), .C(n3180), .Y(n6912) );
  NAND3X1 U6061 ( .A(n4395), .B(n2380), .C(n3182), .Y(n6911) );
  NAND3X1 U6062 ( .A(n4397), .B(n2382), .C(n3184), .Y(n6910) );
  NAND3X1 U6063 ( .A(n4399), .B(n2384), .C(n3186), .Y(n6909) );
  NAND3X1 U6064 ( .A(n4401), .B(n2386), .C(n3188), .Y(n6908) );
  NAND3X1 U6065 ( .A(n4403), .B(n2388), .C(n3190), .Y(n6907) );
  NAND3X1 U6066 ( .A(n4405), .B(n2390), .C(n3192), .Y(n6906) );
  NAND3X1 U6067 ( .A(n4407), .B(n2392), .C(n3194), .Y(n6905) );
  NAND3X1 U6068 ( .A(n4409), .B(n2394), .C(n3196), .Y(n6904) );
  NAND3X1 U6069 ( .A(n4411), .B(n2396), .C(n3198), .Y(n6903) );
  NAND3X1 U6070 ( .A(n4413), .B(n2398), .C(n3200), .Y(n6902) );
  NAND3X1 U6071 ( .A(n680), .B(n4415), .C(n1170), .Y(n6901) );
  NAND3X1 U6072 ( .A(n1172), .B(n4417), .C(n682), .Y(n6900) );
  NAND3X1 U6073 ( .A(n1174), .B(n2400), .C(n4419), .Y(n6899) );
  NAND3X1 U6074 ( .A(n1176), .B(n4421), .C(n684), .Y(n6898) );
  NAND3X1 U6075 ( .A(n1178), .B(n4423), .C(n686), .Y(n6897) );
  NAND3X1 U6076 ( .A(n1180), .B(n2402), .C(n4425), .Y(n6896) );
  NAND3X1 U6077 ( .A(n1182), .B(n4427), .C(n688), .Y(n6895) );
  NAND3X1 U6078 ( .A(n1184), .B(n4429), .C(n690), .Y(n6894) );
  NAND3X1 U6079 ( .A(n4431), .B(n2404), .C(n3202), .Y(n6893) );
  NAND3X1 U6080 ( .A(n4433), .B(n2406), .C(n3204), .Y(n6892) );
  NAND3X1 U6081 ( .A(n4435), .B(n2408), .C(n3206), .Y(n6891) );
  NAND3X1 U6082 ( .A(n4437), .B(n2410), .C(n3208), .Y(n6890) );
  NAND3X1 U6083 ( .A(n4439), .B(n2412), .C(n3210), .Y(n6889) );
  NAND3X1 U6084 ( .A(n4441), .B(n2414), .C(n3212), .Y(n6888) );
  NAND3X1 U6085 ( .A(n4443), .B(n2416), .C(n3214), .Y(n6887) );
  NAND3X1 U6086 ( .A(n1186), .B(n2418), .C(n4445), .Y(n6886) );
  NAND3X1 U6087 ( .A(n4447), .B(n2420), .C(n3216), .Y(n6885) );
  NAND3X1 U6088 ( .A(n4449), .B(n2422), .C(n3218), .Y(n6884) );
  NAND3X1 U6089 ( .A(n4451), .B(n2424), .C(n3220), .Y(n6883) );
  NAND3X1 U6090 ( .A(n4453), .B(n2426), .C(n3222), .Y(n6882) );
  NAND3X1 U6091 ( .A(n4455), .B(n2428), .C(n3224), .Y(n6881) );
  NAND3X1 U6092 ( .A(n4457), .B(n2430), .C(n3226), .Y(n6880) );
  NAND3X1 U6093 ( .A(n4459), .B(n2432), .C(n3228), .Y(n6879) );
  NAND3X1 U6094 ( .A(n4461), .B(n2434), .C(n3230), .Y(n6878) );
  NAND3X1 U6095 ( .A(n4463), .B(n2436), .C(n3232), .Y(n6877) );
  NAND3X1 U6096 ( .A(n4465), .B(n2438), .C(n3234), .Y(n6876) );
  NAND3X1 U6097 ( .A(n4467), .B(n2440), .C(n3236), .Y(n6875) );
  NAND3X1 U6098 ( .A(n4469), .B(n2442), .C(n3238), .Y(n6874) );
  NAND3X1 U6099 ( .A(n4471), .B(n2444), .C(n3240), .Y(n6873) );
  NAND3X1 U6100 ( .A(n4473), .B(n2446), .C(n3242), .Y(n6872) );
  NAND3X1 U6101 ( .A(n4475), .B(n2448), .C(n3244), .Y(n6871) );
  NAND3X1 U6102 ( .A(n4477), .B(n2450), .C(n3246), .Y(n6870) );
  NAND3X1 U6103 ( .A(n3768), .B(n2452), .C(n3880), .Y(n6869) );
  NAND3X1 U6104 ( .A(n3770), .B(n2454), .C(n3882), .Y(n6868) );
  NAND3X1 U6105 ( .A(n3772), .B(n2456), .C(n3884), .Y(n6867) );
  NAND3X1 U6106 ( .A(n284), .B(n2458), .C(n3774), .Y(n6866) );
  NAND3X1 U6107 ( .A(n286), .B(n2460), .C(n3776), .Y(n6865) );
  NAND3X1 U6108 ( .A(n288), .B(n2462), .C(n3778), .Y(n6864) );
  NAND3X1 U6109 ( .A(n290), .B(n2464), .C(n3780), .Y(n6863) );
  NAND3X1 U6110 ( .A(n292), .B(n2466), .C(n3782), .Y(n6862) );
  NAND3X1 U6111 ( .A(n1188), .B(n334), .C(n698), .Y(n6861) );
  NAND3X1 U6112 ( .A(n1190), .B(n336), .C(n700), .Y(n6860) );
  NAND3X1 U6113 ( .A(n1192), .B(n338), .C(n702), .Y(n6859) );
  NAND3X1 U6114 ( .A(n1194), .B(n340), .C(n704), .Y(n6858) );
  NAND3X1 U6115 ( .A(n1196), .B(n342), .C(n706), .Y(n6857) );
  NAND3X1 U6116 ( .A(n1198), .B(n344), .C(n708), .Y(n6856) );
  NAND3X1 U6117 ( .A(n1200), .B(n346), .C(n710), .Y(n6855) );
  NAND3X1 U6118 ( .A(n1202), .B(n348), .C(n712), .Y(n6854) );
  NAND3X1 U6119 ( .A(n1204), .B(n350), .C(n3858), .Y(n6853) );
  NAND3X1 U6120 ( .A(n3859), .B(n352), .C(n1206), .Y(n6852) );
  NAND3X1 U6121 ( .A(n1208), .B(n354), .C(n717), .Y(n6851) );
  NAND3X1 U6122 ( .A(n1210), .B(n356), .C(n719), .Y(n6850) );
  NAND3X1 U6123 ( .A(n1212), .B(n358), .C(n721), .Y(n6849) );
  NAND3X1 U6124 ( .A(n1214), .B(n360), .C(n723), .Y(n6848) );
  NAND3X1 U6125 ( .A(n1216), .B(n362), .C(n725), .Y(n6847) );
  NAND3X1 U6126 ( .A(n1218), .B(n364), .C(n727), .Y(n6846) );
  NAND2X1 U6127 ( .A(\mem<45><0> ), .B(n5003), .Y(n6403) );
  NAND3X1 U6128 ( .A(n6403), .B(n1220), .C(n3860), .Y(n6845) );
  NAND2X1 U6129 ( .A(\mem<45><1> ), .B(n5003), .Y(n6404) );
  NAND3X1 U6130 ( .A(n6404), .B(n731), .C(n1222), .Y(n6844) );
  NAND3X1 U6131 ( .A(n3248), .B(n2468), .C(n1224), .Y(n6843) );
  NAND2X1 U6132 ( .A(\mem<45><3> ), .B(n5002), .Y(n6405) );
  NAND3X1 U6133 ( .A(n6405), .B(n1226), .C(n733), .Y(n6842) );
  NAND2X1 U6134 ( .A(\mem<45><4> ), .B(n5002), .Y(n6406) );
  NAND3X1 U6135 ( .A(n6406), .B(n1228), .C(n735), .Y(n6841) );
  NAND3X1 U6136 ( .A(n1230), .B(n2470), .C(n3250), .Y(n6840) );
  NAND2X1 U6137 ( .A(\mem<45><6> ), .B(n5002), .Y(n6407) );
  NAND3X1 U6138 ( .A(n6407), .B(n1232), .C(n737), .Y(n6839) );
  NAND2X1 U6139 ( .A(\mem<45><7> ), .B(n5003), .Y(n6408) );
  NAND3X1 U6140 ( .A(n6408), .B(n1234), .C(n739), .Y(n6838) );
  NAND2X1 U6141 ( .A(\mem<44><0> ), .B(n5005), .Y(n6409) );
  NAND3X1 U6142 ( .A(n6409), .B(n1236), .C(n742), .Y(n6837) );
  NAND2X1 U6143 ( .A(\mem<44><1> ), .B(n5005), .Y(n6410) );
  NAND3X1 U6144 ( .A(n6410), .B(n3861), .C(n1238), .Y(n6836) );
  NAND3X1 U6145 ( .A(n3252), .B(n2472), .C(n1240), .Y(n6835) );
  NAND2X1 U6146 ( .A(\mem<44><3> ), .B(n5004), .Y(n6411) );
  NAND3X1 U6147 ( .A(n6411), .B(n1242), .C(n745), .Y(n6834) );
  NAND2X1 U6148 ( .A(\mem<44><4> ), .B(n5004), .Y(n6412) );
  NAND3X1 U6149 ( .A(n6412), .B(n1244), .C(n747), .Y(n6833) );
  NAND3X1 U6150 ( .A(n1246), .B(n2474), .C(n3254), .Y(n6832) );
  NAND2X1 U6151 ( .A(\mem<44><6> ), .B(n5004), .Y(n6413) );
  NAND3X1 U6152 ( .A(n6413), .B(n1248), .C(n749), .Y(n6831) );
  NAND2X1 U6153 ( .A(\mem<44><7> ), .B(n5005), .Y(n6414) );
  NAND3X1 U6154 ( .A(n6414), .B(n1250), .C(n751), .Y(n6830) );
  NAND2X1 U6155 ( .A(\mem<43><0> ), .B(n5007), .Y(n6415) );
  NAND3X1 U6156 ( .A(n6415), .B(n1252), .C(n754), .Y(n6829) );
  NAND3X1 U6157 ( .A(n1254), .B(n366), .C(n756), .Y(n6828) );
  NAND3X1 U6158 ( .A(n1256), .B(n2476), .C(n3256), .Y(n6827) );
  NAND3X1 U6159 ( .A(n758), .B(n368), .C(n1258), .Y(n6826) );
  NAND3X1 U6160 ( .A(n1260), .B(n370), .C(n760), .Y(n6825) );
  NAND3X1 U6161 ( .A(n1262), .B(n2478), .C(n3258), .Y(n6824) );
  NAND3X1 U6162 ( .A(n1264), .B(n372), .C(n762), .Y(n6823) );
  NAND3X1 U6163 ( .A(n1266), .B(n374), .C(n764), .Y(n6822) );
  NAND2X1 U6164 ( .A(\mem<42><0> ), .B(n5009), .Y(n6416) );
  NAND3X1 U6165 ( .A(n6416), .B(n1268), .C(n3862), .Y(n6821) );
  NAND2X1 U6166 ( .A(\mem<42><1> ), .B(n5009), .Y(n6417) );
  NAND3X1 U6167 ( .A(n6417), .B(n768), .C(n1270), .Y(n6820) );
  NAND3X1 U6168 ( .A(n3260), .B(n2480), .C(n1272), .Y(n6819) );
  NAND2X1 U6169 ( .A(\mem<42><3> ), .B(n5009), .Y(n6418) );
  NAND3X1 U6170 ( .A(n6418), .B(n1274), .C(n770), .Y(n6818) );
  NAND2X1 U6171 ( .A(\mem<42><4> ), .B(n5009), .Y(n6419) );
  NAND3X1 U6172 ( .A(n6419), .B(n1276), .C(n772), .Y(n6817) );
  NAND3X1 U6173 ( .A(n1278), .B(n2482), .C(n3262), .Y(n6816) );
  NAND2X1 U6174 ( .A(\mem<42><6> ), .B(n5009), .Y(n6420) );
  NAND3X1 U6175 ( .A(n6420), .B(n1280), .C(n774), .Y(n6815) );
  NAND2X1 U6176 ( .A(\mem<42><7> ), .B(n5009), .Y(n6421) );
  NAND3X1 U6177 ( .A(n6421), .B(n1282), .C(n776), .Y(n6814) );
  NAND3X1 U6178 ( .A(n294), .B(n3864), .C(n1284), .Y(n6813) );
  NAND3X1 U6179 ( .A(n296), .B(n3866), .C(n1286), .Y(n6812) );
  NAND3X1 U6180 ( .A(n1288), .B(n376), .C(n779), .Y(n6811) );
  NAND3X1 U6181 ( .A(n298), .B(n3868), .C(n1290), .Y(n6810) );
  NAND3X1 U6182 ( .A(n300), .B(n3870), .C(n1292), .Y(n6809) );
  NAND3X1 U6183 ( .A(n781), .B(n378), .C(n1294), .Y(n6808) );
  NAND3X1 U6184 ( .A(n302), .B(n3872), .C(n1296), .Y(n6807) );
  NAND3X1 U6185 ( .A(n304), .B(n3874), .C(n1298), .Y(n6806) );
  OAI21X1 U6186 ( .A(n5751), .B(n6422), .C(n3669), .Y(n6423) );
  NAND3X1 U6187 ( .A(n3784), .B(n2484), .C(n4479), .Y(n6805) );
  NAND3X1 U6188 ( .A(n3786), .B(n2486), .C(n4481), .Y(n6804) );
  NAND3X1 U6189 ( .A(n3788), .B(n2488), .C(n4483), .Y(n6803) );
  NAND3X1 U6190 ( .A(n3790), .B(n2490), .C(n4485), .Y(n6802) );
  NAND3X1 U6191 ( .A(n3792), .B(n2492), .C(n4487), .Y(n6801) );
  NAND3X1 U6192 ( .A(n3794), .B(n2494), .C(n4489), .Y(n6800) );
  NAND3X1 U6193 ( .A(n3796), .B(n2496), .C(n4491), .Y(n6799) );
  NAND3X1 U6194 ( .A(n3798), .B(n2498), .C(n4493), .Y(n6798) );
  NAND3X1 U6195 ( .A(n4495), .B(n787), .C(n785), .Y(n6797) );
  NAND3X1 U6196 ( .A(n4497), .B(n791), .C(n789), .Y(n6796) );
  NAND3X1 U6197 ( .A(n1300), .B(n2500), .C(n3886), .Y(n6795) );
  NAND3X1 U6198 ( .A(n4499), .B(n795), .C(n793), .Y(n6794) );
  NAND3X1 U6199 ( .A(n4501), .B(n799), .C(n797), .Y(n6793) );
  NAND3X1 U6200 ( .A(n1302), .B(n2502), .C(n3888), .Y(n6792) );
  NAND3X1 U6201 ( .A(n4503), .B(n803), .C(n801), .Y(n6791) );
  NAND3X1 U6202 ( .A(n4505), .B(n807), .C(n805), .Y(n6790) );
  NAND3X1 U6203 ( .A(n4507), .B(n2504), .C(n3264), .Y(n6789) );
  NAND3X1 U6204 ( .A(n4509), .B(n2506), .C(n3266), .Y(n6788) );
  NAND3X1 U6205 ( .A(n4511), .B(n2508), .C(n3268), .Y(n6787) );
  NAND3X1 U6206 ( .A(n4513), .B(n2510), .C(n3270), .Y(n6786) );
  NAND3X1 U6207 ( .A(n4515), .B(n2512), .C(n3272), .Y(n6785) );
  NAND3X1 U6208 ( .A(n4517), .B(n2514), .C(n3274), .Y(n6784) );
  NAND3X1 U6209 ( .A(n4519), .B(n2516), .C(n3276), .Y(n6783) );
  NAND3X1 U6210 ( .A(n4521), .B(n2518), .C(n3278), .Y(n6782) );
  NAND3X1 U6211 ( .A(n4523), .B(n2520), .C(n3280), .Y(n6781) );
  NAND3X1 U6212 ( .A(n4525), .B(n2522), .C(n3282), .Y(n6780) );
  NAND3X1 U6213 ( .A(n4527), .B(n2524), .C(n3284), .Y(n6779) );
  NAND3X1 U6214 ( .A(n4529), .B(n2526), .C(n3286), .Y(n6778) );
  NAND3X1 U6215 ( .A(n4531), .B(n2528), .C(n3288), .Y(n6777) );
  NAND3X1 U6216 ( .A(n4533), .B(n2530), .C(n3290), .Y(n6776) );
  NAND3X1 U6217 ( .A(n4535), .B(n2532), .C(n3292), .Y(n6775) );
  NAND3X1 U6218 ( .A(n4537), .B(n2534), .C(n3294), .Y(n6774) );
  NAND3X1 U6219 ( .A(n1304), .B(n2536), .C(n4539), .Y(n6773) );
  NAND3X1 U6220 ( .A(n1306), .B(n2538), .C(n4541), .Y(n6772) );
  NAND3X1 U6221 ( .A(n4543), .B(n2540), .C(n3296), .Y(n6771) );
  NAND3X1 U6222 ( .A(n1308), .B(n2542), .C(n4545), .Y(n6770) );
  NAND3X1 U6223 ( .A(n1310), .B(n2544), .C(n4547), .Y(n6769) );
  NAND3X1 U6224 ( .A(n4549), .B(n2546), .C(n3298), .Y(n6768) );
  NAND3X1 U6225 ( .A(n1312), .B(n2548), .C(n4551), .Y(n6767) );
  NAND3X1 U6226 ( .A(n1314), .B(n2550), .C(n4553), .Y(n6766) );
  NAND3X1 U6227 ( .A(n2552), .B(n1316), .C(n392), .Y(n6765) );
  NAND3X1 U6228 ( .A(n394), .B(n2554), .C(n1318), .Y(n6764) );
  NAND3X1 U6229 ( .A(n3890), .B(n2556), .C(n1320), .Y(n6763) );
  NAND3X1 U6230 ( .A(n1322), .B(n2558), .C(n396), .Y(n6762) );
  NAND3X1 U6231 ( .A(n1324), .B(n2560), .C(n398), .Y(n6761) );
  NAND3X1 U6232 ( .A(n1326), .B(n2562), .C(n3892), .Y(n6760) );
  NAND3X1 U6233 ( .A(n1328), .B(n2564), .C(n400), .Y(n6759) );
  NAND3X1 U6234 ( .A(n1330), .B(n2566), .C(n402), .Y(n6758) );
  NAND3X1 U6235 ( .A(n4039), .B(n380), .C(n1332), .Y(n6757) );
  NAND3X1 U6236 ( .A(n1334), .B(n382), .C(n815), .Y(n6756) );
  NAND3X1 U6237 ( .A(n306), .B(n2568), .C(n1336), .Y(n6755) );
  NAND3X1 U6238 ( .A(n1338), .B(n384), .C(n817), .Y(n6754) );
  NAND3X1 U6239 ( .A(n1340), .B(n386), .C(n819), .Y(n6753) );
  NAND3X1 U6240 ( .A(n308), .B(n2570), .C(n1342), .Y(n6752) );
  NAND3X1 U6241 ( .A(n1344), .B(n388), .C(n821), .Y(n6751) );
  NAND3X1 U6242 ( .A(n1346), .B(n390), .C(n823), .Y(n6750) );
  NAND3X1 U6243 ( .A(n4555), .B(n2572), .C(n3300), .Y(n6749) );
  NAND3X1 U6244 ( .A(n4557), .B(n2574), .C(n3302), .Y(n6748) );
  NAND3X1 U6245 ( .A(n4559), .B(n2576), .C(n3304), .Y(n6747) );
  NAND3X1 U6246 ( .A(n4561), .B(n2578), .C(n3306), .Y(n6746) );
  NAND3X1 U6247 ( .A(n4563), .B(n2580), .C(n3308), .Y(n6745) );
  NAND3X1 U6248 ( .A(n4565), .B(n2582), .C(n3310), .Y(n6744) );
  NAND3X1 U6249 ( .A(n4567), .B(n2584), .C(n3312), .Y(n6743) );
  NAND3X1 U6250 ( .A(n4569), .B(n2586), .C(n3314), .Y(n6742) );
  OAI21X1 U6251 ( .A(n6424), .B(n5750), .C(n3672), .Y(n6425) );
  NAND3X1 U6252 ( .A(n4571), .B(n2588), .C(n3316), .Y(n6741) );
  NAND3X1 U6253 ( .A(n4573), .B(n2590), .C(n3318), .Y(n6740) );
  NAND3X1 U6254 ( .A(n4575), .B(n2592), .C(n3320), .Y(n6739) );
  NAND3X1 U6255 ( .A(n4577), .B(n2594), .C(n3322), .Y(n6738) );
  NAND3X1 U6256 ( .A(n4579), .B(n2596), .C(n3324), .Y(n6737) );
  NAND3X1 U6257 ( .A(n4581), .B(n2598), .C(n3326), .Y(n6736) );
  NAND3X1 U6258 ( .A(n4583), .B(n2600), .C(n3328), .Y(n6735) );
  NAND3X1 U6259 ( .A(n4585), .B(n2602), .C(n1348), .Y(n6734) );
  NAND3X1 U6260 ( .A(n4587), .B(n2604), .C(n3330), .Y(n6733) );
  NAND3X1 U6261 ( .A(n4589), .B(n2606), .C(n3332), .Y(n6732) );
  NAND3X1 U6262 ( .A(n4591), .B(n2608), .C(n3334), .Y(n6731) );
  NAND3X1 U6263 ( .A(n4593), .B(n2610), .C(n3336), .Y(n6730) );
  NAND3X1 U6264 ( .A(n4595), .B(n2612), .C(n3338), .Y(n6729) );
  NAND3X1 U6265 ( .A(n4597), .B(n2614), .C(n3340), .Y(n6728) );
  NAND3X1 U6266 ( .A(n4599), .B(n2616), .C(n3342), .Y(n6727) );
  NAND3X1 U6267 ( .A(n4601), .B(n2618), .C(n3344), .Y(n6726) );
  NAND3X1 U6268 ( .A(n4603), .B(n2620), .C(n3346), .Y(n6725) );
  NAND3X1 U6269 ( .A(n4605), .B(n2622), .C(n3348), .Y(n6724) );
  NAND3X1 U6270 ( .A(n4607), .B(n2624), .C(n3350), .Y(n6723) );
  NAND3X1 U6271 ( .A(n4609), .B(n2626), .C(n3352), .Y(n6722) );
  NAND3X1 U6272 ( .A(n4611), .B(n2628), .C(n3354), .Y(n6721) );
  NAND3X1 U6273 ( .A(n4613), .B(n2630), .C(n3356), .Y(n6720) );
  NAND3X1 U6274 ( .A(n4615), .B(n2632), .C(n3358), .Y(n6719) );
  NAND3X1 U6275 ( .A(n4617), .B(n2634), .C(n3360), .Y(n6718) );
  NAND3X1 U6276 ( .A(n4619), .B(n2636), .C(n3362), .Y(n6717) );
  NAND3X1 U6277 ( .A(n4621), .B(n2638), .C(n3364), .Y(n6716) );
  NAND3X1 U6278 ( .A(n4623), .B(n2640), .C(n3366), .Y(n6715) );
  NAND3X1 U6279 ( .A(n4625), .B(n2642), .C(n3368), .Y(n6714) );
  NAND3X1 U6280 ( .A(n4627), .B(n2644), .C(n3370), .Y(n6713) );
  NAND3X1 U6281 ( .A(n4629), .B(n2646), .C(n3372), .Y(n6712) );
  NAND3X1 U6282 ( .A(n4631), .B(n2648), .C(n3374), .Y(n6711) );
  NAND3X1 U6283 ( .A(n4633), .B(n2650), .C(n3376), .Y(n6710) );
  NAND3X1 U6284 ( .A(n4635), .B(n2652), .C(n3378), .Y(n6709) );
  NAND3X1 U6285 ( .A(n4637), .B(n2654), .C(n3380), .Y(n6708) );
  NAND3X1 U6286 ( .A(n4639), .B(n2656), .C(n3382), .Y(n6707) );
  NAND3X1 U6287 ( .A(n4641), .B(n2658), .C(n3384), .Y(n6706) );
  NAND3X1 U6288 ( .A(n4643), .B(n2660), .C(n3386), .Y(n6705) );
  NAND3X1 U6289 ( .A(n4645), .B(n2662), .C(n3388), .Y(n6704) );
  NAND3X1 U6290 ( .A(n4647), .B(n2664), .C(n3390), .Y(n6703) );
  NAND3X1 U6291 ( .A(n4649), .B(n2666), .C(n3392), .Y(n6702) );
  NAND3X1 U6292 ( .A(n4651), .B(n2668), .C(n3394), .Y(n6701) );
  NAND3X1 U6293 ( .A(n4653), .B(n2670), .C(n3396), .Y(n6700) );
  NAND3X1 U6294 ( .A(n4655), .B(n2672), .C(n3398), .Y(n6699) );
  NAND3X1 U6295 ( .A(n4657), .B(n2674), .C(n3400), .Y(n6698) );
  NAND3X1 U6296 ( .A(n4659), .B(n2676), .C(n3402), .Y(n6697) );
  NAND3X1 U6297 ( .A(n4661), .B(n2678), .C(n3404), .Y(n6696) );
  NAND3X1 U6298 ( .A(n4663), .B(n2680), .C(n3406), .Y(n6695) );
  NAND3X1 U6299 ( .A(n4665), .B(n2682), .C(n3408), .Y(n6694) );
  NAND3X1 U6300 ( .A(n4667), .B(n2684), .C(n3410), .Y(n6693) );
  NAND3X1 U6301 ( .A(n4669), .B(n2686), .C(n3412), .Y(n6692) );
  NAND3X1 U6302 ( .A(n4671), .B(n2688), .C(n3414), .Y(n6691) );
  NAND3X1 U6303 ( .A(n4673), .B(n2690), .C(n3416), .Y(n6690) );
  NAND3X1 U6304 ( .A(n4675), .B(n2692), .C(n3418), .Y(n6689) );
  NAND3X1 U6305 ( .A(n4677), .B(n2694), .C(n3420), .Y(n6688) );
  NAND3X1 U6306 ( .A(n4679), .B(n2696), .C(n3422), .Y(n6687) );
  NAND3X1 U6307 ( .A(n4681), .B(n2698), .C(n3424), .Y(n6686) );
  NAND3X1 U6308 ( .A(n4683), .B(n2700), .C(n3426), .Y(n6685) );
  NAND3X1 U6309 ( .A(n4685), .B(n2702), .C(n3428), .Y(n6684) );
  NAND3X1 U6310 ( .A(n4687), .B(n2704), .C(n3430), .Y(n6683) );
  NAND3X1 U6311 ( .A(n4689), .B(n2706), .C(n3432), .Y(n6682) );
  NAND3X1 U6312 ( .A(n4691), .B(n2708), .C(n3434), .Y(n6681) );
  NAND3X1 U6313 ( .A(n4693), .B(n2710), .C(n3436), .Y(n6680) );
  NAND3X1 U6314 ( .A(n4695), .B(n2712), .C(n3438), .Y(n6679) );
  NAND3X1 U6315 ( .A(n4697), .B(n2714), .C(n3440), .Y(n6678) );
  OAI21X1 U6316 ( .A(n5709), .B(n5750), .C(n70), .Y(n6428) );
  NAND3X1 U6317 ( .A(n3442), .B(n1350), .C(n4699), .Y(n6677) );
  NAND3X1 U6318 ( .A(n1352), .B(n4701), .C(n3444), .Y(n6676) );
  NAND3X1 U6319 ( .A(n1354), .B(n4703), .C(n3446), .Y(n6675) );
  NAND3X1 U6320 ( .A(n1356), .B(n4705), .C(n3448), .Y(n6674) );
  NAND3X1 U6321 ( .A(n1358), .B(n4707), .C(n3450), .Y(n6673) );
  NAND3X1 U6322 ( .A(n1360), .B(n4709), .C(n3452), .Y(n6672) );
  NAND3X1 U6323 ( .A(n1362), .B(n4711), .C(n3454), .Y(n6671) );
  NAND3X1 U6324 ( .A(n1364), .B(n4713), .C(n3456), .Y(n6670) );
  NAND3X1 U6325 ( .A(n4715), .B(n2716), .C(n3458), .Y(n6669) );
  NAND3X1 U6326 ( .A(n4717), .B(n2718), .C(n3460), .Y(n6668) );
  NAND3X1 U6327 ( .A(n4719), .B(n2720), .C(n3462), .Y(n6667) );
  NAND3X1 U6328 ( .A(n4721), .B(n2722), .C(n3464), .Y(n6666) );
  NAND3X1 U6329 ( .A(n4723), .B(n2724), .C(n3466), .Y(n6665) );
  NAND3X1 U6330 ( .A(n4725), .B(n2726), .C(n3468), .Y(n6664) );
  NAND3X1 U6331 ( .A(n4727), .B(n2728), .C(n3470), .Y(n6663) );
  NAND3X1 U6332 ( .A(n4729), .B(n2730), .C(n3472), .Y(n6662) );
  NAND3X1 U6333 ( .A(n4731), .B(n2732), .C(n3474), .Y(n6661) );
  NAND3X1 U6334 ( .A(n4733), .B(n2734), .C(n3476), .Y(n6660) );
  NAND3X1 U6335 ( .A(n4735), .B(n2736), .C(n3478), .Y(n6659) );
  NAND3X1 U6336 ( .A(n4737), .B(n2738), .C(n3480), .Y(n6658) );
  NAND3X1 U6337 ( .A(n4739), .B(n2740), .C(n3482), .Y(n6657) );
  NAND3X1 U6338 ( .A(n4741), .B(n2742), .C(n3484), .Y(n6656) );
  NAND3X1 U6339 ( .A(n4743), .B(n2744), .C(n3486), .Y(n6655) );
  NAND3X1 U6340 ( .A(n4745), .B(n2746), .C(n3488), .Y(n6654) );
  NAND3X1 U6341 ( .A(n4747), .B(n2748), .C(n3490), .Y(n6653) );
  NAND3X1 U6342 ( .A(n4749), .B(n2750), .C(n3492), .Y(n6652) );
  NAND3X1 U6343 ( .A(n4751), .B(n2752), .C(n3494), .Y(n6651) );
  NAND3X1 U6344 ( .A(n4753), .B(n2754), .C(n3496), .Y(n6650) );
  NAND3X1 U6345 ( .A(n4755), .B(n2756), .C(n3498), .Y(n6649) );
  NAND3X1 U6346 ( .A(n4757), .B(n2758), .C(n3500), .Y(n6648) );
  NAND3X1 U6347 ( .A(n4759), .B(n2760), .C(n3502), .Y(n6647) );
  NAND3X1 U6348 ( .A(n4761), .B(n2762), .C(n3504), .Y(n6646) );
  NAND3X1 U6349 ( .A(n4763), .B(n841), .C(n839), .Y(n6645) );
  NAND3X1 U6350 ( .A(n4765), .B(n4040), .C(n843), .Y(n6644) );
  NAND3X1 U6351 ( .A(n4767), .B(n848), .C(n846), .Y(n6643) );
  NAND3X1 U6352 ( .A(n4769), .B(n852), .C(n850), .Y(n6642) );
  NAND3X1 U6353 ( .A(n4771), .B(n856), .C(n854), .Y(n6641) );
  NAND3X1 U6354 ( .A(n4773), .B(n860), .C(n858), .Y(n6640) );
  NAND3X1 U6355 ( .A(n4775), .B(n864), .C(n862), .Y(n6639) );
  NAND3X1 U6356 ( .A(n4777), .B(n868), .C(n866), .Y(n6638) );
  NAND3X1 U6357 ( .A(n4779), .B(n2764), .C(n3506), .Y(n6637) );
  NAND3X1 U6358 ( .A(n4781), .B(n2766), .C(n3508), .Y(n6636) );
  NAND3X1 U6359 ( .A(n4783), .B(n2768), .C(n3510), .Y(n6635) );
  NAND3X1 U6360 ( .A(n4785), .B(n2770), .C(n3512), .Y(n6634) );
  NAND3X1 U6361 ( .A(n4787), .B(n2772), .C(n3514), .Y(n6633) );
  NAND3X1 U6362 ( .A(n4789), .B(n2774), .C(n3516), .Y(n6632) );
  NAND3X1 U6363 ( .A(n4791), .B(n2776), .C(n3518), .Y(n6631) );
  NAND3X1 U6364 ( .A(n4793), .B(n2778), .C(n3520), .Y(n6630) );
  NAND3X1 U6365 ( .A(n4795), .B(n2780), .C(n3522), .Y(n6629) );
  NAND3X1 U6366 ( .A(n4797), .B(n2782), .C(n3524), .Y(n6628) );
  NAND3X1 U6367 ( .A(n4799), .B(n2784), .C(n3526), .Y(n6627) );
  NAND3X1 U6368 ( .A(n4801), .B(n2786), .C(n3528), .Y(n6626) );
  NAND3X1 U6369 ( .A(n4803), .B(n2788), .C(n3530), .Y(n6625) );
  NAND3X1 U6370 ( .A(n4805), .B(n2790), .C(n3532), .Y(n6624) );
  NAND3X1 U6371 ( .A(n4807), .B(n2792), .C(n3534), .Y(n6623) );
  NAND3X1 U6372 ( .A(n4809), .B(n2794), .C(n3536), .Y(n6622) );
  NAND3X1 U6373 ( .A(n4811), .B(n2796), .C(n3538), .Y(n6621) );
  NAND3X1 U6374 ( .A(n4813), .B(n2798), .C(n3540), .Y(n6620) );
  NAND3X1 U6375 ( .A(n4815), .B(n2800), .C(n3542), .Y(n6619) );
  NAND3X1 U6376 ( .A(n4817), .B(n2802), .C(n3544), .Y(n6618) );
  NAND3X1 U6377 ( .A(n4819), .B(n2804), .C(n3546), .Y(n6617) );
  NAND3X1 U6378 ( .A(n4821), .B(n2806), .C(n3548), .Y(n6616) );
  NAND3X1 U6379 ( .A(n4823), .B(n2808), .C(n3550), .Y(n6615) );
  NAND3X1 U6380 ( .A(n4825), .B(n2810), .C(n3552), .Y(n6614) );
  OAI21X1 U6381 ( .A(n30), .B(n5751), .C(n3677), .Y(n6430) );
  NAND2X1 U6382 ( .A(\mem<16><0> ), .B(n5052), .Y(n6431) );
  NAND3X1 U6383 ( .A(n6431), .B(n2812), .C(n3800), .Y(n6613) );
  NAND2X1 U6384 ( .A(\mem<16><1> ), .B(n5052), .Y(n6432) );
  NAND3X1 U6385 ( .A(n6432), .B(n2814), .C(n3802), .Y(n6612) );
  NAND3X1 U6386 ( .A(n1366), .B(n2816), .C(n3804), .Y(n6611) );
  NAND2X1 U6387 ( .A(\mem<16><3> ), .B(n5052), .Y(n6433) );
  NAND3X1 U6388 ( .A(n6433), .B(n2818), .C(n3806), .Y(n6610) );
  NAND2X1 U6389 ( .A(\mem<16><4> ), .B(n5052), .Y(n6434) );
  NAND3X1 U6390 ( .A(n6434), .B(n2820), .C(n3808), .Y(n6609) );
  NAND3X1 U6391 ( .A(n1368), .B(n2822), .C(n3810), .Y(n6608) );
  NAND2X1 U6392 ( .A(\mem<16><6> ), .B(n5052), .Y(n6435) );
  NAND3X1 U6393 ( .A(n6435), .B(n2824), .C(n3812), .Y(n6607) );
  NAND2X1 U6394 ( .A(\mem<16><7> ), .B(n5052), .Y(n6436) );
  NAND3X1 U6395 ( .A(n6436), .B(n2826), .C(n3814), .Y(n6606) );
  NAND3X1 U6396 ( .A(n2828), .B(n1370), .C(n4827), .Y(n6605) );
  NAND3X1 U6397 ( .A(n1372), .B(n2830), .C(n4829), .Y(n6604) );
  NAND3X1 U6398 ( .A(n1374), .B(n2832), .C(n4831), .Y(n6603) );
  NAND3X1 U6399 ( .A(n1376), .B(n2834), .C(n4833), .Y(n6602) );
  NAND3X1 U6400 ( .A(n1378), .B(n2836), .C(n4835), .Y(n6601) );
  NAND3X1 U6401 ( .A(n1380), .B(n2838), .C(n4837), .Y(n6600) );
  NAND3X1 U6402 ( .A(n1382), .B(n2840), .C(n4839), .Y(n6599) );
  NAND3X1 U6403 ( .A(n1384), .B(n2842), .C(n4841), .Y(n6598) );
  NAND3X1 U6404 ( .A(n4843), .B(n2844), .C(n3554), .Y(n6597) );
  NAND3X1 U6405 ( .A(n4845), .B(n2846), .C(n3556), .Y(n6596) );
  NAND3X1 U6406 ( .A(n4847), .B(n2848), .C(n3558), .Y(n6595) );
  NAND3X1 U6407 ( .A(n4849), .B(n2850), .C(n3560), .Y(n6594) );
  NAND3X1 U6408 ( .A(n4851), .B(n2852), .C(n3562), .Y(n6593) );
  NAND3X1 U6409 ( .A(n4853), .B(n2854), .C(n3564), .Y(n6592) );
  NAND3X1 U6410 ( .A(n4855), .B(n2856), .C(n3566), .Y(n6591) );
  NAND3X1 U6411 ( .A(n4857), .B(n2858), .C(n3568), .Y(n6590) );
  NAND3X1 U6412 ( .A(n310), .B(n2908), .C(n1386), .Y(n6565) );
  NAND3X1 U6413 ( .A(n312), .B(n2910), .C(n1388), .Y(n6564) );
  NAND3X1 U6414 ( .A(n314), .B(n2912), .C(n1390), .Y(n6563) );
  NAND3X1 U6415 ( .A(n1392), .B(n2914), .C(n3618), .Y(n6562) );
  NAND3X1 U6416 ( .A(n316), .B(n2916), .C(n1394), .Y(n6561) );
  NAND3X1 U6417 ( .A(n318), .B(n2918), .C(n1396), .Y(n6560) );
  NAND3X1 U6418 ( .A(n320), .B(n2920), .C(n1398), .Y(n6559) );
  NAND3X1 U6419 ( .A(n1400), .B(n2922), .C(n3620), .Y(n6558) );
  OAI21X1 U6420 ( .A(n73), .B(n5751), .C(n3680), .Y(n6440) );
  NAND2X1 U6421 ( .A(\mem<8><0> ), .B(n880), .Y(n6441) );
  NAND3X1 U6422 ( .A(n6441), .B(n1402), .C(n882), .Y(n6549) );
  NAND2X1 U6423 ( .A(\mem<8><1> ), .B(n880), .Y(n6442) );
  NAND3X1 U6424 ( .A(n6442), .B(n1404), .C(n4192), .Y(n6548) );
  NAND2X1 U6425 ( .A(\mem<8><2> ), .B(n880), .Y(n6443) );
  NAND3X1 U6426 ( .A(n6443), .B(n1406), .C(n885), .Y(n6547) );
  NAND2X1 U6427 ( .A(\mem<8><3> ), .B(n880), .Y(n6444) );
  NAND3X1 U6428 ( .A(n6444), .B(n1408), .C(n887), .Y(n6546) );
  NAND2X1 U6429 ( .A(\mem<8><4> ), .B(n880), .Y(n6445) );
  NAND3X1 U6430 ( .A(n6445), .B(n1410), .C(n889), .Y(n6545) );
  NAND2X1 U6431 ( .A(\mem<8><5> ), .B(n880), .Y(n6446) );
  NAND3X1 U6432 ( .A(n6446), .B(n1412), .C(n891), .Y(n6544) );
  NAND2X1 U6433 ( .A(\mem<8><6> ), .B(n880), .Y(n6447) );
  NAND3X1 U6434 ( .A(n6447), .B(n1414), .C(n893), .Y(n6543) );
  NAND2X1 U6435 ( .A(\mem<8><7> ), .B(n880), .Y(n6448) );
  NAND3X1 U6436 ( .A(n6448), .B(n1416), .C(n895), .Y(n6542) );
  NAND3X1 U6437 ( .A(n1418), .B(n4859), .C(n3894), .Y(n6541) );
  NAND3X1 U6438 ( .A(n1420), .B(n4861), .C(n3896), .Y(n6540) );
  NAND3X1 U6439 ( .A(n1422), .B(n4863), .C(n3898), .Y(n6539) );
  NAND3X1 U6440 ( .A(n1424), .B(n4865), .C(n3900), .Y(n6538) );
  NAND3X1 U6441 ( .A(n1426), .B(n4867), .C(n3902), .Y(n6537) );
  NAND3X1 U6442 ( .A(n1428), .B(n4869), .C(n3904), .Y(n6536) );
  NAND3X1 U6443 ( .A(n1430), .B(n4871), .C(n3906), .Y(n6535) );
  NAND3X1 U6444 ( .A(n1432), .B(n4873), .C(n3908), .Y(n6534) );
  NAND3X1 U6445 ( .A(n1434), .B(n2940), .C(n4875), .Y(n6533) );
  NAND3X1 U6446 ( .A(n1436), .B(n2942), .C(n4877), .Y(n6532) );
  NAND3X1 U6447 ( .A(n1438), .B(n2944), .C(n4879), .Y(n6531) );
  NAND3X1 U6448 ( .A(n1440), .B(n2946), .C(n4881), .Y(n6530) );
  NAND3X1 U6449 ( .A(n1442), .B(n2948), .C(n4883), .Y(n6529) );
  NAND3X1 U6450 ( .A(n1444), .B(n2950), .C(n4885), .Y(n6528) );
  NAND3X1 U6451 ( .A(n1446), .B(n2952), .C(n4887), .Y(n6527) );
  NAND3X1 U6452 ( .A(n1448), .B(n2954), .C(n4889), .Y(n6526) );
  NAND3X1 U6453 ( .A(n322), .B(n2956), .C(n1450), .Y(n6525) );
  NAND3X1 U6454 ( .A(n324), .B(n2958), .C(n1452), .Y(n6524) );
  NAND3X1 U6455 ( .A(n1454), .B(n2960), .C(n3638), .Y(n6523) );
  NAND3X1 U6456 ( .A(n326), .B(n2962), .C(n1456), .Y(n6522) );
  NAND3X1 U6457 ( .A(n328), .B(n2964), .C(n1458), .Y(n6521) );
  NAND3X1 U6458 ( .A(n1460), .B(n2966), .C(n3640), .Y(n6520) );
  NAND3X1 U6459 ( .A(n330), .B(n2968), .C(n1462), .Y(n6519) );
  NAND3X1 U6460 ( .A(n332), .B(n2970), .C(n1464), .Y(n6518) );
  NAND3X1 U6461 ( .A(n1466), .B(n2972), .C(n4891), .Y(n6517) );
  NAND3X1 U6462 ( .A(n1468), .B(n2974), .C(n4893), .Y(n6516) );
  NAND3X1 U6463 ( .A(n4895), .B(n1470), .C(n3642), .Y(n6515) );
  NAND3X1 U6464 ( .A(n1472), .B(n2976), .C(n4897), .Y(n6514) );
  NAND3X1 U6465 ( .A(n1474), .B(n2978), .C(n4899), .Y(n6513) );
  NAND3X1 U6466 ( .A(n1476), .B(n4901), .C(n3644), .Y(n6512) );
  NAND3X1 U6467 ( .A(n1478), .B(n2980), .C(n4903), .Y(n6511) );
  NAND3X1 U6468 ( .A(n1480), .B(n2982), .C(n4905), .Y(n6510) );
  NAND3X1 U6469 ( .A(n1482), .B(n2984), .C(n4907), .Y(n6509) );
  NAND3X1 U6470 ( .A(n1484), .B(n2986), .C(n4909), .Y(n6508) );
  NAND3X1 U6471 ( .A(n1486), .B(n2988), .C(n4911), .Y(n6507) );
  NAND3X1 U6472 ( .A(n1488), .B(n2990), .C(n4913), .Y(n6506) );
  NAND3X1 U6473 ( .A(n1490), .B(n2992), .C(n4915), .Y(n6505) );
  NAND3X1 U6474 ( .A(n1492), .B(n2994), .C(n4917), .Y(n6504) );
  NAND3X1 U6475 ( .A(n4919), .B(n1494), .C(n3646), .Y(n6503) );
  NAND3X1 U6476 ( .A(n1496), .B(n4921), .C(n3648), .Y(n6502) );
  NAND3X1 U6477 ( .A(n1498), .B(n2996), .C(n4923), .Y(n6501) );
  NAND3X1 U6478 ( .A(n1500), .B(n2998), .C(n4925), .Y(n6500) );
  NAND3X1 U6479 ( .A(n4927), .B(n1502), .C(n3650), .Y(n6499) );
  NAND3X1 U6480 ( .A(n1504), .B(n3000), .C(n4929), .Y(n6498) );
  NAND3X1 U6481 ( .A(n1506), .B(n3002), .C(n4931), .Y(n6497) );
  NAND3X1 U6482 ( .A(n1508), .B(n4933), .C(n3652), .Y(n6496) );
  NAND3X1 U6483 ( .A(n1510), .B(n3004), .C(n4935), .Y(n6495) );
  NAND3X1 U6484 ( .A(n1512), .B(n3006), .C(n4937), .Y(n6494) );
  INVX2 U6485 ( .A(n3968), .Y(n6460) );
  NAND3X1 U6486 ( .A(n1514), .B(n4236), .C(n4194), .Y(n6493) );
  NAND3X1 U6487 ( .A(n1516), .B(n4238), .C(n4196), .Y(n6492) );
  NAND3X1 U6488 ( .A(n1518), .B(n4240), .C(n4198), .Y(n6491) );
  NAND3X1 U6489 ( .A(n1520), .B(n4242), .C(n4200), .Y(n6490) );
  NAND3X1 U6490 ( .A(n1522), .B(n4244), .C(n4202), .Y(n6489) );
  NAND3X1 U6491 ( .A(n1524), .B(n4246), .C(n4204), .Y(n6488) );
  NAND3X1 U6492 ( .A(n1526), .B(n4248), .C(n4206), .Y(n6487) );
  NAND3X1 U6493 ( .A(n1528), .B(n4250), .C(n4208), .Y(n6486) );
  MUX2X1 U6494 ( .B(n6464), .A(n6463), .S(n47), .Y(n6484) );
  MUX2X1 U6495 ( .B(n6466), .A(n6465), .S(n47), .Y(n6483) );
  MUX2X1 U6496 ( .B(n6468), .A(n6467), .S(n47), .Y(n6482) );
  MUX2X1 U6497 ( .B(n6470), .A(n6469), .S(n47), .Y(n6481) );
  MUX2X1 U6498 ( .B(n6472), .A(n6471), .S(n50), .Y(n6480) );
  MUX2X1 U6499 ( .B(n6476), .A(n6475), .S(n50), .Y(n6478) );
endmodule


module fetch ( clk, rst, halt, .nextPC({\nextPC<15> , \nextPC<14> , 
        \nextPC<13> , \nextPC<12> , \nextPC<11> , \nextPC<10> , \nextPC<9> , 
        \nextPC<8> , \nextPC<7> , \nextPC<6> , \nextPC<5> , \nextPC<4> , 
        \nextPC<3> , \nextPC<2> , \nextPC<1> , \nextPC<0> }), .PC2({\PC2<15> , 
        \PC2<14> , \PC2<13> , \PC2<12> , \PC2<11> , \PC2<10> , \PC2<9> , 
        \PC2<8> , \PC2<7> , \PC2<6> , \PC2<5> , \PC2<4> , \PC2<3> , \PC2<2> , 
        \PC2<1> , \PC2<0> }), .instr({\instr<15> , \instr<14> , \instr<13> , 
        \instr<12> , \instr<11> , \instr<10> , \instr<9> , \instr<8> , 
        \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> , \instr<2> , 
        \instr<1> , \instr<0> }), err );
  input clk, rst, halt, \nextPC<15> , \nextPC<14> , \nextPC<13> , \nextPC<12> ,
         \nextPC<11> , \nextPC<10> , \nextPC<9> , \nextPC<8> , \nextPC<7> ,
         \nextPC<6> , \nextPC<5> , \nextPC<4> , \nextPC<3> , \nextPC<2> ,
         \nextPC<1> , \nextPC<0> ;
  output \PC2<15> , \PC2<14> , \PC2<13> , \PC2<12> , \PC2<11> , \PC2<10> ,
         \PC2<9> , \PC2<8> , \PC2<7> , \PC2<6> , \PC2<5> , \PC2<4> , \PC2<3> ,
         \PC2<2> , \PC2<1> , \PC2<0> , \instr<15> , \instr<14> , \instr<13> ,
         \instr<12> , \instr<11> , \instr<10> , \instr<9> , \instr<8> ,
         \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> ,
         \instr<2> , \instr<1> , \instr<0> , err;
  wire   \currentPC<15> , \currentPC<14> , \currentPC<13> , \currentPC<12> ,
         \currentPC<11> , \currentPC<10> , \currentPC<9> , \currentPC<8> ,
         \currentPC<7> , \currentPC<6> , \currentPC<5> , \currentPC<4> ,
         \currentPC<3> , \currentPC<2> , \currentPC<1> , \currentPC<0> , n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18;
  assign err = 1'b0;

  dff_128 \pc[0]  ( .q(\currentPC<0> ), .d(\nextPC<0> ), .clk(clk), .rst(n17)
         );
  dff_129 \pc[1]  ( .q(\currentPC<1> ), .d(\nextPC<1> ), .clk(clk), .rst(n17)
         );
  dff_130 \pc[2]  ( .q(\currentPC<2> ), .d(\nextPC<2> ), .clk(clk), .rst(rst)
         );
  dff_131 \pc[3]  ( .q(\currentPC<3> ), .d(\nextPC<3> ), .clk(clk), .rst(rst)
         );
  dff_132 \pc[4]  ( .q(\currentPC<4> ), .d(\nextPC<4> ), .clk(clk), .rst(rst)
         );
  dff_133 \pc[5]  ( .q(\currentPC<5> ), .d(\nextPC<5> ), .clk(clk), .rst(rst)
         );
  dff_134 \pc[6]  ( .q(\currentPC<6> ), .d(\nextPC<6> ), .clk(clk), .rst(n17)
         );
  dff_135 \pc[7]  ( .q(\currentPC<7> ), .d(\nextPC<7> ), .clk(clk), .rst(n17)
         );
  dff_136 \pc[8]  ( .q(\currentPC<8> ), .d(\nextPC<8> ), .clk(clk), .rst(n17)
         );
  dff_137 \pc[9]  ( .q(\currentPC<9> ), .d(\nextPC<9> ), .clk(clk), .rst(n17)
         );
  dff_138 \pc[10]  ( .q(\currentPC<10> ), .d(\nextPC<10> ), .clk(clk), .rst(
        n17) );
  dff_139 \pc[11]  ( .q(\currentPC<11> ), .d(\nextPC<11> ), .clk(clk), .rst(
        n17) );
  dff_140 \pc[12]  ( .q(\currentPC<12> ), .d(\nextPC<12> ), .clk(clk), .rst(
        n17) );
  dff_141 \pc[13]  ( .q(\currentPC<13> ), .d(\nextPC<13> ), .clk(clk), .rst(
        n17) );
  dff_142 \pc[14]  ( .q(\currentPC<14> ), .d(\nextPC<14> ), .clk(clk), .rst(
        n17) );
  dff_143 \pc[15]  ( .q(\currentPC<15> ), .d(\nextPC<15> ), .clk(clk), .rst(
        n17) );
  memory2c_1 instrmem ( .data_out({\instr<15> , \instr<14> , \instr<13> , 
        \instr<12> , \instr<11> , \instr<10> , \instr<9> , \instr<8> , 
        \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> , \instr<2> , 
        \instr<1> , \instr<0> }), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .addr({
        \currentPC<15> , \currentPC<14> , \currentPC<13> , \currentPC<12> , 
        \currentPC<11> , \currentPC<10> , \currentPC<9> , \currentPC<8> , 
        \currentPC<7> , \currentPC<6> , n6, n13, \currentPC<3> , 
        \currentPC<2> , \currentPC<1> , \currentPC<0> }), .enable(1'b1), .wr(
        1'b0), .createdump(1'b0), .clk(clk), .rst(n17) );
  adder_2 pcAdd ( .A({n11, n10, n4, \currentPC<12> , \currentPC<11> , 
        \currentPC<10> , n14, \currentPC<8> , \currentPC<7> , \currentPC<6> , 
        n3, n13, n9, n8, n16, n7}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0}), .Cin(
        1'b0), .Overflow(), .Cout(), .Sum({\PC2<15> , \PC2<14> , \PC2<13> , 
        \PC2<12> , \PC2<11> , \PC2<10> , \PC2<9> , \PC2<8> , \PC2<7> , 
        \PC2<6> , \PC2<5> , \PC2<4> , \PC2<3> , \PC2<2> , \PC2<1> , \PC2<0> })
         );
  INVX1 U4 ( .A(n18), .Y(n17) );
  INVX1 U5 ( .A(rst), .Y(n18) );
  INVX1 U6 ( .A(n6), .Y(n2) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  BUFX2 U8 ( .A(\currentPC<13> ), .Y(n4) );
  INVX4 U9 ( .A(\currentPC<5> ), .Y(n5) );
  INVX8 U10 ( .A(n5), .Y(n6) );
  BUFX2 U11 ( .A(\currentPC<0> ), .Y(n7) );
  BUFX2 U12 ( .A(\currentPC<2> ), .Y(n8) );
  BUFX2 U13 ( .A(\currentPC<3> ), .Y(n9) );
  BUFX2 U14 ( .A(\currentPC<14> ), .Y(n10) );
  BUFX2 U15 ( .A(\currentPC<15> ), .Y(n11) );
  INVX4 U16 ( .A(\currentPC<4> ), .Y(n12) );
  INVX8 U17 ( .A(n12), .Y(n13) );
  BUFX2 U18 ( .A(\currentPC<9> ), .Y(n14) );
  INVX1 U19 ( .A(\currentPC<1> ), .Y(n15) );
  INVX1 U20 ( .A(n15), .Y(n16) );
endmodule


module decode ( clk, rst, .instr({\instr<15> , \instr<14> , \instr<13> , 
        \instr<12> , \instr<11> , \instr<10> , \instr<9> , \instr<8> , 
        \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> , \instr<2> , 
        \instr<1> , \instr<0> }), .PC({\PC<15> , \PC<14> , \PC<13> , \PC<12> , 
        \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> , 
        \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> }), .writeBackData({
        \writeBackData<15> , \writeBackData<14> , \writeBackData<13> , 
        \writeBackData<12> , \writeBackData<11> , \writeBackData<10> , 
        \writeBackData<9> , \writeBackData<8> , \writeBackData<7> , 
        \writeBackData<6> , \writeBackData<5> , \writeBackData<4> , 
        \writeBackData<3> , \writeBackData<2> , \writeBackData<1> , 
        \writeBackData<0> }), .readdata1({\readdata1<15> , \readdata1<14> , 
        \readdata1<13> , \readdata1<12> , \readdata1<11> , \readdata1<10> , 
        \readdata1<9> , \readdata1<8> , \readdata1<7> , \readdata1<6> , 
        \readdata1<5> , \readdata1<4> , \readdata1<3> , \readdata1<2> , 
        \readdata1<1> , \readdata1<0> }), .readdata2({\readdata2<15> , 
        \readdata2<14> , \readdata2<13> , \readdata2<12> , \readdata2<11> , 
        \readdata2<10> , \readdata2<9> , \readdata2<8> , \readdata2<7> , 
        \readdata2<6> , \readdata2<5> , \readdata2<4> , \readdata2<3> , 
        \readdata2<2> , \readdata2<1> , \readdata2<0> }), .immediate({
        \immediate<15> , \immediate<14> , \immediate<13> , \immediate<12> , 
        \immediate<11> , \immediate<10> , \immediate<9> , \immediate<8> , 
        \immediate<7> , \immediate<6> , \immediate<5> , \immediate<4> , 
        \immediate<3> , \immediate<2> , \immediate<1> , \immediate<0> }), jump, 
        jumpReg, branch, .branchOp({\branchOp<1> , \branchOp<0> }), memRead, 
        memWrite, memToReg, .ALUOp({\ALUOp<3> , \ALUOp<2> , \ALUOp<1> , 
        \ALUOp<0> }), ALUSrc, invSrc1, invSrc2, sub, halt, passthrough, 
        reverse, err );
  input clk, rst, \instr<15> , \instr<14> , \instr<13> , \instr<12> ,
         \instr<11> , \instr<10> , \instr<9> , \instr<8> , \instr<7> ,
         \instr<6> , \instr<5> , \instr<4> , \instr<3> , \instr<2> ,
         \instr<1> , \instr<0> , \PC<15> , \PC<14> , \PC<13> , \PC<12> ,
         \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> ,
         \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> , \writeBackData<15> ,
         \writeBackData<14> , \writeBackData<13> , \writeBackData<12> ,
         \writeBackData<11> , \writeBackData<10> , \writeBackData<9> ,
         \writeBackData<8> , \writeBackData<7> , \writeBackData<6> ,
         \writeBackData<5> , \writeBackData<4> , \writeBackData<3> ,
         \writeBackData<2> , \writeBackData<1> , \writeBackData<0> ;
  output \readdata1<15> , \readdata1<14> , \readdata1<13> , \readdata1<12> ,
         \readdata1<11> , \readdata1<10> , \readdata1<9> , \readdata1<8> ,
         \readdata1<7> , \readdata1<6> , \readdata1<5> , \readdata1<4> ,
         \readdata1<3> , \readdata1<2> , \readdata1<1> , \readdata1<0> ,
         \readdata2<15> , \readdata2<14> , \readdata2<13> , \readdata2<12> ,
         \readdata2<11> , \readdata2<10> , \readdata2<9> , \readdata2<8> ,
         \readdata2<7> , \readdata2<6> , \readdata2<5> , \readdata2<4> ,
         \readdata2<3> , \readdata2<2> , \readdata2<1> , \readdata2<0> ,
         \immediate<15> , \immediate<14> , \immediate<13> , \immediate<12> ,
         \immediate<11> , \immediate<10> , \immediate<9> , \immediate<8> ,
         \immediate<7> , \immediate<6> , \immediate<5> , \immediate<4> ,
         \immediate<3> , \immediate<2> , \immediate<1> , \immediate<0> , jump,
         jumpReg, branch, \branchOp<1> , \branchOp<0> , memRead, memWrite,
         memToReg, \ALUOp<3> , \ALUOp<2> , \ALUOp<1> , \ALUOp<0> , ALUSrc,
         invSrc1, invSrc2, sub, halt, passthrough, reverse, err;
  wire   n138, \regDst<1> , \regDst<0> , \writereg<2> , \writereg<1> ,
         \writereg<0> , \whichImm<1> , \whichImm<0> , toExt, regWrite, n28,
         n29, n32, n34, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n30,
         n31, n33, n35, n36, n37, n39, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n83, n85, n87, n88, n90, n91, n92, n93, n95,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n129, n130, n131, n132, n133, n134, n135,
         n136;
  assign \readdata1<15>  = 1'b0;
  assign \readdata1<14>  = 1'b0;
  assign \readdata1<13>  = 1'b0;
  assign \readdata1<12>  = 1'b0;
  assign \readdata1<11>  = 1'b0;
  assign \readdata1<10>  = 1'b0;
  assign \readdata1<9>  = 1'b0;
  assign \readdata1<8>  = 1'b0;
  assign \readdata1<7>  = 1'b0;
  assign \readdata1<6>  = 1'b0;
  assign \readdata1<5>  = 1'b0;
  assign \readdata1<4>  = 1'b0;
  assign \readdata1<3>  = 1'b0;
  assign \readdata1<2>  = 1'b0;
  assign \readdata1<1>  = 1'b0;
  assign \readdata1<0>  = 1'b0;
  assign \readdata2<15>  = 1'b0;
  assign \readdata2<14>  = 1'b0;
  assign \readdata2<13>  = 1'b0;
  assign \readdata2<12>  = 1'b0;
  assign \readdata2<11>  = 1'b0;
  assign \readdata2<10>  = 1'b0;
  assign \readdata2<9>  = 1'b0;
  assign \readdata2<8>  = 1'b0;
  assign \readdata2<7>  = 1'b0;
  assign \readdata2<6>  = 1'b0;
  assign \readdata2<5>  = 1'b0;
  assign \readdata2<4>  = 1'b0;
  assign \readdata2<3>  = 1'b0;
  assign \readdata2<2>  = 1'b0;
  assign \readdata2<1>  = 1'b0;
  assign \readdata2<0>  = 1'b0;
  assign err = 1'b0;

  NAND3X1 U30 ( .A(n65), .B(n102), .C(n68), .Y(\writereg<2> ) );
  AOI22X1 U31 ( .A(\immediate<4> ), .B(n126), .C(n48), .D(\regDst<0> ), .Y(n29) );
  NAND3X1 U33 ( .A(n63), .B(n101), .C(n67), .Y(\writereg<1> ) );
  AOI22X1 U34 ( .A(\immediate<3> ), .B(n126), .C(n47), .D(\regDst<0> ), .Y(n32) );
  NAND3X1 U36 ( .A(n61), .B(n101), .C(n66), .Y(\writereg<0> ) );
  AOI22X1 U37 ( .A(\immediate<2> ), .B(n126), .C(n46), .D(\regDst<0> ), .Y(n34) );
  control ctrl ( .instr({\instr<15> , \instr<14> , \instr<13> , \instr<12> , 
        \instr<11> }), .func({n5, n31}), .regDst({\regDst<1> , \regDst<0> }), 
        .regWrite(regWrite), .whichImm({\whichImm<1> , \whichImm<0> }), 
        .toExt(toExt), .jump(jump), .jumpReg(jumpReg), .branch(branch), 
        .branchOp({\branchOp<1> , \branchOp<0> }), .memRead(memRead), 
        .memWrite(memWrite), .memToReg(memToReg), .ALUOp({\ALUOp<3> , 
        \ALUOp<2> , \ALUOp<1> , \ALUOp<0> }), .ALUSrc(ALUSrc), .invSrc1(
        invSrc1), .invSrc2(n138), .sub(sub), .halt(halt), .passthrough(
        passthrough), .reverse(reverse), .err() );
  rf register ( .read1data(), .read2data(), .err(), .clk(clk), .rst(rst), 
        .read1regsel({\instr<10> , \instr<9> , \instr<8> }), .read2regsel({
        \instr<7> , \instr<6> , \instr<5> }), .writeregsel({\writereg<2> , 
        \writereg<1> , \writereg<0> }), .writedata({n129, n130, n131, n132, 
        n133, n134, n135, n136, n54, n51, n10, n77, n16, n7, n19, n13}), 
        .write(regWrite) );
  INVX1 U3 ( .A(\PC<0> ), .Y(n14) );
  INVX1 U4 ( .A(\PC<11> ), .Y(n110) );
  INVX1 U5 ( .A(\instr<8> ), .Y(n123) );
  INVX1 U6 ( .A(\PC<6> ), .Y(n52) );
  INVX1 U7 ( .A(\PC<1> ), .Y(n20) );
  INVX1 U8 ( .A(\PC<3> ), .Y(n17) );
  INVX1 U9 ( .A(\PC<9> ), .Y(n106) );
  INVX1 U10 ( .A(\PC<12> ), .Y(n112) );
  INVX1 U11 ( .A(\PC<2> ), .Y(n8) );
  INVX1 U12 ( .A(\PC<15> ), .Y(n118) );
  INVX1 U13 ( .A(\PC<5> ), .Y(n11) );
  INVX1 U14 ( .A(\PC<7> ), .Y(n55) );
  INVX1 U15 ( .A(\PC<8> ), .Y(n104) );
  INVX1 U16 ( .A(\PC<10> ), .Y(n108) );
  INVX1 U17 ( .A(\PC<13> ), .Y(n114) );
  INVX1 U18 ( .A(\PC<14> ), .Y(n116) );
  BUFX2 U19 ( .A(n28), .Y(n101) );
  INVX1 U20 ( .A(n28), .Y(n2) );
  INVX1 U21 ( .A(n28), .Y(n1) );
  INVX1 U22 ( .A(n28), .Y(n3) );
  MUX2X1 U23 ( .B(n9), .A(n8), .S(n1), .Y(n7) );
  MUX2X1 U24 ( .B(n15), .A(n14), .S(n2), .Y(n13) );
  MUX2X1 U25 ( .B(n56), .A(n55), .S(n3), .Y(n54) );
  MUX2X1 U26 ( .B(n53), .A(n52), .S(n6), .Y(n51) );
  BUFX2 U27 ( .A(n93), .Y(n4) );
  MUX2X1 U28 ( .B(n12), .A(n11), .S(n6), .Y(n10) );
  INVX1 U29 ( .A(n28), .Y(n6) );
  INVX1 U32 ( .A(n93), .Y(n5) );
  MUX2X1 U35 ( .B(n21), .A(n20), .S(n6), .Y(n19) );
  INVX1 U38 ( .A(\writeBackData<2> ), .Y(n9) );
  MUX2X1 U39 ( .B(n18), .A(n17), .S(n1), .Y(n16) );
  INVX1 U40 ( .A(\writeBackData<5> ), .Y(n12) );
  INVX1 U41 ( .A(\writeBackData<0> ), .Y(n15) );
  INVX1 U42 ( .A(\writeBackData<3> ), .Y(n18) );
  INVX1 U43 ( .A(\writeBackData<1> ), .Y(n21) );
  AND2X2 U44 ( .A(n27), .B(n44), .Y(n22) );
  INVX1 U45 ( .A(n22), .Y(\immediate<5> ) );
  OR2X2 U46 ( .A(n80), .B(\whichImm<1> ), .Y(n24) );
  INVX1 U47 ( .A(n24), .Y(n25) );
  AND2X2 U48 ( .A(n87), .B(n57), .Y(n26) );
  INVX1 U49 ( .A(n26), .Y(n27) );
  BUFX2 U50 ( .A(\regDst<1> ), .Y(n30) );
  BUFX2 U51 ( .A(\instr<0> ), .Y(n31) );
  AND2X2 U52 ( .A(\instr<10> ), .B(n25), .Y(n33) );
  INVX1 U53 ( .A(n33), .Y(n35) );
  INVX1 U54 ( .A(n33), .Y(n36) );
  BUFX2 U55 ( .A(\instr<4> ), .Y(n37) );
  BUFX2 U56 ( .A(n138), .Y(invSrc2) );
  AND2X2 U57 ( .A(n42), .B(n35), .Y(n39) );
  INVX1 U58 ( .A(n39), .Y(\immediate<13> ) );
  INVX1 U59 ( .A(n39), .Y(n41) );
  BUFX2 U60 ( .A(n125), .Y(n42) );
  AND2X2 U61 ( .A(n50), .B(n90), .Y(n43) );
  INVX1 U62 ( .A(n43), .Y(n44) );
  INVX1 U63 ( .A(n43), .Y(n45) );
  INVX1 U64 ( .A(n120), .Y(n46) );
  INVX1 U65 ( .A(n121), .Y(n47) );
  INVX1 U66 ( .A(n122), .Y(n48) );
  INVX1 U67 ( .A(n122), .Y(n49) );
  INVX1 U68 ( .A(\instr<7> ), .Y(n122) );
  INVX1 U69 ( .A(n91), .Y(n50) );
  INVX1 U70 ( .A(\writeBackData<6> ), .Y(n53) );
  INVX1 U71 ( .A(\writeBackData<7> ), .Y(n56) );
  BUFX2 U72 ( .A(n41), .Y(\immediate<15> ) );
  INVX2 U73 ( .A(n83), .Y(\immediate<3> ) );
  INVX1 U74 ( .A(\whichImm<0> ), .Y(n57) );
  INVX1 U75 ( .A(\instr<3> ), .Y(n83) );
  BUFX2 U76 ( .A(n28), .Y(n102) );
  AND2X2 U77 ( .A(\PC<4> ), .B(n3), .Y(n58) );
  INVX1 U78 ( .A(n58), .Y(n59) );
  AND2X2 U79 ( .A(\instr<8> ), .B(n71), .Y(n60) );
  INVX1 U80 ( .A(n60), .Y(n61) );
  AND2X2 U81 ( .A(\instr<9> ), .B(n72), .Y(n62) );
  INVX1 U82 ( .A(n62), .Y(n63) );
  AND2X2 U83 ( .A(\instr<10> ), .B(n70), .Y(n64) );
  INVX1 U84 ( .A(n64), .Y(n65) );
  INVX1 U85 ( .A(\instr<2> ), .Y(n81) );
  BUFX2 U86 ( .A(n34), .Y(n66) );
  BUFX2 U87 ( .A(n32), .Y(n67) );
  BUFX2 U88 ( .A(n29), .Y(n68) );
  INVX1 U89 ( .A(\instr<6> ), .Y(n121) );
  OR2X2 U90 ( .A(n126), .B(\regDst<0> ), .Y(n69) );
  INVX1 U91 ( .A(n69), .Y(n70) );
  INVX1 U92 ( .A(n69), .Y(n71) );
  INVX1 U93 ( .A(n69), .Y(n72) );
  AOI21X1 U94 ( .A(\instr<9> ), .B(n73), .C(n76), .Y(n74) );
  INVX1 U95 ( .A(n124), .Y(n73) );
  INVX1 U96 ( .A(n74), .Y(\immediate<9> ) );
  OAI21X1 U97 ( .A(n75), .B(n3), .C(n59), .Y(n77) );
  INVX1 U98 ( .A(\writeBackData<4> ), .Y(n75) );
  INVX1 U99 ( .A(n42), .Y(n76) );
  INVX1 U100 ( .A(n95), .Y(\immediate<11> ) );
  INVX1 U101 ( .A(n124), .Y(n78) );
  INVX1 U102 ( .A(n78), .Y(n79) );
  INVX1 U103 ( .A(n91), .Y(n80) );
  INVX1 U104 ( .A(n95), .Y(\immediate<10> ) );
  INVX4 U105 ( .A(n81), .Y(\immediate<2> ) );
  INVX1 U106 ( .A(n37), .Y(n85) );
  INVX4 U107 ( .A(n85), .Y(\immediate<4> ) );
  INVX1 U108 ( .A(n4), .Y(\immediate<1> ) );
  INVX1 U109 ( .A(n120), .Y(n87) );
  INVX1 U110 ( .A(\instr<5> ), .Y(n120) );
  INVX1 U111 ( .A(n31), .Y(n88) );
  INVX1 U112 ( .A(n88), .Y(\immediate<0> ) );
  AND2X2 U113 ( .A(n37), .B(toExt), .Y(n90) );
  INVX1 U114 ( .A(\instr<1> ), .Y(n93) );
  INVX1 U115 ( .A(\writeBackData<13> ), .Y(n115) );
  INVX1 U116 ( .A(\writeBackData<15> ), .Y(n119) );
  INVX1 U117 ( .A(\writeBackData<14> ), .Y(n117) );
  INVX1 U118 ( .A(\writeBackData<12> ), .Y(n113) );
  INVX1 U119 ( .A(\writeBackData<11> ), .Y(n111) );
  INVX1 U120 ( .A(\writeBackData<10> ), .Y(n109) );
  INVX1 U121 ( .A(\writeBackData<9> ), .Y(n107) );
  INVX1 U122 ( .A(\whichImm<0> ), .Y(n91) );
  INVX1 U123 ( .A(n57), .Y(n92) );
  INVX1 U124 ( .A(\writeBackData<8> ), .Y(n105) );
  AND2X2 U125 ( .A(n36), .B(n42), .Y(n95) );
  INVX1 U126 ( .A(n95), .Y(\immediate<14> ) );
  INVX1 U127 ( .A(n95), .Y(\immediate<12> ) );
  INVX2 U128 ( .A(\regDst<0> ), .Y(n103) );
  OR2X2 U129 ( .A(n30), .B(n103), .Y(n28) );
  MUX2X1 U130 ( .B(n105), .A(n104), .S(n3), .Y(n136) );
  MUX2X1 U131 ( .B(n107), .A(n106), .S(n1), .Y(n135) );
  MUX2X1 U132 ( .B(n109), .A(n108), .S(n3), .Y(n134) );
  MUX2X1 U133 ( .B(n111), .A(n110), .S(n2), .Y(n133) );
  MUX2X1 U134 ( .B(n113), .A(n112), .S(n3), .Y(n132) );
  MUX2X1 U135 ( .B(n115), .A(n114), .S(n3), .Y(n131) );
  MUX2X1 U136 ( .B(n117), .A(n116), .S(n3), .Y(n130) );
  MUX2X1 U137 ( .B(n119), .A(n118), .S(n3), .Y(n129) );
  OAI21X1 U138 ( .A(n50), .B(n121), .C(n45), .Y(\immediate<6> ) );
  OAI21X1 U139 ( .A(n50), .B(n122), .C(n45), .Y(\immediate<7> ) );
  OR2X2 U140 ( .A(n80), .B(\whichImm<1> ), .Y(n124) );
  AOI22X1 U141 ( .A(n90), .B(n92), .C(n49), .D(\whichImm<1> ), .Y(n125) );
  OAI21X1 U142 ( .A(n79), .B(n123), .C(n42), .Y(\immediate<8> ) );
  INVX2 U143 ( .A(n30), .Y(n126) );
endmodule


module execute ( .readdata1({\readdata1<15> , \readdata1<14> , \readdata1<13> , 
        \readdata1<12> , \readdata1<11> , \readdata1<10> , \readdata1<9> , 
        \readdata1<8> , \readdata1<7> , \readdata1<6> , \readdata1<5> , 
        \readdata1<4> , \readdata1<3> , \readdata1<2> , \readdata1<1> , 
        \readdata1<0> }), .readdata2({\readdata2<15> , \readdata2<14> , 
        \readdata2<13> , \readdata2<12> , \readdata2<11> , \readdata2<10> , 
        \readdata2<9> , \readdata2<8> , \readdata2<7> , \readdata2<6> , 
        \readdata2<5> , \readdata2<4> , \readdata2<3> , \readdata2<2> , 
        \readdata2<1> , \readdata2<0> }), .immediate({\immediate<15> , 
        \immediate<14> , \immediate<13> , \immediate<12> , \immediate<11> , 
        \immediate<10> , \immediate<9> , \immediate<8> , \immediate<7> , 
        \immediate<6> , \immediate<5> , \immediate<4> , \immediate<3> , 
        \immediate<2> , \immediate<1> , \immediate<0> }), .BranchOP({
        \BranchOP<1> , \BranchOP<0> }), .ALUOp({\ALUOp<3> , \ALUOp<2> , 
        \ALUOp<1> , \ALUOp<0> }), ALUSrc, invSrc1, invSrc2, sub, .PC({\PC<15> , 
        \PC<14> , \PC<13> , \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , 
        \PC<7> , \PC<6> , \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> 
        }), jump, jumpReg, branch, .nextPC({\nextPC<15> , \nextPC<14> , 
        \nextPC<13> , \nextPC<12> , \nextPC<11> , \nextPC<10> , \nextPC<9> , 
        \nextPC<8> , \nextPC<7> , \nextPC<6> , \nextPC<5> , \nextPC<4> , 
        \nextPC<3> , \nextPC<2> , \nextPC<1> , \nextPC<0> }), .ALURes({
        \ALURes<15> , \ALURes<14> , \ALURes<13> , \ALURes<12> , \ALURes<11> , 
        \ALURes<10> , \ALURes<9> , \ALURes<8> , \ALURes<7> , \ALURes<6> , 
        \ALURes<5> , \ALURes<4> , \ALURes<3> , \ALURes<2> , \ALURes<1> , 
        \ALURes<0> }), passthrough, reverse, err );
  input \readdata1<15> , \readdata1<14> , \readdata1<13> , \readdata1<12> ,
         \readdata1<11> , \readdata1<10> , \readdata1<9> , \readdata1<8> ,
         \readdata1<7> , \readdata1<6> , \readdata1<5> , \readdata1<4> ,
         \readdata1<3> , \readdata1<2> , \readdata1<1> , \readdata1<0> ,
         \readdata2<15> , \readdata2<14> , \readdata2<13> , \readdata2<12> ,
         \readdata2<11> , \readdata2<10> , \readdata2<9> , \readdata2<8> ,
         \readdata2<7> , \readdata2<6> , \readdata2<5> , \readdata2<4> ,
         \readdata2<3> , \readdata2<2> , \readdata2<1> , \readdata2<0> ,
         \immediate<15> , \immediate<14> , \immediate<13> , \immediate<12> ,
         \immediate<11> , \immediate<10> , \immediate<9> , \immediate<8> ,
         \immediate<7> , \immediate<6> , \immediate<5> , \immediate<4> ,
         \immediate<3> , \immediate<2> , \immediate<1> , \immediate<0> ,
         \BranchOP<1> , \BranchOP<0> , \ALUOp<3> , \ALUOp<2> , \ALUOp<1> ,
         \ALUOp<0> , ALUSrc, invSrc1, invSrc2, sub, \PC<15> , \PC<14> ,
         \PC<13> , \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> ,
         \PC<6> , \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> , jump,
         jumpReg, branch, passthrough, reverse;
  output \nextPC<15> , \nextPC<14> , \nextPC<13> , \nextPC<12> , \nextPC<11> ,
         \nextPC<10> , \nextPC<9> , \nextPC<8> , \nextPC<7> , \nextPC<6> ,
         \nextPC<5> , \nextPC<4> , \nextPC<3> , \nextPC<2> , \nextPC<1> ,
         \nextPC<0> , \ALURes<15> , \ALURes<14> , \ALURes<13> , \ALURes<12> ,
         \ALURes<11> , \ALURes<10> , \ALURes<9> , \ALURes<8> , \ALURes<7> ,
         \ALURes<6> , \ALURes<5> , \ALURes<4> , \ALURes<3> , \ALURes<2> ,
         \ALURes<1> , \ALURes<0> , err;
  wire   n225, n226, n227, n228, n229, zero, \pcImmAddSum<15> ,
         \pcImmAddSum<14> , \pcImmAddSum<13> , \pcImmAddSum<12> ,
         \pcImmAddSum<11> , \pcImmAddSum<10> , \pcImmAddSum<9> ,
         \pcImmAddSum<8> , \pcImmAddSum<7> , \pcImmAddSum<6> ,
         \pcImmAddSum<5> , \pcImmAddSum<4> , \pcImmAddSum<3> ,
         \pcImmAddSum<2> , \pcImmAddSum<1> , \pcImmAddSum<0> , n78, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n92, n93,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224;
  assign err = 1'b0;

  NOR3X1 U93 ( .A(n2), .B(n140), .C(\ALUOp<1> ), .Y(n78) );
  alu ALU ( .A({\readdata1<15> , \readdata1<14> , \readdata1<13> , 
        \readdata1<12> , \readdata1<11> , \readdata1<10> , \readdata1<9> , 
        \readdata1<8> , \readdata1<7> , \readdata1<6> , \readdata1<5> , 
        \readdata1<4> , \readdata1<3> , \readdata1<2> , \readdata1<1> , 
        \readdata1<0> }), .B({n92, n211, n156, n212, n213, n214, n215, n216, 
        n217, n218, n219, n220, n221, n222, n223, n14}), .Cin(sub), .Op({n88, 
        \ALUOp<2> , \ALUOp<1> , \ALUOp<0> }), .passthrough(passthrough), 
        .reverse(reverse), .invA(invSrc1), .invB(invSrc2), .sign(n78), .Out({
        n225, \ALURes<14> , n226, \ALURes<12> , \ALURes<11> , n227, n228, 
        \ALURes<8> , n229, \ALURes<6> , \ALURes<5> , \ALURes<4> , \ALURes<3> , 
        \ALURes<2> , \ALURes<1> , \ALURes<0> }), .Ofl(), .zero(zero) );
  adder_1 pcImmAdd ( .A({\PC<15> , \PC<14> , \PC<13> , \PC<12> , \PC<11> , 
        \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> , \PC<4> , 
        \PC<3> , \PC<2> , \PC<1> , \PC<0> }), .B({n155, n148, n102, n161, n100, 
        n149, n160, n158, n145, n151, n157, \immediate<4> , \immediate<3> , 
        \immediate<2> , \immediate<1> , \immediate<0> }), .Cin(1'b0), 
        .Overflow(), .Cout(), .Sum({\pcImmAddSum<15> , \pcImmAddSum<14> , 
        \pcImmAddSum<13> , \pcImmAddSum<12> , \pcImmAddSum<11> , 
        \pcImmAddSum<10> , \pcImmAddSum<9> , \pcImmAddSum<8> , 
        \pcImmAddSum<7> , \pcImmAddSum<6> , \pcImmAddSum<5> , \pcImmAddSum<4> , 
        \pcImmAddSum<3> , \pcImmAddSum<2> , \pcImmAddSum<1> , \pcImmAddSum<0> }) );
  BUFX2 U3 ( .A(\ALUOp<2> ), .Y(n2) );
  BUFX2 U4 ( .A(\ALUOp<0> ), .Y(n3) );
  INVX4 U5 ( .A(n163), .Y(n218) );
  BUFX4 U6 ( .A(n229), .Y(\ALURes<7> ) );
  INVX1 U7 ( .A(\readdata2<9> ), .Y(n180) );
  INVX1 U8 ( .A(\readdata2<4> ), .Y(n176) );
  INVX1 U9 ( .A(\readdata2<1> ), .Y(n170) );
  INVX1 U10 ( .A(\readdata2<2> ), .Y(n172) );
  INVX1 U11 ( .A(\readdata2<5> ), .Y(n178) );
  INVX1 U12 ( .A(\readdata2<12> ), .Y(n182) );
  INVX1 U13 ( .A(\BranchOP<0> ), .Y(n99) );
  INVX1 U14 ( .A(\readdata2<14> ), .Y(n185) );
  INVX1 U15 ( .A(n162), .Y(n217) );
  INVX1 U16 ( .A(\readdata2<3> ), .Y(n174) );
  AND2X1 U17 ( .A(n97), .B(n224), .Y(n139) );
  INVX2 U18 ( .A(n12), .Y(n4) );
  INVX2 U19 ( .A(n12), .Y(n5) );
  INVX2 U20 ( .A(n12), .Y(n13) );
  AND2X2 U21 ( .A(n194), .B(n10), .Y(n6) );
  AND2X2 U22 ( .A(n194), .B(n10), .Y(n7) );
  BUFX2 U23 ( .A(\ALURes<3> ), .Y(n8) );
  BUFX4 U24 ( .A(n225), .Y(\ALURes<15> ) );
  INVX1 U25 ( .A(n193), .Y(n9) );
  INVX1 U26 ( .A(n9), .Y(n10) );
  OR2X2 U27 ( .A(n193), .B(jumpReg), .Y(n12) );
  MUX2X1 U28 ( .B(n169), .A(n170), .S(n153), .Y(n223) );
  BUFX2 U29 ( .A(n228), .Y(\ALURes<9> ) );
  BUFX4 U30 ( .A(n96), .Y(n152) );
  BUFX4 U31 ( .A(n152), .Y(n11) );
  AND2X2 U32 ( .A(n22), .B(n20), .Y(n14) );
  AND2X2 U33 ( .A(n101), .B(n11), .Y(n15) );
  INVX1 U34 ( .A(n15), .Y(n16) );
  AND2X2 U35 ( .A(n186), .B(n11), .Y(n17) );
  INVX1 U36 ( .A(n17), .Y(n18) );
  AND2X2 U37 ( .A(n167), .B(n152), .Y(n19) );
  INVX1 U38 ( .A(n19), .Y(n20) );
  AND2X2 U39 ( .A(n168), .B(n153), .Y(n21) );
  INVX1 U40 ( .A(n21), .Y(n22) );
  AND2X2 U41 ( .A(\pcImmAddSum<0> ), .B(n93), .Y(n23) );
  INVX1 U42 ( .A(n23), .Y(n24) );
  AND2X2 U43 ( .A(\pcImmAddSum<1> ), .B(n7), .Y(n25) );
  INVX1 U44 ( .A(n25), .Y(n26) );
  AND2X2 U45 ( .A(\pcImmAddSum<2> ), .B(n93), .Y(n27) );
  INVX1 U46 ( .A(n27), .Y(n28) );
  AND2X2 U47 ( .A(\pcImmAddSum<3> ), .B(n7), .Y(n29) );
  INVX1 U48 ( .A(n29), .Y(n30) );
  AND2X2 U49 ( .A(\pcImmAddSum<4> ), .B(n7), .Y(n31) );
  INVX1 U50 ( .A(n31), .Y(n32) );
  AND2X2 U51 ( .A(\pcImmAddSum<5> ), .B(n6), .Y(n33) );
  INVX1 U52 ( .A(n33), .Y(n34) );
  AND2X2 U53 ( .A(\pcImmAddSum<6> ), .B(n7), .Y(n35) );
  INVX1 U54 ( .A(n35), .Y(n36) );
  AND2X2 U55 ( .A(\pcImmAddSum<7> ), .B(n6), .Y(n37) );
  INVX1 U56 ( .A(n37), .Y(n38) );
  AND2X2 U57 ( .A(\pcImmAddSum<8> ), .B(n6), .Y(n39) );
  INVX1 U58 ( .A(n39), .Y(n40) );
  AND2X2 U59 ( .A(\pcImmAddSum<9> ), .B(n93), .Y(n41) );
  INVX1 U60 ( .A(n41), .Y(n42) );
  AND2X2 U61 ( .A(\pcImmAddSum<10> ), .B(n6), .Y(n43) );
  INVX1 U62 ( .A(n43), .Y(n44) );
  AND2X2 U63 ( .A(\pcImmAddSum<11> ), .B(n93), .Y(n45) );
  INVX1 U64 ( .A(n45), .Y(n46) );
  AND2X2 U65 ( .A(\pcImmAddSum<12> ), .B(n93), .Y(n47) );
  INVX1 U66 ( .A(n47), .Y(n48) );
  AND2X2 U67 ( .A(\pcImmAddSum<13> ), .B(n7), .Y(n49) );
  INVX1 U68 ( .A(n49), .Y(n50) );
  AND2X2 U69 ( .A(\pcImmAddSum<14> ), .B(n93), .Y(n51) );
  INVX1 U70 ( .A(n51), .Y(n52) );
  AND2X2 U71 ( .A(\pcImmAddSum<15> ), .B(n6), .Y(n53) );
  INVX1 U72 ( .A(n53), .Y(n54) );
  AND2X2 U73 ( .A(\PC<0> ), .B(n4), .Y(n55) );
  INVX1 U74 ( .A(n55), .Y(n56) );
  AND2X2 U75 ( .A(\PC<1> ), .B(n5), .Y(n57) );
  INVX1 U76 ( .A(n57), .Y(n58) );
  AND2X2 U77 ( .A(\PC<2> ), .B(n13), .Y(n59) );
  INVX1 U78 ( .A(n59), .Y(n60) );
  AND2X2 U79 ( .A(\PC<3> ), .B(n5), .Y(n61) );
  INVX1 U80 ( .A(n61), .Y(n62) );
  AND2X2 U81 ( .A(\PC<4> ), .B(n4), .Y(n63) );
  INVX1 U82 ( .A(n63), .Y(n64) );
  AND2X2 U83 ( .A(\PC<5> ), .B(n4), .Y(n65) );
  INVX1 U84 ( .A(n65), .Y(n66) );
  AND2X2 U85 ( .A(\PC<6> ), .B(n13), .Y(n67) );
  INVX1 U86 ( .A(n67), .Y(n68) );
  AND2X2 U87 ( .A(\PC<7> ), .B(n13), .Y(n69) );
  INVX1 U88 ( .A(n69), .Y(n70) );
  AND2X2 U89 ( .A(\PC<8> ), .B(n5), .Y(n71) );
  INVX1 U90 ( .A(n71), .Y(n72) );
  AND2X2 U91 ( .A(\PC<9> ), .B(n4), .Y(n73) );
  INVX1 U92 ( .A(n73), .Y(n74) );
  AND2X2 U94 ( .A(\PC<10> ), .B(n5), .Y(n75) );
  INVX1 U95 ( .A(n75), .Y(n76) );
  AND2X2 U96 ( .A(\PC<11> ), .B(n4), .Y(n77) );
  INVX1 U97 ( .A(n77), .Y(n79) );
  AND2X2 U98 ( .A(\PC<12> ), .B(n5), .Y(n80) );
  INVX1 U99 ( .A(n80), .Y(n81) );
  AND2X2 U100 ( .A(\PC<13> ), .B(n5), .Y(n82) );
  INVX1 U101 ( .A(n82), .Y(n83) );
  AND2X2 U102 ( .A(\PC<14> ), .B(n4), .Y(n84) );
  INVX1 U103 ( .A(n84), .Y(n85) );
  AND2X2 U104 ( .A(\PC<15> ), .B(n13), .Y(n86) );
  INVX1 U105 ( .A(n86), .Y(n87) );
  BUFX2 U106 ( .A(\ALUOp<3> ), .Y(n88) );
  BUFX2 U107 ( .A(n226), .Y(\ALURes<13> ) );
  BUFX2 U108 ( .A(n227), .Y(\ALURes<10> ) );
  AND2X2 U109 ( .A(n18), .B(n106), .Y(n92) );
  AND2X2 U110 ( .A(n194), .B(n10), .Y(n93) );
  BUFX2 U111 ( .A(ALUSrc), .Y(n96) );
  BUFX2 U112 ( .A(n88), .Y(n97) );
  BUFX2 U113 ( .A(\ALURes<15> ), .Y(n98) );
  MUX2X1 U114 ( .B(\immediate<8> ), .A(\readdata2<8> ), .S(n159), .Y(n164) );
  AND2X2 U115 ( .A(\ALURes<4> ), .B(jumpReg), .Y(n115) );
  XNOR2X1 U116 ( .A(zero), .B(n99), .Y(n189) );
  BUFX2 U117 ( .A(\immediate<11> ), .Y(n100) );
  INVX2 U118 ( .A(n164), .Y(n216) );
  INVX1 U119 ( .A(\immediate<9> ), .Y(n179) );
  INVX1 U120 ( .A(\immediate<13> ), .Y(n101) );
  INVX1 U121 ( .A(n101), .Y(n102) );
  INVX1 U122 ( .A(jumpReg), .Y(n194) );
  AND2X1 U123 ( .A(n143), .B(jumpReg), .Y(n117) );
  AND2X2 U124 ( .A(n183), .B(n159), .Y(n103) );
  INVX1 U125 ( .A(n103), .Y(n104) );
  AND2X2 U126 ( .A(n187), .B(n159), .Y(n105) );
  INVX1 U127 ( .A(n105), .Y(n106) );
  AND2X2 U128 ( .A(jumpReg), .B(n154), .Y(n107) );
  INVX1 U129 ( .A(n107), .Y(n108) );
  AND2X2 U130 ( .A(jumpReg), .B(\ALURes<1> ), .Y(n109) );
  INVX1 U131 ( .A(n109), .Y(n110) );
  AND2X2 U132 ( .A(jumpReg), .B(n144), .Y(n111) );
  INVX1 U133 ( .A(n111), .Y(n112) );
  AND2X2 U134 ( .A(n8), .B(jumpReg), .Y(n113) );
  INVX1 U135 ( .A(n113), .Y(n114) );
  INVX1 U136 ( .A(n115), .Y(n116) );
  INVX1 U137 ( .A(n117), .Y(n118) );
  AND2X2 U138 ( .A(\ALURes<6> ), .B(jumpReg), .Y(n119) );
  INVX1 U139 ( .A(n119), .Y(n120) );
  AND2X2 U140 ( .A(jumpReg), .B(\ALURes<7> ), .Y(n121) );
  INVX1 U141 ( .A(n121), .Y(n122) );
  AND2X2 U142 ( .A(\ALURes<8> ), .B(jumpReg), .Y(n123) );
  INVX1 U143 ( .A(n123), .Y(n124) );
  AND2X2 U144 ( .A(jumpReg), .B(n142), .Y(n125) );
  INVX1 U145 ( .A(n125), .Y(n126) );
  AND2X2 U146 ( .A(\ALURes<10> ), .B(jumpReg), .Y(n127) );
  INVX1 U147 ( .A(n127), .Y(n128) );
  AND2X2 U148 ( .A(jumpReg), .B(\ALURes<11> ), .Y(n129) );
  INVX1 U149 ( .A(n129), .Y(n130) );
  AND2X2 U150 ( .A(\ALURes<12> ), .B(jumpReg), .Y(n131) );
  INVX1 U151 ( .A(n131), .Y(n132) );
  AND2X2 U152 ( .A(jumpReg), .B(n146), .Y(n133) );
  INVX1 U153 ( .A(n133), .Y(n134) );
  AND2X2 U154 ( .A(\ALURes<14> ), .B(jumpReg), .Y(n135) );
  INVX1 U155 ( .A(n135), .Y(n136) );
  AND2X2 U156 ( .A(jumpReg), .B(n98), .Y(n137) );
  INVX1 U157 ( .A(n137), .Y(n138) );
  INVX1 U158 ( .A(n139), .Y(n140) );
  OAI21X1 U159 ( .A(n191), .B(n192), .C(n190), .Y(n193) );
  INVX1 U160 ( .A(jump), .Y(n190) );
  INVX1 U161 ( .A(\ALURes<9> ), .Y(n141) );
  INVX1 U162 ( .A(n141), .Y(n142) );
  BUFX2 U163 ( .A(\ALURes<5> ), .Y(n143) );
  BUFX2 U164 ( .A(\ALURes<2> ), .Y(n144) );
  BUFX2 U165 ( .A(\immediate<7> ), .Y(n145) );
  BUFX2 U166 ( .A(\ALURes<13> ), .Y(n146) );
  INVX1 U167 ( .A(\immediate<3> ), .Y(n173) );
  INVX1 U168 ( .A(\immediate<2> ), .Y(n171) );
  INVX2 U169 ( .A(n166), .Y(n213) );
  INVX1 U170 ( .A(n96), .Y(n153) );
  INVX1 U171 ( .A(\immediate<14> ), .Y(n147) );
  INVX1 U172 ( .A(n147), .Y(n148) );
  BUFX2 U173 ( .A(\immediate<10> ), .Y(n149) );
  INVX1 U174 ( .A(\immediate<6> ), .Y(n150) );
  INVX1 U175 ( .A(n150), .Y(n151) );
  BUFX2 U176 ( .A(\immediate<8> ), .Y(n158) );
  INVX1 U177 ( .A(\readdata2<0> ), .Y(n168) );
  INVX1 U178 ( .A(branch), .Y(n191) );
  BUFX2 U179 ( .A(\ALURes<0> ), .Y(n154) );
  INVX4 U180 ( .A(n186), .Y(n155) );
  AND2X2 U181 ( .A(n16), .B(n104), .Y(n156) );
  INVX1 U182 ( .A(n177), .Y(n157) );
  INVX1 U183 ( .A(\immediate<5> ), .Y(n177) );
  INVX1 U184 ( .A(n11), .Y(n159) );
  INVX1 U185 ( .A(\readdata2<13> ), .Y(n183) );
  INVX1 U186 ( .A(n179), .Y(n160) );
  INVX2 U187 ( .A(n165), .Y(n214) );
  INVX1 U188 ( .A(\immediate<4> ), .Y(n175) );
  INVX1 U189 ( .A(n181), .Y(n161) );
  INVX1 U190 ( .A(\immediate<12> ), .Y(n181) );
  INVX1 U191 ( .A(\readdata2<15> ), .Y(n187) );
  INVX1 U192 ( .A(\immediate<15> ), .Y(n186) );
  MUX2X1 U193 ( .B(\readdata2<7> ), .A(\immediate<7> ), .S(n11), .Y(n162) );
  MUX2X1 U194 ( .B(\readdata2<6> ), .A(\immediate<6> ), .S(n11), .Y(n163) );
  INVX1 U195 ( .A(\immediate<14> ), .Y(n184) );
  INVX1 U196 ( .A(\immediate<1> ), .Y(n169) );
  MUX2X1 U197 ( .B(\readdata2<10> ), .A(\immediate<10> ), .S(n11), .Y(n165) );
  INVX1 U198 ( .A(\immediate<0> ), .Y(n167) );
  MUX2X1 U199 ( .B(\readdata2<11> ), .A(\immediate<11> ), .S(n11), .Y(n166) );
  INVX1 U200 ( .A(n3), .Y(n224) );
  MUX2X1 U201 ( .B(n172), .A(n171), .S(n152), .Y(n222) );
  MUX2X1 U202 ( .B(n174), .A(n173), .S(n11), .Y(n221) );
  MUX2X1 U203 ( .B(n176), .A(n175), .S(n11), .Y(n220) );
  MUX2X1 U204 ( .B(n178), .A(n177), .S(n11), .Y(n219) );
  MUX2X1 U205 ( .B(n180), .A(n179), .S(n11), .Y(n215) );
  MUX2X1 U206 ( .B(n182), .A(n181), .S(n11), .Y(n212) );
  MUX2X1 U207 ( .B(n185), .A(n184), .S(n11), .Y(n211) );
  XOR2X1 U208 ( .A(\BranchOP<0> ), .B(\readdata1<15> ), .Y(n188) );
  MUX2X1 U209 ( .B(n189), .A(n188), .S(\BranchOP<1> ), .Y(n192) );
  NAND3X1 U210 ( .A(n24), .B(n108), .C(n56), .Y(\nextPC<0> ) );
  NAND3X1 U211 ( .A(n26), .B(n110), .C(n58), .Y(\nextPC<1> ) );
  NAND3X1 U212 ( .A(n28), .B(n112), .C(n60), .Y(\nextPC<2> ) );
  NAND3X1 U213 ( .A(n30), .B(n114), .C(n62), .Y(\nextPC<3> ) );
  NAND3X1 U214 ( .A(n32), .B(n116), .C(n64), .Y(\nextPC<4> ) );
  NAND3X1 U215 ( .A(n34), .B(n118), .C(n66), .Y(\nextPC<5> ) );
  NAND3X1 U216 ( .A(n36), .B(n120), .C(n68), .Y(\nextPC<6> ) );
  NAND3X1 U217 ( .A(n38), .B(n122), .C(n70), .Y(\nextPC<7> ) );
  NAND3X1 U218 ( .A(n40), .B(n124), .C(n72), .Y(\nextPC<8> ) );
  NAND3X1 U219 ( .A(n42), .B(n126), .C(n74), .Y(\nextPC<9> ) );
  NAND3X1 U220 ( .A(n44), .B(n128), .C(n76), .Y(\nextPC<10> ) );
  NAND3X1 U221 ( .A(n46), .B(n130), .C(n79), .Y(\nextPC<11> ) );
  NAND3X1 U222 ( .A(n48), .B(n132), .C(n81), .Y(\nextPC<12> ) );
  NAND3X1 U223 ( .A(n50), .B(n134), .C(n83), .Y(\nextPC<13> ) );
  NAND3X1 U224 ( .A(n52), .B(n136), .C(n85), .Y(\nextPC<14> ) );
  NAND3X1 U225 ( .A(n54), .B(n138), .C(n87), .Y(\nextPC<15> ) );
endmodule


module memory ( clk, rst, .addr({\addr<15> , \addr<14> , \addr<13> , 
        \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , 
        \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , 
        \addr<0> }), .writeData({\writeData<15> , \writeData<14> , 
        \writeData<13> , \writeData<12> , \writeData<11> , \writeData<10> , 
        \writeData<9> , \writeData<8> , \writeData<7> , \writeData<6> , 
        \writeData<5> , \writeData<4> , \writeData<3> , \writeData<2> , 
        \writeData<1> , \writeData<0> }), halt, memWrite, memRead, .readData({
        \readData<15> , \readData<14> , \readData<13> , \readData<12> , 
        \readData<11> , \readData<10> , \readData<9> , \readData<8> , 
        \readData<7> , \readData<6> , \readData<5> , \readData<4> , 
        \readData<3> , \readData<2> , \readData<1> , \readData<0> }), err );
  input clk, rst, \addr<15> , \addr<14> , \addr<13> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> ,
         \writeData<15> , \writeData<14> , \writeData<13> , \writeData<12> ,
         \writeData<11> , \writeData<10> , \writeData<9> , \writeData<8> ,
         \writeData<7> , \writeData<6> , \writeData<5> , \writeData<4> ,
         \writeData<3> , \writeData<2> , \writeData<1> , \writeData<0> , halt,
         memWrite, memRead;
  output \readData<15> , \readData<14> , \readData<13> , \readData<12> ,
         \readData<11> , \readData<10> , \readData<9> , \readData<8> ,
         \readData<7> , \readData<6> , \readData<5> , \readData<4> ,
         \readData<3> , \readData<2> , \readData<1> , \readData<0> , err;
  wire   n1;
  assign err = 1'b0;

  memory2c_0 instrmem ( .data_out({\readData<15> , \readData<14> , 
        \readData<13> , \readData<12> , \readData<11> , \readData<10> , 
        \readData<9> , \readData<8> , \readData<7> , \readData<6> , 
        \readData<5> , \readData<4> , \readData<3> , \readData<2> , 
        \readData<1> , \readData<0> }), .data_in({\writeData<15> , 
        \writeData<14> , \writeData<13> , \writeData<12> , \writeData<11> , 
        \writeData<10> , \writeData<9> , \writeData<8> , \writeData<7> , 
        \writeData<6> , \writeData<5> , \writeData<4> , \writeData<3> , 
        \writeData<2> , \writeData<1> , \writeData<0> }), .addr({\addr<15> , 
        \addr<14> , \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), .enable(n1), .wr(memWrite), 
        .createdump(halt), .clk(clk), .rst(rst) );
  INVX2 U2 ( .A(halt), .Y(n1) );
endmodule


module writeBack ( .memData({\memData<15> , \memData<14> , \memData<13> , 
        \memData<12> , \memData<11> , \memData<10> , \memData<9> , 
        \memData<8> , \memData<7> , \memData<6> , \memData<5> , \memData<4> , 
        \memData<3> , \memData<2> , \memData<1> , \memData<0> }), .ALUData({
        \ALUData<15> , \ALUData<14> , \ALUData<13> , \ALUData<12> , 
        \ALUData<11> , \ALUData<10> , \ALUData<9> , \ALUData<8> , \ALUData<7> , 
        \ALUData<6> , \ALUData<5> , \ALUData<4> , \ALUData<3> , \ALUData<2> , 
        \ALUData<1> , \ALUData<0> }), memToReg, .writeBackData({
        \writeBackData<15> , \writeBackData<14> , \writeBackData<13> , 
        \writeBackData<12> , \writeBackData<11> , \writeBackData<10> , 
        \writeBackData<9> , \writeBackData<8> , \writeBackData<7> , 
        \writeBackData<6> , \writeBackData<5> , \writeBackData<4> , 
        \writeBackData<3> , \writeBackData<2> , \writeBackData<1> , 
        \writeBackData<0> }), err );
  input \memData<15> , \memData<14> , \memData<13> , \memData<12> ,
         \memData<11> , \memData<10> , \memData<9> , \memData<8> ,
         \memData<7> , \memData<6> , \memData<5> , \memData<4> , \memData<3> ,
         \memData<2> , \memData<1> , \memData<0> , \ALUData<15> ,
         \ALUData<14> , \ALUData<13> , \ALUData<12> , \ALUData<11> ,
         \ALUData<10> , \ALUData<9> , \ALUData<8> , \ALUData<7> , \ALUData<6> ,
         \ALUData<5> , \ALUData<4> , \ALUData<3> , \ALUData<2> , \ALUData<1> ,
         \ALUData<0> , memToReg;
  output \writeBackData<15> , \writeBackData<14> , \writeBackData<13> ,
         \writeBackData<12> , \writeBackData<11> , \writeBackData<10> ,
         \writeBackData<9> , \writeBackData<8> , \writeBackData<7> ,
         \writeBackData<6> , \writeBackData<5> , \writeBackData<4> ,
         \writeBackData<3> , \writeBackData<2> , \writeBackData<1> ,
         \writeBackData<0> , err;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52;
  assign err = 1'b0;

  INVX1 U2 ( .A(n25), .Y(n20) );
  INVX1 U3 ( .A(n25), .Y(n1) );
  INVX1 U4 ( .A(n25), .Y(n22) );
  INVX1 U5 ( .A(n25), .Y(n23) );
  INVX1 U6 ( .A(n25), .Y(n19) );
  INVX2 U7 ( .A(n25), .Y(n21) );
  INVX1 U8 ( .A(n25), .Y(n18) );
  INVX2 U9 ( .A(memToReg), .Y(n24) );
  INVX1 U10 ( .A(n25), .Y(n29) );
  INVX1 U11 ( .A(n25), .Y(n27) );
  MUX2X1 U12 ( .B(n41), .A(n42), .S(n1), .Y(\writeBackData<10> ) );
  AND2X2 U13 ( .A(\ALUData<0> ), .B(n35), .Y(n2) );
  INVX1 U14 ( .A(n2), .Y(n3) );
  AND2X2 U15 ( .A(\ALUData<1> ), .B(n35), .Y(n4) );
  INVX1 U16 ( .A(n4), .Y(n5) );
  AND2X2 U17 ( .A(\ALUData<2> ), .B(n35), .Y(n6) );
  INVX1 U18 ( .A(n6), .Y(n7) );
  AND2X2 U19 ( .A(\ALUData<3> ), .B(n35), .Y(n8) );
  INVX1 U20 ( .A(n8), .Y(n9) );
  AND2X2 U21 ( .A(\ALUData<4> ), .B(n35), .Y(n10) );
  INVX1 U22 ( .A(n10), .Y(n11) );
  AND2X2 U23 ( .A(\ALUData<5> ), .B(n35), .Y(n12) );
  INVX1 U24 ( .A(n12), .Y(n13) );
  AND2X2 U25 ( .A(\ALUData<6> ), .B(n35), .Y(n14) );
  INVX1 U26 ( .A(n14), .Y(n15) );
  AND2X2 U27 ( .A(\ALUData<7> ), .B(n35), .Y(n16) );
  INVX1 U28 ( .A(n16), .Y(n17) );
  MUX2X1 U29 ( .B(n45), .A(n46), .S(n18), .Y(\writeBackData<12> ) );
  INVX1 U30 ( .A(\ALUData<12> ), .Y(n46) );
  MUX2X1 U31 ( .B(n39), .A(n40), .S(n19), .Y(\writeBackData<9> ) );
  MUX2X1 U32 ( .B(n37), .A(n38), .S(n20), .Y(\writeBackData<8> ) );
  MUX2X1 U33 ( .B(n43), .A(n44), .S(n21), .Y(\writeBackData<11> ) );
  MUX2X1 U34 ( .B(n47), .A(n48), .S(n22), .Y(\writeBackData<13> ) );
  MUX2X1 U35 ( .B(n51), .A(n52), .S(n27), .Y(\writeBackData<15> ) );
  MUX2X1 U36 ( .B(n49), .A(n50), .S(n23), .Y(\writeBackData<14> ) );
  INVX1 U37 ( .A(\memData<15> ), .Y(n51) );
  INVX1 U38 ( .A(\memData<10> ), .Y(n41) );
  INVX1 U39 ( .A(\ALUData<15> ), .Y(n52) );
  INVX1 U40 ( .A(\memData<14> ), .Y(n49) );
  INVX1 U41 ( .A(\memData<13> ), .Y(n47) );
  INVX1 U42 ( .A(\memData<12> ), .Y(n45) );
  INVX1 U43 ( .A(\memData<11> ), .Y(n43) );
  INVX1 U44 ( .A(\ALUData<9> ), .Y(n40) );
  INVX1 U45 ( .A(\memData<9> ), .Y(n39) );
  INVX1 U46 ( .A(\memData<8> ), .Y(n37) );
  INVX1 U47 ( .A(\ALUData<10> ), .Y(n42) );
  INVX1 U48 ( .A(\memData<3> ), .Y(n31) );
  INVX1 U49 ( .A(\memData<2> ), .Y(n30) );
  INVX1 U50 ( .A(\memData<1> ), .Y(n28) );
  INVX1 U51 ( .A(\memData<0> ), .Y(n26) );
  INVX1 U52 ( .A(\memData<7> ), .Y(n36) );
  INVX1 U53 ( .A(\memData<5> ), .Y(n33) );
  INVX1 U54 ( .A(\memData<6> ), .Y(n34) );
  INVX1 U55 ( .A(\ALUData<14> ), .Y(n50) );
  INVX1 U56 ( .A(\memData<4> ), .Y(n32) );
  INVX1 U57 ( .A(\ALUData<13> ), .Y(n48) );
  INVX1 U58 ( .A(\ALUData<8> ), .Y(n38) );
  INVX1 U59 ( .A(\ALUData<11> ), .Y(n44) );
  INVX8 U60 ( .A(n24), .Y(n25) );
  INVX2 U61 ( .A(memToReg), .Y(n35) );
  AOI22X1 U62 ( .A(n3), .B(n27), .C(n3), .D(n26), .Y(\writeBackData<0> ) );
  AOI22X1 U63 ( .A(n5), .B(n29), .C(n5), .D(n28), .Y(\writeBackData<1> ) );
  AOI22X1 U64 ( .A(n7), .B(n29), .C(n7), .D(n30), .Y(\writeBackData<2> ) );
  AOI22X1 U65 ( .A(n9), .B(n29), .C(n9), .D(n31), .Y(\writeBackData<3> ) );
  AOI22X1 U66 ( .A(n11), .B(n18), .C(n11), .D(n32), .Y(\writeBackData<4> ) );
  AOI22X1 U67 ( .A(n13), .B(n29), .C(n13), .D(n33), .Y(\writeBackData<5> ) );
  AOI22X1 U68 ( .A(n15), .B(n29), .C(n15), .D(n34), .Y(\writeBackData<6> ) );
  AOI22X1 U69 ( .A(n17), .B(n29), .C(n17), .D(n36), .Y(\writeBackData<7> ) );
endmodule


module proc ( err, clk, rst );
  input clk, rst;
  output err;
  wire   decodeErr, halt, \nextPC<15> , \nextPC<14> , \nextPC<13> ,
         \nextPC<12> , \nextPC<11> , \nextPC<10> , \nextPC<9> , \nextPC<8> ,
         \nextPC<7> , \nextPC<6> , \nextPC<5> , \nextPC<4> , \nextPC<3> ,
         \nextPC<2> , \nextPC<1> , \nextPC<0> , \PC<15> , \PC<14> , \PC<13> ,
         \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> ,
         \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> , \instr<15> ,
         \instr<14> , \instr<13> , \instr<12> , \instr<11> , \instr<10> ,
         \instr<9> , \instr<8> , \instr<7> , \instr<6> , \instr<5> ,
         \instr<4> , \instr<3> , \instr<2> , \instr<1> , \instr<0> ,
         \writeBackData<15> , \writeBackData<14> , \writeBackData<13> ,
         \writeBackData<12> , \writeBackData<11> , \writeBackData<10> ,
         \writeBackData<9> , \writeBackData<8> , \writeBackData<7> ,
         \writeBackData<6> , \writeBackData<5> , \writeBackData<4> ,
         \writeBackData<3> , \writeBackData<2> , \writeBackData<1> ,
         \writeBackData<0> , \readdata1<15> , \readdata1<14> , \readdata1<13> ,
         \readdata1<12> , \readdata1<11> , \readdata1<10> , \readdata1<9> ,
         \readdata1<8> , \readdata1<7> , \readdata1<6> , \readdata1<5> ,
         \readdata1<4> , \readdata1<3> , \readdata1<2> , \readdata1<1> ,
         \readdata1<0> , \readdata2<15> , \readdata2<14> , \readdata2<13> ,
         \readdata2<12> , \readdata2<11> , \readdata2<10> , \readdata2<9> ,
         \readdata2<8> , \readdata2<7> , \readdata2<6> , \readdata2<5> ,
         \readdata2<4> , \readdata2<3> , \readdata2<2> , \readdata2<1> ,
         \readdata2<0> , \immediate<15> , \immediate<14> , \immediate<13> ,
         \immediate<12> , \immediate<11> , \immediate<10> , \immediate<9> ,
         \immediate<8> , \immediate<7> , \immediate<6> , \immediate<5> ,
         \immediate<4> , \immediate<3> , \immediate<2> , \immediate<1> ,
         \immediate<0> , jump, jumpReg, branch, \branchOp<1> , \branchOp<0> ,
         memRead, memWrite, memToReg, \ALUOp<3> , \ALUOp<2> , \ALUOp<1> ,
         \ALUOp<0> , ALUSrc, invSrc1, invSrc2, sub, passthrough, reverse,
         \ALURes<15> , \ALURes<14> , \ALURes<13> , \ALURes<12> , \ALURes<11> ,
         \ALURes<10> , \ALURes<9> , \ALURes<8> , \ALURes<7> , \ALURes<6> ,
         \ALURes<5> , \ALURes<4> , \ALURes<3> , \ALURes<2> , \ALURes<1> ,
         \ALURes<0> , \readData<15> , \readData<14> , \readData<13> ,
         \readData<12> , \readData<11> , \readData<10> , \readData<9> ,
         \readData<8> , \readData<7> , \readData<6> , \readData<5> ,
         \readData<4> , \readData<3> , \readData<2> , \readData<1> ,
         \readData<0> , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n19, n20;
  assign err = 1'b0;

  fetch fetch0 ( .clk(clk), .rst(n19), .halt(halt), .nextPC({\nextPC<15> , 
        \nextPC<14> , \nextPC<13> , \nextPC<12> , \nextPC<11> , \nextPC<10> , 
        \nextPC<9> , \nextPC<8> , \nextPC<7> , \nextPC<6> , \nextPC<5> , 
        \nextPC<4> , \nextPC<3> , \nextPC<2> , \nextPC<1> , \nextPC<0> }), 
        .PC2({\PC<15> , \PC<14> , \PC<13> , \PC<12> , \PC<11> , \PC<10> , 
        \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> , \PC<4> , \PC<3> , \PC<2> , 
        \PC<1> , \PC<0> }), .instr({\instr<15> , \instr<14> , \instr<13> , 
        \instr<12> , \instr<11> , \instr<10> , \instr<9> , \instr<8> , 
        \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> , \instr<2> , 
        \instr<1> , \instr<0> }), .err() );
  decode decode0 ( .clk(clk), .rst(n19), .instr({\instr<15> , \instr<14> , 
        \instr<13> , \instr<12> , \instr<11> , \instr<10> , \instr<9> , 
        \instr<8> , \instr<7> , \instr<6> , \instr<5> , \instr<4> , \instr<3> , 
        \instr<2> , \instr<1> , \instr<0> }), .PC({\PC<15> , \PC<14> , 
        \PC<13> , \PC<12> , \PC<11> , \PC<10> , \PC<9> , \PC<8> , \PC<7> , 
        \PC<6> , \PC<5> , \PC<4> , \PC<3> , \PC<2> , \PC<1> , \PC<0> }), 
        .writeBackData({\writeBackData<15> , \writeBackData<14> , 
        \writeBackData<13> , \writeBackData<12> , \writeBackData<11> , 
        \writeBackData<10> , \writeBackData<9> , \writeBackData<8> , 
        \writeBackData<7> , \writeBackData<6> , \writeBackData<5> , 
        \writeBackData<4> , \writeBackData<3> , \writeBackData<2> , 
        \writeBackData<1> , \writeBackData<0> }), .readdata1({\readdata1<15> , 
        \readdata1<14> , \readdata1<13> , \readdata1<12> , \readdata1<11> , 
        \readdata1<10> , \readdata1<9> , \readdata1<8> , \readdata1<7> , 
        \readdata1<6> , \readdata1<5> , \readdata1<4> , \readdata1<3> , 
        \readdata1<2> , \readdata1<1> , \readdata1<0> }), .readdata2({
        \readdata2<15> , \readdata2<14> , \readdata2<13> , \readdata2<12> , 
        \readdata2<11> , \readdata2<10> , \readdata2<9> , \readdata2<8> , 
        \readdata2<7> , \readdata2<6> , \readdata2<5> , \readdata2<4> , 
        \readdata2<3> , \readdata2<2> , \readdata2<1> , \readdata2<0> }), 
        .immediate({\immediate<15> , \immediate<14> , \immediate<13> , 
        \immediate<12> , \immediate<11> , \immediate<10> , \immediate<9> , 
        \immediate<8> , \immediate<7> , \immediate<6> , \immediate<5> , 
        \immediate<4> , \immediate<3> , \immediate<2> , \immediate<1> , 
        \immediate<0> }), .jump(jump), .jumpReg(jumpReg), .branch(branch), 
        .branchOp({\branchOp<1> , \branchOp<0> }), .memRead(memRead), 
        .memWrite(memWrite), .memToReg(memToReg), .ALUOp({\ALUOp<3> , 
        \ALUOp<2> , \ALUOp<1> , \ALUOp<0> }), .ALUSrc(ALUSrc), .invSrc1(
        invSrc1), .invSrc2(invSrc2), .sub(sub), .halt(halt), .passthrough(
        passthrough), .reverse(reverse), .err(decodeErr) );
  execute ex0 ( .readdata1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .readdata2({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .immediate({\immediate<12> , \immediate<14> , 
        \immediate<13> , \immediate<12> , \immediate<11> , \immediate<10> , 
        \immediate<9> , \immediate<8> , \immediate<7> , \immediate<6> , 
        \immediate<5> , \immediate<4> , \immediate<3> , \immediate<2> , 
        \immediate<1> , \immediate<0> }), .BranchOP({\branchOp<1> , 
        \branchOp<0> }), .ALUOp({\ALUOp<3> , \ALUOp<2> , \ALUOp<1> , 
        \ALUOp<0> }), .ALUSrc(ALUSrc), .invSrc1(invSrc1), .invSrc2(invSrc2), 
        .sub(sub), .PC({\PC<15> , \PC<14> , \PC<13> , \PC<12> , \PC<11> , 
        \PC<10> , \PC<9> , \PC<8> , \PC<7> , \PC<6> , \PC<5> , \PC<4> , 
        \PC<3> , \PC<2> , \PC<1> , \PC<0> }), .jump(jump), .jumpReg(jumpReg), 
        .branch(branch), .nextPC({\nextPC<15> , \nextPC<14> , \nextPC<13> , 
        \nextPC<12> , \nextPC<11> , \nextPC<10> , \nextPC<9> , \nextPC<8> , 
        \nextPC<7> , \nextPC<6> , \nextPC<5> , \nextPC<4> , \nextPC<3> , 
        \nextPC<2> , \nextPC<1> , \nextPC<0> }), .ALURes({\ALURes<15> , 
        \ALURes<14> , \ALURes<13> , \ALURes<12> , \ALURes<11> , \ALURes<10> , 
        \ALURes<9> , \ALURes<8> , \ALURes<7> , \ALURes<6> , \ALURes<5> , 
        \ALURes<4> , \ALURes<3> , \ALURes<2> , \ALURes<1> , \ALURes<0> }), 
        .passthrough(passthrough), .reverse(reverse), .err() );
  memory memory0 ( .clk(clk), .rst(n19), .addr({\ALURes<15> , \ALURes<14> , 
        \ALURes<13> , \ALURes<12> , \ALURes<11> , \ALURes<10> , \ALURes<9> , 
        \ALURes<8> , \ALURes<7> , \ALURes<6> , \ALURes<5> , \ALURes<4> , 
        \ALURes<3> , \ALURes<2> , \ALURes<1> , \ALURes<0> }), .writeData({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .halt(halt), .memWrite(memWrite), .memRead(memRead), .readData({\readData<15> , \readData<14> , \readData<13> , \readData<12> , 
        \readData<11> , \readData<10> , \readData<9> , \readData<8> , 
        \readData<7> , \readData<6> , \readData<5> , \readData<4> , 
        \readData<3> , \readData<2> , \readData<1> , \readData<0> }), .err()
         );
  writeBack wb0 ( .memData({\readData<15> , \readData<14> , \readData<13> , 
        \readData<12> , \readData<11> , \readData<10> , \readData<9> , 
        \readData<8> , \readData<7> , \readData<6> , \readData<5> , 
        \readData<4> , \readData<3> , \readData<2> , \readData<1> , 
        \readData<0> }), .ALUData({n6, n13, n12, \ALURes<12> , \ALURes<11> , 
        n17, \ALURes<9> , \ALURes<8> , n11, n15, n10, \ALURes<4> , n4, n5, n8, 
        n14}), .memToReg(memToReg), .writeBackData({\writeBackData<15> , 
        \writeBackData<14> , \writeBackData<13> , \writeBackData<12> , 
        \writeBackData<11> , \writeBackData<10> , \writeBackData<9> , 
        \writeBackData<8> , \writeBackData<7> , \writeBackData<6> , 
        \writeBackData<5> , \writeBackData<4> , \writeBackData<3> , 
        \writeBackData<2> , \writeBackData<1> , \writeBackData<0> }), .err()
         );
  INVX1 U5 ( .A(n20), .Y(n19) );
  INVX1 U6 ( .A(rst), .Y(n20) );
  BUFX2 U7 ( .A(\ALURes<3> ), .Y(n4) );
  BUFX2 U8 ( .A(\ALURes<2> ), .Y(n5) );
  BUFX2 U9 ( .A(\ALURes<15> ), .Y(n6) );
  INVX1 U10 ( .A(\ALURes<1> ), .Y(n7) );
  INVX1 U11 ( .A(n7), .Y(n8) );
  INVX1 U12 ( .A(\ALURes<5> ), .Y(n9) );
  INVX1 U13 ( .A(n9), .Y(n10) );
  BUFX2 U14 ( .A(\ALURes<7> ), .Y(n11) );
  BUFX2 U15 ( .A(\ALURes<13> ), .Y(n12) );
  BUFX2 U16 ( .A(\ALURes<14> ), .Y(n13) );
  BUFX2 U17 ( .A(\ALURes<0> ), .Y(n14) );
  INVX1 U18 ( .A(n16), .Y(n15) );
  INVX1 U19 ( .A(\ALURes<6> ), .Y(n16) );
  BUFX2 U20 ( .A(\ALURes<10> ), .Y(n17) );
endmodule

