module execute(readdata1, readdata2, immediate, ALUOp, ALUSrc, jump, jumpReg, branch, nextPC, ALURes, err);
	
endmodule
