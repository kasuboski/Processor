library verilog;
use verilog.vl_types.all;
entity comparator_tb is
end comparator_tb;
